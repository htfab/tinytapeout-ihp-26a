module tt_um_herald (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _00000_;
 wire _00001_;
 wire _00002_;
 wire _00003_;
 wire _00004_;
 wire _00005_;
 wire _00006_;
 wire _00007_;
 wire _00008_;
 wire _00009_;
 wire _00010_;
 wire _00011_;
 wire _00012_;
 wire _00013_;
 wire _00014_;
 wire _00015_;
 wire _00016_;
 wire _00017_;
 wire _00018_;
 wire _00019_;
 wire _00020_;
 wire _00021_;
 wire _00022_;
 wire _00023_;
 wire _00024_;
 wire _00025_;
 wire _00026_;
 wire _00027_;
 wire _00028_;
 wire _00029_;
 wire _00030_;
 wire _00031_;
 wire _00032_;
 wire _00033_;
 wire _00034_;
 wire _00035_;
 wire _00036_;
 wire _00037_;
 wire _00038_;
 wire _00039_;
 wire _00040_;
 wire _00041_;
 wire _00042_;
 wire _00043_;
 wire _00044_;
 wire _00045_;
 wire _00046_;
 wire _00047_;
 wire _00048_;
 wire _00049_;
 wire _00050_;
 wire _00051_;
 wire _00052_;
 wire _00053_;
 wire _00054_;
 wire _00055_;
 wire _00056_;
 wire _00057_;
 wire _00058_;
 wire _00059_;
 wire _00060_;
 wire _00061_;
 wire _00062_;
 wire _00063_;
 wire _00064_;
 wire _00065_;
 wire _00066_;
 wire _00067_;
 wire _00068_;
 wire _00069_;
 wire _00070_;
 wire _00071_;
 wire _00072_;
 wire _00073_;
 wire _00074_;
 wire _00075_;
 wire _00076_;
 wire _00077_;
 wire _00078_;
 wire _00079_;
 wire _00080_;
 wire _00081_;
 wire _00082_;
 wire _00083_;
 wire _00084_;
 wire _00085_;
 wire _00086_;
 wire _00087_;
 wire _00088_;
 wire _00089_;
 wire _00090_;
 wire _00091_;
 wire _00092_;
 wire _00093_;
 wire _00094_;
 wire _00095_;
 wire _00096_;
 wire _00097_;
 wire _00098_;
 wire _00099_;
 wire _00100_;
 wire _00101_;
 wire _00102_;
 wire _00103_;
 wire _00104_;
 wire _00105_;
 wire _00106_;
 wire _00107_;
 wire _00108_;
 wire _00109_;
 wire _00110_;
 wire _00111_;
 wire _00112_;
 wire _00113_;
 wire _00114_;
 wire _00115_;
 wire _00116_;
 wire _00117_;
 wire _00118_;
 wire _00119_;
 wire _00120_;
 wire _00121_;
 wire _00122_;
 wire _00123_;
 wire _00124_;
 wire _00125_;
 wire _00126_;
 wire _00127_;
 wire _00128_;
 wire _00129_;
 wire _00130_;
 wire _00131_;
 wire _00132_;
 wire _00133_;
 wire _00134_;
 wire _00135_;
 wire _00136_;
 wire _00137_;
 wire _00138_;
 wire _00139_;
 wire _00140_;
 wire _00141_;
 wire _00142_;
 wire _00143_;
 wire _00144_;
 wire _00145_;
 wire _00146_;
 wire _00147_;
 wire _00148_;
 wire _00149_;
 wire _00150_;
 wire _00151_;
 wire _00152_;
 wire _00153_;
 wire _00154_;
 wire _00155_;
 wire _00156_;
 wire _00157_;
 wire _00158_;
 wire _00159_;
 wire _00160_;
 wire _00161_;
 wire _00162_;
 wire _00163_;
 wire _00164_;
 wire _00165_;
 wire _00166_;
 wire _00167_;
 wire _00168_;
 wire _00169_;
 wire _00170_;
 wire _00171_;
 wire _00172_;
 wire _00173_;
 wire _00174_;
 wire _00175_;
 wire _00176_;
 wire _00177_;
 wire _00178_;
 wire _00179_;
 wire _00180_;
 wire _00181_;
 wire _00182_;
 wire _00183_;
 wire _00184_;
 wire _00185_;
 wire _00186_;
 wire _00187_;
 wire _00188_;
 wire _00189_;
 wire _00190_;
 wire _00191_;
 wire _00192_;
 wire _00193_;
 wire _00194_;
 wire _00195_;
 wire _00196_;
 wire _00197_;
 wire _00198_;
 wire _00199_;
 wire _00200_;
 wire _00201_;
 wire _00202_;
 wire _00203_;
 wire _00204_;
 wire _00205_;
 wire _00206_;
 wire _00207_;
 wire _00208_;
 wire _00209_;
 wire _00210_;
 wire _00211_;
 wire _00212_;
 wire _00213_;
 wire _00214_;
 wire _00215_;
 wire _00216_;
 wire _00217_;
 wire _00218_;
 wire _00219_;
 wire _00220_;
 wire _00221_;
 wire _00222_;
 wire _00223_;
 wire _00224_;
 wire _00225_;
 wire _00226_;
 wire _00227_;
 wire _00228_;
 wire _00229_;
 wire _00230_;
 wire _00231_;
 wire _00232_;
 wire _00233_;
 wire _00234_;
 wire _00235_;
 wire _00236_;
 wire _00237_;
 wire _00238_;
 wire _00239_;
 wire _00240_;
 wire _00241_;
 wire _00242_;
 wire _00243_;
 wire _00244_;
 wire _00245_;
 wire _00246_;
 wire _00247_;
 wire _00248_;
 wire _00249_;
 wire _00250_;
 wire _00251_;
 wire _00252_;
 wire _00253_;
 wire _00254_;
 wire _00255_;
 wire _00256_;
 wire _00257_;
 wire _00258_;
 wire _00259_;
 wire _00260_;
 wire _00261_;
 wire _00262_;
 wire _00263_;
 wire _00264_;
 wire _00265_;
 wire _00266_;
 wire _00267_;
 wire _00268_;
 wire _00269_;
 wire _00270_;
 wire _00271_;
 wire _00272_;
 wire _00273_;
 wire _00274_;
 wire _00275_;
 wire _00276_;
 wire _00277_;
 wire _00278_;
 wire _00279_;
 wire _00280_;
 wire _00281_;
 wire _00282_;
 wire _00283_;
 wire _00284_;
 wire _00285_;
 wire _00286_;
 wire _00287_;
 wire _00288_;
 wire _00289_;
 wire _00290_;
 wire _00291_;
 wire _00292_;
 wire _00293_;
 wire _00294_;
 wire _00295_;
 wire _00296_;
 wire _00297_;
 wire _00298_;
 wire _00299_;
 wire _00300_;
 wire _00301_;
 wire _00302_;
 wire _00303_;
 wire _00304_;
 wire _00305_;
 wire _00306_;
 wire _00307_;
 wire _00308_;
 wire _00309_;
 wire _00310_;
 wire _00311_;
 wire _00312_;
 wire _00313_;
 wire _00314_;
 wire _00315_;
 wire _00316_;
 wire _00317_;
 wire _00318_;
 wire _00319_;
 wire _00320_;
 wire _00321_;
 wire _00322_;
 wire _00323_;
 wire _00324_;
 wire _00325_;
 wire _00326_;
 wire _00327_;
 wire _00328_;
 wire _00329_;
 wire _00330_;
 wire _00331_;
 wire _00332_;
 wire _00333_;
 wire _00334_;
 wire _00335_;
 wire _00336_;
 wire _00337_;
 wire _00338_;
 wire _00339_;
 wire _00340_;
 wire _00341_;
 wire _00342_;
 wire _00343_;
 wire _00344_;
 wire _00345_;
 wire _00346_;
 wire _00347_;
 wire _00348_;
 wire _00349_;
 wire _00350_;
 wire _00351_;
 wire _00352_;
 wire _00353_;
 wire _00354_;
 wire _00355_;
 wire _00356_;
 wire _00357_;
 wire _00358_;
 wire _00359_;
 wire _00360_;
 wire _00361_;
 wire _00362_;
 wire _00363_;
 wire _00364_;
 wire _00365_;
 wire _00366_;
 wire _00367_;
 wire _00368_;
 wire _00369_;
 wire _00370_;
 wire _00371_;
 wire _00372_;
 wire _00373_;
 wire _00374_;
 wire _00375_;
 wire _00376_;
 wire _00377_;
 wire _00378_;
 wire _00379_;
 wire _00380_;
 wire _00381_;
 wire _00382_;
 wire _00383_;
 wire _00384_;
 wire _00385_;
 wire _00386_;
 wire _00387_;
 wire _00388_;
 wire _00389_;
 wire _00390_;
 wire _00391_;
 wire _00392_;
 wire _00393_;
 wire _00394_;
 wire _00395_;
 wire _00396_;
 wire _00397_;
 wire _00398_;
 wire _00399_;
 wire _00400_;
 wire _00401_;
 wire _00402_;
 wire _00403_;
 wire _00404_;
 wire _00405_;
 wire _00406_;
 wire _00407_;
 wire _00408_;
 wire _00409_;
 wire _00410_;
 wire _00411_;
 wire _00412_;
 wire _00413_;
 wire _00414_;
 wire _00415_;
 wire _00416_;
 wire _00417_;
 wire _00418_;
 wire _00419_;
 wire _00420_;
 wire _00421_;
 wire _00422_;
 wire _00423_;
 wire _00424_;
 wire _00425_;
 wire _00426_;
 wire _00427_;
 wire _00428_;
 wire _00429_;
 wire _00430_;
 wire _00431_;
 wire _00432_;
 wire _00433_;
 wire _00434_;
 wire _00435_;
 wire _00436_;
 wire _00437_;
 wire _00438_;
 wire _00439_;
 wire _00440_;
 wire _00441_;
 wire _00442_;
 wire _00443_;
 wire _00444_;
 wire _00445_;
 wire _00446_;
 wire _00447_;
 wire _00448_;
 wire _00449_;
 wire _00450_;
 wire _00451_;
 wire _00452_;
 wire _00453_;
 wire _00454_;
 wire _00455_;
 wire _00456_;
 wire _00457_;
 wire _00458_;
 wire _00459_;
 wire _00460_;
 wire _00461_;
 wire _00462_;
 wire _00463_;
 wire _00464_;
 wire _00465_;
 wire _00466_;
 wire _00467_;
 wire _00468_;
 wire _00469_;
 wire _00470_;
 wire _00471_;
 wire _00472_;
 wire _00473_;
 wire _00474_;
 wire _00475_;
 wire _00476_;
 wire _00477_;
 wire _00478_;
 wire _00479_;
 wire _00480_;
 wire _00481_;
 wire _00482_;
 wire _00483_;
 wire _00484_;
 wire _00485_;
 wire _00486_;
 wire _00487_;
 wire _00488_;
 wire _00489_;
 wire _00490_;
 wire _00491_;
 wire _00492_;
 wire _00493_;
 wire _00494_;
 wire _00495_;
 wire _00496_;
 wire _00497_;
 wire _00498_;
 wire _00499_;
 wire _00500_;
 wire _00501_;
 wire _00502_;
 wire _00503_;
 wire _00504_;
 wire _00505_;
 wire _00506_;
 wire _00507_;
 wire _00508_;
 wire _00509_;
 wire _00510_;
 wire _00511_;
 wire _00512_;
 wire _00513_;
 wire _00514_;
 wire _00515_;
 wire _00516_;
 wire _00517_;
 wire _00518_;
 wire _00519_;
 wire _00520_;
 wire _00521_;
 wire _00522_;
 wire _00523_;
 wire _00524_;
 wire _00525_;
 wire _00526_;
 wire _00527_;
 wire _00528_;
 wire _00529_;
 wire _00530_;
 wire _00531_;
 wire _00532_;
 wire _00533_;
 wire _00534_;
 wire _00535_;
 wire _00536_;
 wire _00537_;
 wire _00538_;
 wire _00539_;
 wire _00540_;
 wire _00541_;
 wire _00542_;
 wire _00543_;
 wire _00544_;
 wire _00545_;
 wire _00546_;
 wire _00547_;
 wire _00548_;
 wire _00549_;
 wire _00550_;
 wire _00551_;
 wire _00552_;
 wire _00553_;
 wire _00554_;
 wire _00555_;
 wire _00556_;
 wire _00557_;
 wire _00558_;
 wire _00559_;
 wire _00560_;
 wire _00561_;
 wire _00562_;
 wire _00563_;
 wire _00564_;
 wire _00565_;
 wire _00566_;
 wire _00567_;
 wire _00568_;
 wire _00569_;
 wire _00570_;
 wire _00571_;
 wire _00572_;
 wire _00573_;
 wire _00574_;
 wire _00575_;
 wire _00576_;
 wire _00577_;
 wire _00578_;
 wire _00579_;
 wire _00580_;
 wire _00581_;
 wire _00582_;
 wire _00583_;
 wire _00584_;
 wire _00585_;
 wire _00586_;
 wire _00587_;
 wire _00588_;
 wire _00589_;
 wire _00590_;
 wire _00591_;
 wire _00592_;
 wire _00593_;
 wire _00594_;
 wire _00595_;
 wire _00596_;
 wire _00597_;
 wire _00598_;
 wire _00599_;
 wire _00600_;
 wire _00601_;
 wire _00602_;
 wire _00603_;
 wire _00604_;
 wire _00605_;
 wire _00606_;
 wire _00607_;
 wire _00608_;
 wire _00609_;
 wire _00610_;
 wire _00611_;
 wire _00612_;
 wire _00613_;
 wire _00614_;
 wire _00615_;
 wire _00616_;
 wire _00617_;
 wire _00618_;
 wire _00619_;
 wire _00620_;
 wire _00621_;
 wire _00622_;
 wire _00623_;
 wire _00624_;
 wire _00625_;
 wire _00626_;
 wire _00627_;
 wire _00628_;
 wire _00629_;
 wire _00630_;
 wire _00631_;
 wire _00632_;
 wire _00633_;
 wire _00634_;
 wire _00635_;
 wire _00636_;
 wire _00637_;
 wire _00638_;
 wire _00639_;
 wire _00640_;
 wire _00641_;
 wire _00642_;
 wire _00643_;
 wire _00644_;
 wire _00645_;
 wire _00646_;
 wire _00647_;
 wire _00648_;
 wire _00649_;
 wire _00650_;
 wire _00651_;
 wire _00652_;
 wire _00653_;
 wire _00654_;
 wire _00655_;
 wire _00656_;
 wire _00657_;
 wire _00658_;
 wire _00659_;
 wire _00660_;
 wire _00661_;
 wire _00662_;
 wire _00663_;
 wire _00664_;
 wire _00665_;
 wire _00666_;
 wire _00667_;
 wire _00668_;
 wire _00669_;
 wire _00670_;
 wire _00671_;
 wire _00672_;
 wire _00673_;
 wire _00674_;
 wire _00675_;
 wire _00676_;
 wire _00677_;
 wire _00678_;
 wire _00679_;
 wire _00680_;
 wire _00681_;
 wire _00682_;
 wire _00683_;
 wire _00684_;
 wire _00685_;
 wire _00686_;
 wire _00687_;
 wire _00688_;
 wire _00689_;
 wire _00690_;
 wire _00691_;
 wire _00692_;
 wire _00693_;
 wire _00694_;
 wire _00695_;
 wire _00696_;
 wire _00697_;
 wire _00698_;
 wire _00699_;
 wire _00700_;
 wire _00701_;
 wire _00702_;
 wire _00703_;
 wire _00704_;
 wire _00705_;
 wire _00706_;
 wire _00707_;
 wire _00708_;
 wire _00709_;
 wire _00710_;
 wire _00711_;
 wire _00712_;
 wire _00713_;
 wire _00714_;
 wire _00715_;
 wire _00716_;
 wire _00717_;
 wire _00718_;
 wire _00719_;
 wire _00720_;
 wire _00721_;
 wire _00722_;
 wire _00723_;
 wire _00724_;
 wire _00725_;
 wire _00726_;
 wire _00727_;
 wire _00728_;
 wire _00729_;
 wire _00730_;
 wire _00731_;
 wire _00732_;
 wire _00733_;
 wire _00734_;
 wire _00735_;
 wire _00736_;
 wire _00737_;
 wire _00738_;
 wire _00739_;
 wire _00740_;
 wire _00741_;
 wire _00742_;
 wire _00743_;
 wire _00744_;
 wire _00745_;
 wire _00746_;
 wire _00747_;
 wire _00748_;
 wire _00749_;
 wire _00750_;
 wire _00751_;
 wire _00752_;
 wire _00753_;
 wire _00754_;
 wire _00755_;
 wire _00756_;
 wire _00757_;
 wire _00758_;
 wire _00759_;
 wire _00760_;
 wire _00761_;
 wire _00762_;
 wire _00763_;
 wire _00764_;
 wire _00765_;
 wire _00766_;
 wire _00767_;
 wire _00768_;
 wire _00769_;
 wire _00770_;
 wire _00771_;
 wire _00772_;
 wire _00773_;
 wire _00774_;
 wire _00775_;
 wire _00776_;
 wire _00777_;
 wire _00778_;
 wire _00779_;
 wire _00780_;
 wire _00781_;
 wire _00782_;
 wire _00783_;
 wire _00784_;
 wire _00785_;
 wire _00786_;
 wire _00787_;
 wire _00788_;
 wire _00789_;
 wire _00790_;
 wire _00791_;
 wire _00792_;
 wire _00793_;
 wire _00794_;
 wire _00795_;
 wire _00796_;
 wire _00797_;
 wire _00798_;
 wire _00799_;
 wire _00800_;
 wire _00801_;
 wire _00802_;
 wire _00803_;
 wire _00804_;
 wire _00805_;
 wire _00806_;
 wire _00807_;
 wire _00808_;
 wire _00809_;
 wire _00810_;
 wire _00811_;
 wire _00812_;
 wire _00813_;
 wire _00814_;
 wire _00815_;
 wire _00816_;
 wire _00817_;
 wire _00818_;
 wire _00819_;
 wire _00820_;
 wire _00821_;
 wire _00822_;
 wire _00823_;
 wire _00824_;
 wire _00825_;
 wire _00826_;
 wire _00827_;
 wire _00828_;
 wire _00829_;
 wire _00830_;
 wire _00831_;
 wire _00832_;
 wire _00833_;
 wire _00834_;
 wire _00835_;
 wire _00836_;
 wire _00837_;
 wire _00838_;
 wire _00839_;
 wire _00840_;
 wire _00841_;
 wire _00842_;
 wire _00843_;
 wire _00844_;
 wire _00845_;
 wire _00846_;
 wire _00847_;
 wire _00848_;
 wire _00849_;
 wire _00850_;
 wire _00851_;
 wire _00852_;
 wire _00853_;
 wire _00854_;
 wire _00855_;
 wire _00856_;
 wire _00857_;
 wire _00858_;
 wire _00859_;
 wire _00860_;
 wire _00861_;
 wire _00862_;
 wire _00863_;
 wire _00864_;
 wire _00865_;
 wire _00866_;
 wire _00867_;
 wire _00868_;
 wire _00869_;
 wire _00870_;
 wire _00871_;
 wire _00872_;
 wire _00873_;
 wire _00874_;
 wire _00875_;
 wire _00876_;
 wire _00877_;
 wire _00878_;
 wire _00879_;
 wire _00880_;
 wire _00881_;
 wire _00882_;
 wire _00883_;
 wire _00884_;
 wire _00885_;
 wire _00886_;
 wire _00887_;
 wire _00888_;
 wire _00889_;
 wire _00890_;
 wire _00891_;
 wire _00892_;
 wire _00893_;
 wire _00894_;
 wire _00895_;
 wire _00896_;
 wire _00897_;
 wire _00898_;
 wire _00899_;
 wire _00900_;
 wire _00901_;
 wire _00902_;
 wire _00903_;
 wire _00904_;
 wire _00905_;
 wire _00906_;
 wire _00907_;
 wire _00908_;
 wire _00909_;
 wire _00910_;
 wire _00911_;
 wire _00912_;
 wire _00913_;
 wire _00914_;
 wire _00915_;
 wire _00916_;
 wire _00917_;
 wire _00918_;
 wire _00919_;
 wire _00920_;
 wire _00921_;
 wire _00922_;
 wire _00923_;
 wire _00924_;
 wire _00925_;
 wire _00926_;
 wire _00927_;
 wire _00928_;
 wire _00929_;
 wire _00930_;
 wire _00931_;
 wire _00932_;
 wire _00933_;
 wire _00934_;
 wire _00935_;
 wire _00936_;
 wire _00937_;
 wire _00938_;
 wire _00939_;
 wire _00940_;
 wire _00941_;
 wire _00942_;
 wire _00943_;
 wire _00944_;
 wire _00945_;
 wire _00946_;
 wire _00947_;
 wire _00948_;
 wire _00949_;
 wire _00950_;
 wire _00951_;
 wire _00952_;
 wire _00953_;
 wire _00954_;
 wire _00955_;
 wire _00956_;
 wire _00957_;
 wire _00958_;
 wire _00959_;
 wire _00960_;
 wire _00961_;
 wire _00962_;
 wire _00963_;
 wire _00964_;
 wire _00965_;
 wire _00966_;
 wire _00967_;
 wire _00968_;
 wire _00969_;
 wire _00970_;
 wire _00971_;
 wire _00972_;
 wire _00973_;
 wire _00974_;
 wire _00975_;
 wire _00976_;
 wire _00977_;
 wire _00978_;
 wire _00979_;
 wire _00980_;
 wire _00981_;
 wire _00982_;
 wire _00983_;
 wire _00984_;
 wire _00985_;
 wire _00986_;
 wire _00987_;
 wire _00988_;
 wire _00989_;
 wire _00990_;
 wire _00991_;
 wire _00992_;
 wire _00993_;
 wire _00994_;
 wire _00995_;
 wire _00996_;
 wire _00997_;
 wire _00998_;
 wire _00999_;
 wire _01000_;
 wire _01001_;
 wire _01002_;
 wire _01003_;
 wire _01004_;
 wire _01005_;
 wire _01006_;
 wire _01007_;
 wire _01008_;
 wire _01009_;
 wire _01010_;
 wire _01011_;
 wire _01012_;
 wire _01013_;
 wire _01014_;
 wire _01015_;
 wire _01016_;
 wire _01017_;
 wire _01018_;
 wire _01019_;
 wire _01020_;
 wire _01021_;
 wire _01022_;
 wire _01023_;
 wire _01024_;
 wire _01025_;
 wire _01026_;
 wire _01027_;
 wire _01028_;
 wire _01029_;
 wire _01030_;
 wire _01031_;
 wire _01032_;
 wire _01033_;
 wire _01034_;
 wire _01035_;
 wire _01036_;
 wire _01037_;
 wire _01038_;
 wire _01039_;
 wire _01040_;
 wire _01041_;
 wire _01042_;
 wire _01043_;
 wire _01044_;
 wire _01045_;
 wire _01046_;
 wire _01047_;
 wire _01048_;
 wire _01049_;
 wire _01050_;
 wire _01051_;
 wire _01052_;
 wire _01053_;
 wire _01054_;
 wire _01055_;
 wire _01056_;
 wire _01057_;
 wire _01058_;
 wire _01059_;
 wire _01060_;
 wire _01061_;
 wire _01062_;
 wire _01063_;
 wire _01064_;
 wire _01065_;
 wire _01066_;
 wire _01067_;
 wire _01068_;
 wire _01069_;
 wire _01070_;
 wire _01071_;
 wire _01072_;
 wire _01073_;
 wire _01074_;
 wire _01075_;
 wire _01076_;
 wire _01077_;
 wire _01078_;
 wire _01079_;
 wire _01080_;
 wire _01081_;
 wire _01082_;
 wire _01083_;
 wire _01084_;
 wire _01085_;
 wire _01086_;
 wire _01087_;
 wire _01088_;
 wire _01089_;
 wire _01090_;
 wire _01091_;
 wire _01092_;
 wire _01093_;
 wire _01094_;
 wire _01095_;
 wire _01096_;
 wire _01097_;
 wire _01098_;
 wire _01099_;
 wire _01100_;
 wire _01101_;
 wire _01102_;
 wire _01103_;
 wire _01104_;
 wire _01105_;
 wire _01106_;
 wire _01107_;
 wire _01108_;
 wire _01109_;
 wire _01110_;
 wire _01111_;
 wire _01112_;
 wire _01113_;
 wire _01114_;
 wire _01115_;
 wire _01116_;
 wire _01117_;
 wire _01118_;
 wire _01119_;
 wire _01120_;
 wire _01121_;
 wire _01122_;
 wire _01123_;
 wire _01124_;
 wire _01125_;
 wire _01126_;
 wire _01127_;
 wire _01128_;
 wire _01129_;
 wire _01130_;
 wire _01131_;
 wire _01132_;
 wire _01133_;
 wire _01134_;
 wire _01135_;
 wire _01136_;
 wire _01137_;
 wire _01138_;
 wire _01139_;
 wire _01140_;
 wire _01141_;
 wire _01142_;
 wire _01143_;
 wire _01144_;
 wire _01145_;
 wire _01146_;
 wire _01147_;
 wire _01148_;
 wire _01149_;
 wire _01150_;
 wire _01151_;
 wire _01152_;
 wire _01153_;
 wire _01154_;
 wire _01155_;
 wire _01156_;
 wire _01157_;
 wire _01158_;
 wire _01159_;
 wire _01160_;
 wire _01161_;
 wire _01162_;
 wire _01163_;
 wire _01164_;
 wire _01165_;
 wire _01166_;
 wire _01167_;
 wire _01168_;
 wire _01169_;
 wire _01170_;
 wire _01171_;
 wire _01172_;
 wire _01173_;
 wire _01174_;
 wire _01175_;
 wire _01176_;
 wire _01177_;
 wire _01178_;
 wire _01179_;
 wire _01180_;
 wire _01181_;
 wire _01182_;
 wire _01183_;
 wire _01184_;
 wire _01185_;
 wire _01186_;
 wire _01187_;
 wire _01188_;
 wire _01189_;
 wire _01190_;
 wire _01191_;
 wire _01192_;
 wire _01193_;
 wire _01194_;
 wire _01195_;
 wire _01196_;
 wire _01197_;
 wire _01198_;
 wire _01199_;
 wire _01200_;
 wire _01201_;
 wire _01202_;
 wire _01203_;
 wire _01204_;
 wire _01205_;
 wire _01206_;
 wire _01207_;
 wire _01208_;
 wire _01209_;
 wire _01210_;
 wire _01211_;
 wire _01212_;
 wire _01213_;
 wire _01214_;
 wire _01215_;
 wire _01216_;
 wire _01217_;
 wire _01218_;
 wire _01219_;
 wire _01220_;
 wire _01221_;
 wire _01222_;
 wire _01223_;
 wire _01224_;
 wire _01225_;
 wire _01226_;
 wire _01227_;
 wire _01228_;
 wire _01229_;
 wire _01230_;
 wire _01231_;
 wire _01232_;
 wire _01233_;
 wire _01234_;
 wire _01235_;
 wire _01236_;
 wire _01237_;
 wire _01238_;
 wire _01239_;
 wire _01240_;
 wire _01241_;
 wire _01242_;
 wire _01243_;
 wire _01244_;
 wire _01245_;
 wire _01246_;
 wire _01247_;
 wire _01248_;
 wire _01249_;
 wire _01250_;
 wire _01251_;
 wire _01252_;
 wire _01253_;
 wire _01254_;
 wire _01255_;
 wire _01256_;
 wire _01257_;
 wire _01258_;
 wire _01259_;
 wire _01260_;
 wire _01261_;
 wire _01262_;
 wire _01263_;
 wire _01264_;
 wire _01265_;
 wire _01266_;
 wire _01267_;
 wire _01268_;
 wire _01269_;
 wire _01270_;
 wire _01271_;
 wire _01272_;
 wire _01273_;
 wire _01274_;
 wire _01275_;
 wire _01276_;
 wire _01277_;
 wire _01278_;
 wire _01279_;
 wire _01280_;
 wire _01281_;
 wire _01282_;
 wire _01283_;
 wire _01284_;
 wire _01285_;
 wire _01286_;
 wire _01287_;
 wire _01288_;
 wire _01289_;
 wire _01290_;
 wire _01291_;
 wire _01292_;
 wire _01293_;
 wire _01294_;
 wire _01295_;
 wire _01296_;
 wire _01297_;
 wire _01298_;
 wire _01299_;
 wire _01300_;
 wire _01301_;
 wire _01302_;
 wire _01303_;
 wire _01304_;
 wire _01305_;
 wire _01306_;
 wire _01307_;
 wire _01308_;
 wire _01309_;
 wire _01310_;
 wire _01311_;
 wire _01312_;
 wire _01313_;
 wire _01314_;
 wire _01315_;
 wire _01316_;
 wire _01317_;
 wire _01318_;
 wire _01319_;
 wire _01320_;
 wire _01321_;
 wire _01322_;
 wire _01323_;
 wire _01324_;
 wire _01325_;
 wire _01326_;
 wire _01327_;
 wire _01328_;
 wire _01329_;
 wire _01330_;
 wire _01331_;
 wire _01332_;
 wire _01333_;
 wire _01334_;
 wire _01335_;
 wire _01336_;
 wire _01337_;
 wire _01338_;
 wire _01339_;
 wire _01340_;
 wire _01341_;
 wire _01342_;
 wire _01343_;
 wire _01344_;
 wire _01345_;
 wire _01346_;
 wire _01347_;
 wire _01348_;
 wire _01349_;
 wire _01350_;
 wire _01351_;
 wire _01352_;
 wire _01353_;
 wire _01354_;
 wire _01355_;
 wire _01356_;
 wire _01357_;
 wire _01358_;
 wire _01359_;
 wire _01360_;
 wire _01361_;
 wire _01362_;
 wire _01363_;
 wire _01364_;
 wire _01365_;
 wire _01366_;
 wire _01367_;
 wire _01368_;
 wire _01369_;
 wire _01370_;
 wire _01371_;
 wire _01372_;
 wire _01373_;
 wire _01374_;
 wire _01375_;
 wire _01376_;
 wire _01377_;
 wire _01378_;
 wire _01379_;
 wire _01380_;
 wire _01381_;
 wire _01382_;
 wire _01383_;
 wire _01384_;
 wire _01385_;
 wire _01386_;
 wire _01387_;
 wire _01388_;
 wire _01389_;
 wire _01390_;
 wire _01391_;
 wire _01392_;
 wire _01393_;
 wire _01394_;
 wire _01395_;
 wire _01396_;
 wire _01397_;
 wire _01398_;
 wire _01399_;
 wire _01400_;
 wire _01401_;
 wire _01402_;
 wire _01403_;
 wire _01404_;
 wire _01405_;
 wire _01406_;
 wire _01407_;
 wire _01408_;
 wire _01409_;
 wire _01410_;
 wire _01411_;
 wire _01412_;
 wire _01413_;
 wire _01414_;
 wire _01415_;
 wire _01416_;
 wire _01417_;
 wire _01418_;
 wire _01419_;
 wire _01420_;
 wire _01421_;
 wire _01422_;
 wire _01423_;
 wire _01424_;
 wire _01425_;
 wire _01426_;
 wire _01427_;
 wire _01428_;
 wire _01429_;
 wire _01430_;
 wire _01431_;
 wire _01432_;
 wire _01433_;
 wire _01434_;
 wire _01435_;
 wire _01436_;
 wire _01437_;
 wire _01438_;
 wire _01439_;
 wire _01440_;
 wire _01441_;
 wire _01442_;
 wire _01443_;
 wire _01444_;
 wire _01445_;
 wire _01446_;
 wire _01447_;
 wire _01448_;
 wire _01449_;
 wire _01450_;
 wire _01451_;
 wire _01452_;
 wire _01453_;
 wire _01454_;
 wire _01455_;
 wire _01456_;
 wire _01457_;
 wire _01458_;
 wire _01459_;
 wire _01460_;
 wire _01461_;
 wire _01462_;
 wire _01463_;
 wire _01464_;
 wire _01465_;
 wire _01466_;
 wire _01467_;
 wire _01468_;
 wire _01469_;
 wire _01470_;
 wire _01471_;
 wire _01472_;
 wire _01473_;
 wire _01474_;
 wire _01475_;
 wire _01476_;
 wire _01477_;
 wire _01478_;
 wire _01479_;
 wire _01480_;
 wire _01481_;
 wire _01482_;
 wire _01483_;
 wire _01484_;
 wire _01485_;
 wire _01486_;
 wire _01487_;
 wire _01488_;
 wire _01489_;
 wire _01490_;
 wire _01491_;
 wire _01492_;
 wire _01493_;
 wire _01494_;
 wire _01495_;
 wire _01496_;
 wire _01497_;
 wire _01498_;
 wire _01499_;
 wire _01500_;
 wire _01501_;
 wire _01502_;
 wire _01503_;
 wire _01504_;
 wire _01505_;
 wire _01506_;
 wire _01507_;
 wire _01508_;
 wire _01509_;
 wire _01510_;
 wire _01511_;
 wire _01512_;
 wire _01513_;
 wire _01514_;
 wire _01515_;
 wire _01516_;
 wire _01517_;
 wire _01518_;
 wire _01519_;
 wire _01520_;
 wire _01521_;
 wire _01522_;
 wire _01523_;
 wire _01524_;
 wire _01525_;
 wire _01526_;
 wire _01527_;
 wire _01528_;
 wire _01529_;
 wire _01530_;
 wire _01531_;
 wire _01532_;
 wire _01533_;
 wire _01534_;
 wire _01535_;
 wire _01536_;
 wire _01537_;
 wire _01538_;
 wire _01539_;
 wire _01540_;
 wire _01541_;
 wire _01542_;
 wire _01543_;
 wire _01544_;
 wire _01545_;
 wire _01546_;
 wire _01547_;
 wire _01548_;
 wire _01549_;
 wire _01550_;
 wire _01551_;
 wire _01552_;
 wire _01553_;
 wire _01554_;
 wire _01555_;
 wire _01556_;
 wire _01557_;
 wire _01558_;
 wire _01559_;
 wire _01560_;
 wire _01561_;
 wire _01562_;
 wire _01563_;
 wire _01564_;
 wire _01565_;
 wire _01566_;
 wire _01567_;
 wire _01568_;
 wire _01569_;
 wire _01570_;
 wire _01571_;
 wire _01572_;
 wire _01573_;
 wire _01574_;
 wire _01575_;
 wire _01576_;
 wire _01577_;
 wire _01578_;
 wire _01579_;
 wire _01580_;
 wire _01581_;
 wire _01582_;
 wire _01583_;
 wire _01584_;
 wire _01585_;
 wire _01586_;
 wire _01587_;
 wire _01588_;
 wire _01589_;
 wire _01590_;
 wire _01591_;
 wire _01592_;
 wire _01593_;
 wire _01594_;
 wire _01595_;
 wire _01596_;
 wire _01597_;
 wire _01598_;
 wire _01599_;
 wire _01600_;
 wire _01601_;
 wire _01602_;
 wire _01603_;
 wire _01604_;
 wire _01605_;
 wire _01606_;
 wire _01607_;
 wire _01608_;
 wire _01609_;
 wire _01610_;
 wire _01611_;
 wire _01612_;
 wire _01613_;
 wire _01614_;
 wire _01615_;
 wire _01616_;
 wire _01617_;
 wire _01618_;
 wire _01619_;
 wire _01620_;
 wire _01621_;
 wire _01622_;
 wire _01623_;
 wire _01624_;
 wire _01625_;
 wire _01626_;
 wire _01627_;
 wire _01628_;
 wire _01629_;
 wire _01630_;
 wire _01631_;
 wire _01632_;
 wire _01633_;
 wire _01634_;
 wire _01635_;
 wire _01636_;
 wire _01637_;
 wire _01638_;
 wire _01639_;
 wire _01640_;
 wire _01641_;
 wire _01642_;
 wire _01643_;
 wire _01644_;
 wire _01645_;
 wire _01646_;
 wire _01647_;
 wire _01648_;
 wire _01649_;
 wire _01650_;
 wire _01651_;
 wire _01652_;
 wire _01653_;
 wire _01654_;
 wire _01655_;
 wire _01656_;
 wire _01657_;
 wire _01658_;
 wire _01659_;
 wire _01660_;
 wire _01661_;
 wire _01662_;
 wire _01663_;
 wire _01664_;
 wire _01665_;
 wire _01666_;
 wire _01667_;
 wire _01668_;
 wire _01669_;
 wire _01670_;
 wire _01671_;
 wire _01672_;
 wire _01673_;
 wire _01674_;
 wire _01675_;
 wire _01676_;
 wire _01677_;
 wire _01678_;
 wire _01679_;
 wire _01680_;
 wire _01681_;
 wire _01682_;
 wire _01683_;
 wire _01684_;
 wire _01685_;
 wire _01686_;
 wire _01687_;
 wire _01688_;
 wire _01689_;
 wire _01690_;
 wire _01691_;
 wire _01692_;
 wire _01693_;
 wire _01694_;
 wire _01695_;
 wire _01696_;
 wire _01697_;
 wire _01698_;
 wire _01699_;
 wire _01700_;
 wire _01701_;
 wire _01702_;
 wire _01703_;
 wire _01704_;
 wire _01705_;
 wire _01706_;
 wire _01707_;
 wire _01708_;
 wire _01709_;
 wire _01710_;
 wire _01711_;
 wire _01712_;
 wire _01713_;
 wire _01714_;
 wire _01715_;
 wire _01716_;
 wire _01717_;
 wire _01718_;
 wire _01719_;
 wire _01720_;
 wire _01721_;
 wire _01722_;
 wire _01723_;
 wire _01724_;
 wire _01725_;
 wire _01726_;
 wire _01727_;
 wire _01728_;
 wire _01729_;
 wire _01730_;
 wire _01731_;
 wire _01732_;
 wire _01733_;
 wire _01734_;
 wire _01735_;
 wire _01736_;
 wire _01737_;
 wire _01738_;
 wire _01739_;
 wire _01740_;
 wire _01741_;
 wire _01742_;
 wire _01743_;
 wire _01744_;
 wire _01745_;
 wire _01746_;
 wire _01747_;
 wire _01748_;
 wire _01749_;
 wire _01750_;
 wire _01751_;
 wire _01752_;
 wire _01753_;
 wire _01754_;
 wire _01755_;
 wire _01756_;
 wire _01757_;
 wire _01758_;
 wire _01759_;
 wire _01760_;
 wire _01761_;
 wire _01762_;
 wire _01763_;
 wire _01764_;
 wire _01765_;
 wire _01766_;
 wire _01767_;
 wire _01768_;
 wire _01769_;
 wire _01770_;
 wire _01771_;
 wire _01772_;
 wire _01773_;
 wire _01774_;
 wire _01775_;
 wire _01776_;
 wire _01777_;
 wire _01778_;
 wire _01779_;
 wire _01780_;
 wire _01781_;
 wire _01782_;
 wire _01783_;
 wire _01784_;
 wire _01785_;
 wire _01786_;
 wire _01787_;
 wire _01788_;
 wire _01789_;
 wire _01790_;
 wire _01791_;
 wire _01792_;
 wire _01793_;
 wire _01794_;
 wire _01795_;
 wire _01796_;
 wire _01797_;
 wire _01798_;
 wire _01799_;
 wire _01800_;
 wire _01801_;
 wire _01802_;
 wire _01803_;
 wire _01804_;
 wire _01805_;
 wire _01806_;
 wire _01807_;
 wire _01808_;
 wire _01809_;
 wire _01810_;
 wire _01811_;
 wire _01812_;
 wire _01813_;
 wire _01814_;
 wire _01815_;
 wire _01816_;
 wire _01817_;
 wire _01818_;
 wire _01819_;
 wire _01820_;
 wire _01821_;
 wire _01822_;
 wire _01823_;
 wire _01824_;
 wire _01825_;
 wire _01826_;
 wire _01827_;
 wire _01828_;
 wire _01829_;
 wire _01830_;
 wire _01831_;
 wire _01832_;
 wire _01833_;
 wire _01834_;
 wire _01835_;
 wire _01836_;
 wire _01837_;
 wire _01838_;
 wire _01839_;
 wire _01840_;
 wire _01841_;
 wire _01842_;
 wire _01843_;
 wire _01844_;
 wire _01845_;
 wire _01846_;
 wire _01847_;
 wire _01848_;
 wire _01849_;
 wire _01850_;
 wire _01851_;
 wire _01852_;
 wire _01853_;
 wire _01854_;
 wire _01855_;
 wire _01856_;
 wire _01857_;
 wire _01858_;
 wire _01859_;
 wire _01860_;
 wire _01861_;
 wire _01862_;
 wire _01863_;
 wire _01864_;
 wire _01865_;
 wire _01866_;
 wire _01867_;
 wire _01868_;
 wire _01869_;
 wire _01870_;
 wire _01871_;
 wire _01872_;
 wire _01873_;
 wire _01874_;
 wire _01875_;
 wire _01876_;
 wire _01877_;
 wire _01878_;
 wire _01879_;
 wire _01880_;
 wire _01881_;
 wire _01882_;
 wire _01883_;
 wire _01884_;
 wire _01885_;
 wire _01886_;
 wire _01887_;
 wire _01888_;
 wire _01889_;
 wire _01890_;
 wire _01891_;
 wire _01892_;
 wire _01893_;
 wire _01894_;
 wire _01895_;
 wire _01896_;
 wire _01897_;
 wire _01898_;
 wire _01899_;
 wire _01900_;
 wire _01901_;
 wire _01902_;
 wire _01903_;
 wire _01904_;
 wire _01905_;
 wire _01906_;
 wire _01907_;
 wire _01908_;
 wire _01909_;
 wire _01910_;
 wire _01911_;
 wire _01912_;
 wire _01913_;
 wire _01914_;
 wire _01915_;
 wire _01916_;
 wire _01917_;
 wire _01918_;
 wire _01919_;
 wire _01920_;
 wire _01921_;
 wire _01922_;
 wire _01923_;
 wire _01924_;
 wire _01925_;
 wire _01926_;
 wire _01927_;
 wire _01928_;
 wire _01929_;
 wire _01930_;
 wire _01931_;
 wire _01932_;
 wire _01933_;
 wire _01934_;
 wire _01935_;
 wire _01936_;
 wire _01937_;
 wire _01938_;
 wire _01939_;
 wire _01940_;
 wire _01941_;
 wire _01942_;
 wire _01943_;
 wire _01944_;
 wire _01945_;
 wire _01946_;
 wire _01947_;
 wire _01948_;
 wire _01949_;
 wire _01950_;
 wire _01951_;
 wire _01952_;
 wire _01953_;
 wire _01954_;
 wire _01955_;
 wire _01956_;
 wire _01957_;
 wire _01958_;
 wire _01959_;
 wire _01960_;
 wire _01961_;
 wire _01962_;
 wire _01963_;
 wire _01964_;
 wire _01965_;
 wire _01966_;
 wire _01967_;
 wire _01968_;
 wire _01969_;
 wire _01970_;
 wire _01971_;
 wire _01972_;
 wire _01973_;
 wire _01974_;
 wire _01975_;
 wire _01976_;
 wire _01977_;
 wire _01978_;
 wire _01979_;
 wire _01980_;
 wire _01981_;
 wire _01982_;
 wire _01983_;
 wire _01984_;
 wire _01985_;
 wire _01986_;
 wire _01987_;
 wire _01988_;
 wire _01989_;
 wire _01990_;
 wire _01991_;
 wire _01992_;
 wire _01993_;
 wire _01994_;
 wire _01995_;
 wire _01996_;
 wire _01997_;
 wire _01998_;
 wire _01999_;
 wire _02000_;
 wire _02001_;
 wire _02002_;
 wire _02003_;
 wire _02004_;
 wire _02005_;
 wire _02006_;
 wire _02007_;
 wire _02008_;
 wire _02009_;
 wire _02010_;
 wire _02011_;
 wire _02012_;
 wire _02013_;
 wire _02014_;
 wire _02015_;
 wire _02016_;
 wire _02017_;
 wire _02018_;
 wire _02019_;
 wire _02020_;
 wire _02021_;
 wire _02022_;
 wire _02023_;
 wire _02024_;
 wire _02025_;
 wire _02026_;
 wire _02027_;
 wire _02028_;
 wire _02029_;
 wire _02030_;
 wire _02031_;
 wire _02032_;
 wire _02033_;
 wire _02034_;
 wire _02035_;
 wire _02036_;
 wire _02037_;
 wire _02038_;
 wire _02039_;
 wire _02040_;
 wire _02041_;
 wire _02042_;
 wire _02043_;
 wire _02044_;
 wire _02045_;
 wire _02046_;
 wire _02047_;
 wire _02048_;
 wire _02049_;
 wire _02050_;
 wire _02051_;
 wire _02052_;
 wire _02053_;
 wire _02054_;
 wire _02055_;
 wire _02056_;
 wire _02057_;
 wire _02058_;
 wire _02059_;
 wire _02060_;
 wire _02061_;
 wire _02062_;
 wire _02063_;
 wire _02064_;
 wire _02065_;
 wire _02066_;
 wire _02067_;
 wire _02068_;
 wire _02069_;
 wire _02070_;
 wire _02071_;
 wire _02072_;
 wire _02073_;
 wire _02074_;
 wire _02075_;
 wire _02076_;
 wire _02077_;
 wire _02078_;
 wire _02079_;
 wire _02080_;
 wire _02081_;
 wire _02082_;
 wire _02083_;
 wire _02084_;
 wire _02085_;
 wire _02086_;
 wire _02087_;
 wire _02088_;
 wire _02089_;
 wire _02090_;
 wire _02091_;
 wire _02092_;
 wire _02093_;
 wire _02094_;
 wire _02095_;
 wire _02096_;
 wire _02097_;
 wire _02098_;
 wire _02099_;
 wire _02100_;
 wire _02101_;
 wire _02102_;
 wire _02103_;
 wire _02104_;
 wire _02105_;
 wire _02106_;
 wire _02107_;
 wire _02108_;
 wire _02109_;
 wire _02110_;
 wire _02111_;
 wire _02112_;
 wire _02113_;
 wire _02114_;
 wire _02115_;
 wire _02116_;
 wire _02117_;
 wire _02118_;
 wire _02119_;
 wire _02120_;
 wire _02121_;
 wire _02122_;
 wire _02123_;
 wire _02124_;
 wire _02125_;
 wire _02126_;
 wire _02127_;
 wire _02128_;
 wire _02129_;
 wire _02130_;
 wire _02131_;
 wire _02132_;
 wire _02133_;
 wire _02134_;
 wire _02135_;
 wire _02136_;
 wire _02137_;
 wire _02138_;
 wire _02139_;
 wire _02140_;
 wire _02141_;
 wire _02142_;
 wire _02143_;
 wire _02144_;
 wire _02145_;
 wire _02146_;
 wire _02147_;
 wire _02148_;
 wire _02149_;
 wire _02150_;
 wire _02151_;
 wire _02152_;
 wire _02153_;
 wire _02154_;
 wire _02155_;
 wire _02156_;
 wire _02157_;
 wire _02158_;
 wire _02159_;
 wire _02160_;
 wire _02161_;
 wire _02162_;
 wire _02163_;
 wire _02164_;
 wire _02165_;
 wire _02166_;
 wire _02167_;
 wire _02168_;
 wire _02169_;
 wire _02170_;
 wire _02171_;
 wire _02172_;
 wire _02173_;
 wire _02174_;
 wire _02175_;
 wire _02176_;
 wire _02177_;
 wire _02178_;
 wire _02179_;
 wire _02180_;
 wire _02181_;
 wire _02182_;
 wire _02183_;
 wire _02184_;
 wire _02185_;
 wire _02186_;
 wire _02187_;
 wire _02188_;
 wire _02189_;
 wire _02190_;
 wire _02191_;
 wire _02192_;
 wire _02193_;
 wire _02194_;
 wire _02195_;
 wire _02196_;
 wire _02197_;
 wire _02198_;
 wire _02199_;
 wire _02200_;
 wire _02201_;
 wire _02202_;
 wire _02203_;
 wire _02204_;
 wire _02205_;
 wire _02206_;
 wire _02207_;
 wire _02208_;
 wire _02209_;
 wire _02210_;
 wire _02211_;
 wire _02212_;
 wire _02213_;
 wire _02214_;
 wire _02215_;
 wire _02216_;
 wire _02217_;
 wire _02218_;
 wire _02219_;
 wire _02220_;
 wire _02221_;
 wire _02222_;
 wire _02223_;
 wire _02224_;
 wire _02225_;
 wire _02226_;
 wire _02227_;
 wire _02228_;
 wire _02229_;
 wire _02230_;
 wire _02231_;
 wire _02232_;
 wire _02233_;
 wire _02234_;
 wire _02235_;
 wire _02236_;
 wire _02237_;
 wire _02238_;
 wire _02239_;
 wire _02240_;
 wire _02241_;
 wire _02242_;
 wire _02243_;
 wire _02244_;
 wire _02245_;
 wire _02246_;
 wire _02247_;
 wire _02248_;
 wire _02249_;
 wire _02250_;
 wire _02251_;
 wire _02252_;
 wire _02253_;
 wire _02254_;
 wire _02255_;
 wire _02256_;
 wire _02257_;
 wire _02258_;
 wire _02259_;
 wire _02260_;
 wire _02261_;
 wire _02262_;
 wire _02263_;
 wire _02264_;
 wire _02265_;
 wire _02266_;
 wire _02267_;
 wire _02268_;
 wire _02269_;
 wire _02270_;
 wire _02271_;
 wire _02272_;
 wire _02273_;
 wire _02274_;
 wire _02275_;
 wire _02276_;
 wire _02277_;
 wire _02278_;
 wire _02279_;
 wire _02280_;
 wire _02281_;
 wire _02282_;
 wire _02283_;
 wire _02284_;
 wire _02285_;
 wire _02286_;
 wire _02287_;
 wire _02288_;
 wire _02289_;
 wire _02290_;
 wire _02291_;
 wire _02292_;
 wire _02293_;
 wire _02294_;
 wire _02295_;
 wire _02296_;
 wire _02297_;
 wire _02298_;
 wire _02299_;
 wire _02300_;
 wire _02301_;
 wire _02302_;
 wire _02303_;
 wire _02304_;
 wire _02305_;
 wire _02306_;
 wire _02307_;
 wire _02308_;
 wire _02309_;
 wire _02310_;
 wire _02311_;
 wire _02312_;
 wire _02313_;
 wire _02314_;
 wire _02315_;
 wire _02316_;
 wire _02317_;
 wire _02318_;
 wire _02319_;
 wire _02320_;
 wire _02321_;
 wire _02322_;
 wire _02323_;
 wire _02324_;
 wire _02325_;
 wire _02326_;
 wire _02327_;
 wire _02328_;
 wire _02329_;
 wire _02330_;
 wire _02331_;
 wire _02332_;
 wire _02333_;
 wire _02334_;
 wire _02335_;
 wire _02336_;
 wire _02337_;
 wire _02338_;
 wire _02339_;
 wire _02340_;
 wire _02341_;
 wire _02342_;
 wire _02343_;
 wire _02344_;
 wire _02345_;
 wire _02346_;
 wire _02347_;
 wire _02348_;
 wire _02349_;
 wire _02350_;
 wire _02351_;
 wire _02352_;
 wire _02353_;
 wire _02354_;
 wire _02355_;
 wire _02356_;
 wire _02357_;
 wire _02358_;
 wire _02359_;
 wire _02360_;
 wire _02361_;
 wire _02362_;
 wire _02363_;
 wire _02364_;
 wire _02365_;
 wire _02366_;
 wire _02367_;
 wire _02368_;
 wire _02369_;
 wire _02370_;
 wire _02371_;
 wire _02372_;
 wire _02373_;
 wire _02374_;
 wire _02375_;
 wire _02376_;
 wire _02377_;
 wire _02378_;
 wire _02379_;
 wire _02380_;
 wire _02381_;
 wire _02382_;
 wire _02383_;
 wire _02384_;
 wire _02385_;
 wire _02386_;
 wire _02387_;
 wire _02388_;
 wire _02389_;
 wire _02390_;
 wire _02391_;
 wire _02392_;
 wire _02393_;
 wire _02394_;
 wire _02395_;
 wire _02396_;
 wire _02397_;
 wire _02398_;
 wire _02399_;
 wire _02400_;
 wire _02401_;
 wire _02402_;
 wire _02403_;
 wire _02404_;
 wire _02405_;
 wire _02406_;
 wire _02407_;
 wire _02408_;
 wire _02409_;
 wire _02410_;
 wire _02411_;
 wire _02412_;
 wire _02413_;
 wire _02414_;
 wire _02415_;
 wire _02416_;
 wire _02417_;
 wire _02418_;
 wire _02419_;
 wire _02420_;
 wire _02421_;
 wire _02422_;
 wire _02423_;
 wire _02424_;
 wire _02425_;
 wire _02426_;
 wire _02427_;
 wire _02428_;
 wire _02429_;
 wire _02430_;
 wire _02431_;
 wire _02432_;
 wire _02433_;
 wire _02434_;
 wire _02435_;
 wire _02436_;
 wire _02437_;
 wire _02438_;
 wire _02439_;
 wire _02440_;
 wire _02441_;
 wire _02442_;
 wire _02443_;
 wire _02444_;
 wire _02445_;
 wire _02446_;
 wire _02447_;
 wire _02448_;
 wire _02449_;
 wire _02450_;
 wire _02451_;
 wire _02452_;
 wire _02453_;
 wire _02454_;
 wire _02455_;
 wire _02456_;
 wire _02457_;
 wire _02458_;
 wire _02459_;
 wire _02460_;
 wire _02461_;
 wire _02462_;
 wire _02463_;
 wire _02464_;
 wire _02465_;
 wire _02466_;
 wire _02467_;
 wire _02468_;
 wire _02469_;
 wire _02470_;
 wire _02471_;
 wire _02472_;
 wire _02473_;
 wire _02474_;
 wire _02475_;
 wire _02476_;
 wire _02477_;
 wire _02478_;
 wire _02479_;
 wire _02480_;
 wire _02481_;
 wire _02482_;
 wire _02483_;
 wire _02484_;
 wire _02485_;
 wire _02486_;
 wire _02487_;
 wire _02488_;
 wire _02489_;
 wire _02490_;
 wire _02491_;
 wire _02492_;
 wire _02493_;
 wire _02494_;
 wire _02495_;
 wire _02496_;
 wire _02497_;
 wire _02498_;
 wire _02499_;
 wire _02500_;
 wire _02501_;
 wire _02502_;
 wire _02503_;
 wire _02504_;
 wire _02505_;
 wire _02506_;
 wire _02507_;
 wire _02508_;
 wire _02509_;
 wire _02510_;
 wire _02511_;
 wire _02512_;
 wire _02513_;
 wire _02514_;
 wire _02515_;
 wire _02516_;
 wire _02517_;
 wire _02518_;
 wire _02519_;
 wire _02520_;
 wire _02521_;
 wire _02522_;
 wire _02523_;
 wire _02524_;
 wire _02525_;
 wire _02526_;
 wire _02527_;
 wire _02528_;
 wire _02529_;
 wire _02530_;
 wire _02531_;
 wire _02532_;
 wire _02533_;
 wire _02534_;
 wire _02535_;
 wire _02536_;
 wire _02537_;
 wire _02538_;
 wire _02539_;
 wire _02540_;
 wire _02541_;
 wire _02542_;
 wire _02543_;
 wire _02544_;
 wire _02545_;
 wire _02546_;
 wire _02547_;
 wire _02548_;
 wire _02549_;
 wire _02550_;
 wire _02551_;
 wire _02552_;
 wire _02553_;
 wire _02554_;
 wire _02555_;
 wire _02556_;
 wire _02557_;
 wire _02558_;
 wire _02559_;
 wire _02560_;
 wire _02561_;
 wire _02562_;
 wire _02563_;
 wire _02564_;
 wire _02565_;
 wire _02566_;
 wire _02567_;
 wire _02568_;
 wire _02569_;
 wire _02570_;
 wire _02571_;
 wire _02572_;
 wire _02573_;
 wire _02574_;
 wire _02575_;
 wire _02576_;
 wire _02577_;
 wire _02578_;
 wire _02579_;
 wire _02580_;
 wire _02581_;
 wire _02582_;
 wire _02583_;
 wire _02584_;
 wire _02585_;
 wire _02586_;
 wire _02587_;
 wire _02588_;
 wire _02589_;
 wire _02590_;
 wire _02591_;
 wire _02592_;
 wire _02593_;
 wire _02594_;
 wire _02595_;
 wire _02596_;
 wire _02597_;
 wire _02598_;
 wire _02599_;
 wire _02600_;
 wire _02601_;
 wire _02602_;
 wire _02603_;
 wire _02604_;
 wire _02605_;
 wire _02606_;
 wire _02607_;
 wire _02608_;
 wire _02609_;
 wire _02610_;
 wire _02611_;
 wire _02612_;
 wire _02613_;
 wire _02614_;
 wire _02615_;
 wire _02616_;
 wire _02617_;
 wire _02618_;
 wire _02619_;
 wire _02620_;
 wire _02621_;
 wire _02622_;
 wire _02623_;
 wire _02624_;
 wire _02625_;
 wire _02626_;
 wire _02627_;
 wire _02628_;
 wire _02629_;
 wire _02630_;
 wire _02631_;
 wire _02632_;
 wire _02633_;
 wire _02634_;
 wire _02635_;
 wire _02636_;
 wire _02637_;
 wire _02638_;
 wire _02639_;
 wire _02640_;
 wire _02641_;
 wire _02642_;
 wire _02643_;
 wire _02644_;
 wire _02645_;
 wire _02646_;
 wire _02647_;
 wire _02648_;
 wire _02649_;
 wire _02650_;
 wire _02651_;
 wire _02652_;
 wire _02653_;
 wire _02654_;
 wire _02655_;
 wire _02656_;
 wire _02657_;
 wire _02658_;
 wire _02659_;
 wire _02660_;
 wire _02661_;
 wire _02662_;
 wire _02663_;
 wire _02664_;
 wire _02665_;
 wire _02666_;
 wire _02667_;
 wire _02668_;
 wire _02669_;
 wire _02670_;
 wire _02671_;
 wire _02672_;
 wire _02673_;
 wire _02674_;
 wire _02675_;
 wire _02676_;
 wire _02677_;
 wire _02678_;
 wire _02679_;
 wire _02680_;
 wire _02681_;
 wire _02682_;
 wire _02683_;
 wire _02684_;
 wire _02685_;
 wire _02686_;
 wire _02687_;
 wire _02688_;
 wire _02689_;
 wire _02690_;
 wire _02691_;
 wire _02692_;
 wire _02693_;
 wire _02694_;
 wire _02695_;
 wire _02696_;
 wire _02697_;
 wire _02698_;
 wire _02699_;
 wire _02700_;
 wire _02701_;
 wire _02702_;
 wire _02703_;
 wire _02704_;
 wire _02705_;
 wire _02706_;
 wire _02707_;
 wire _02708_;
 wire _02709_;
 wire _02710_;
 wire _02711_;
 wire _02712_;
 wire _02713_;
 wire _02714_;
 wire _02715_;
 wire _02716_;
 wire _02717_;
 wire _02718_;
 wire _02719_;
 wire _02720_;
 wire _02721_;
 wire _02722_;
 wire _02723_;
 wire _02724_;
 wire _02725_;
 wire _02726_;
 wire _02727_;
 wire _02728_;
 wire _02729_;
 wire _02730_;
 wire _02731_;
 wire _02732_;
 wire _02733_;
 wire _02734_;
 wire _02735_;
 wire _02736_;
 wire _02737_;
 wire _02738_;
 wire _02739_;
 wire _02740_;
 wire _02741_;
 wire _02742_;
 wire _02743_;
 wire _02744_;
 wire _02745_;
 wire _02746_;
 wire _02747_;
 wire _02748_;
 wire _02749_;
 wire _02750_;
 wire _02751_;
 wire _02752_;
 wire _02753_;
 wire _02754_;
 wire _02755_;
 wire _02756_;
 wire _02757_;
 wire _02758_;
 wire _02759_;
 wire _02760_;
 wire _02761_;
 wire _02762_;
 wire _02763_;
 wire _02764_;
 wire _02765_;
 wire _02766_;
 wire _02767_;
 wire _02768_;
 wire _02769_;
 wire _02770_;
 wire _02771_;
 wire _02772_;
 wire _02773_;
 wire _02774_;
 wire _02775_;
 wire _02776_;
 wire _02777_;
 wire _02778_;
 wire _02779_;
 wire _02780_;
 wire _02781_;
 wire _02782_;
 wire _02783_;
 wire _02784_;
 wire _02785_;
 wire _02786_;
 wire _02787_;
 wire _02788_;
 wire _02789_;
 wire _02790_;
 wire _02791_;
 wire _02792_;
 wire _02793_;
 wire _02794_;
 wire _02795_;
 wire _02796_;
 wire _02797_;
 wire _02798_;
 wire _02799_;
 wire _02800_;
 wire _02801_;
 wire _02802_;
 wire _02803_;
 wire _02804_;
 wire _02805_;
 wire _02806_;
 wire _02807_;
 wire _02808_;
 wire _02809_;
 wire _02810_;
 wire _02811_;
 wire _02812_;
 wire _02813_;
 wire _02814_;
 wire _02815_;
 wire _02816_;
 wire _02817_;
 wire _02818_;
 wire _02819_;
 wire _02820_;
 wire _02821_;
 wire _02822_;
 wire _02823_;
 wire _02824_;
 wire _02825_;
 wire _02826_;
 wire _02827_;
 wire _02828_;
 wire _02829_;
 wire _02830_;
 wire _02831_;
 wire _02832_;
 wire _02833_;
 wire _02834_;
 wire _02835_;
 wire _02836_;
 wire _02837_;
 wire _02838_;
 wire _02839_;
 wire _02840_;
 wire _02841_;
 wire _02842_;
 wire _02843_;
 wire _02844_;
 wire _02845_;
 wire _02846_;
 wire _02847_;
 wire _02848_;
 wire _02849_;
 wire _02850_;
 wire _02851_;
 wire _02852_;
 wire _02853_;
 wire _02854_;
 wire _02855_;
 wire _02856_;
 wire _02857_;
 wire _02858_;
 wire _02859_;
 wire _02860_;
 wire _02861_;
 wire _02862_;
 wire _02863_;
 wire _02864_;
 wire _02865_;
 wire _02866_;
 wire _02867_;
 wire _02868_;
 wire _02869_;
 wire _02870_;
 wire _02871_;
 wire _02872_;
 wire _02873_;
 wire _02874_;
 wire _02875_;
 wire _02876_;
 wire _02877_;
 wire _02878_;
 wire _02879_;
 wire _02880_;
 wire _02881_;
 wire _02882_;
 wire _02883_;
 wire _02884_;
 wire _02885_;
 wire _02886_;
 wire _02887_;
 wire _02888_;
 wire _02889_;
 wire _02890_;
 wire _02891_;
 wire _02892_;
 wire _02893_;
 wire _02894_;
 wire _02895_;
 wire _02896_;
 wire _02897_;
 wire _02898_;
 wire _02899_;
 wire _02900_;
 wire _02901_;
 wire _02902_;
 wire _02903_;
 wire _02904_;
 wire _02905_;
 wire _02906_;
 wire _02907_;
 wire _02908_;
 wire _02909_;
 wire _02910_;
 wire _02911_;
 wire _02912_;
 wire _02913_;
 wire _02914_;
 wire _02915_;
 wire _02916_;
 wire _02917_;
 wire _02918_;
 wire _02919_;
 wire _02920_;
 wire _02921_;
 wire _02922_;
 wire _02923_;
 wire _02924_;
 wire _02925_;
 wire _02926_;
 wire _02927_;
 wire _02928_;
 wire _02929_;
 wire _02930_;
 wire _02931_;
 wire _02932_;
 wire _02933_;
 wire _02934_;
 wire _02935_;
 wire _02936_;
 wire _02937_;
 wire _02938_;
 wire _02939_;
 wire _02940_;
 wire _02941_;
 wire _02942_;
 wire _02943_;
 wire _02944_;
 wire _02945_;
 wire _02946_;
 wire _02947_;
 wire _02948_;
 wire _02949_;
 wire _02950_;
 wire _02951_;
 wire _02952_;
 wire _02953_;
 wire _02954_;
 wire _02955_;
 wire _02956_;
 wire _02957_;
 wire _02958_;
 wire _02959_;
 wire _02960_;
 wire _02961_;
 wire _02962_;
 wire _02963_;
 wire _02964_;
 wire _02965_;
 wire _02966_;
 wire _02967_;
 wire _02968_;
 wire _02969_;
 wire _02970_;
 wire _02971_;
 wire _02972_;
 wire _02973_;
 wire _02974_;
 wire _02975_;
 wire _02976_;
 wire _02977_;
 wire _02978_;
 wire _02979_;
 wire _02980_;
 wire _02981_;
 wire _02982_;
 wire _02983_;
 wire _02984_;
 wire _02985_;
 wire _02986_;
 wire _02987_;
 wire _02988_;
 wire _02989_;
 wire _02990_;
 wire _02991_;
 wire _02992_;
 wire _02993_;
 wire _02994_;
 wire _02995_;
 wire _02996_;
 wire _02997_;
 wire _02998_;
 wire _02999_;
 wire _03000_;
 wire _03001_;
 wire _03002_;
 wire _03003_;
 wire _03004_;
 wire _03005_;
 wire _03006_;
 wire _03007_;
 wire _03008_;
 wire _03009_;
 wire _03010_;
 wire _03011_;
 wire _03012_;
 wire _03013_;
 wire _03014_;
 wire _03015_;
 wire _03016_;
 wire _03017_;
 wire _03018_;
 wire _03019_;
 wire _03020_;
 wire _03021_;
 wire _03022_;
 wire _03023_;
 wire _03024_;
 wire _03025_;
 wire _03026_;
 wire _03027_;
 wire _03028_;
 wire _03029_;
 wire _03030_;
 wire _03031_;
 wire _03032_;
 wire _03033_;
 wire _03034_;
 wire _03035_;
 wire _03036_;
 wire _03037_;
 wire _03038_;
 wire _03039_;
 wire _03040_;
 wire _03041_;
 wire _03042_;
 wire _03043_;
 wire _03044_;
 wire _03045_;
 wire _03046_;
 wire _03047_;
 wire _03048_;
 wire _03049_;
 wire _03050_;
 wire _03051_;
 wire _03052_;
 wire _03053_;
 wire _03054_;
 wire _03055_;
 wire _03056_;
 wire _03057_;
 wire _03058_;
 wire _03059_;
 wire _03060_;
 wire _03061_;
 wire _03062_;
 wire _03063_;
 wire _03064_;
 wire _03065_;
 wire _03066_;
 wire _03067_;
 wire _03068_;
 wire _03069_;
 wire _03070_;
 wire _03071_;
 wire _03072_;
 wire _03073_;
 wire _03074_;
 wire _03075_;
 wire _03076_;
 wire _03077_;
 wire _03078_;
 wire _03079_;
 wire _03080_;
 wire _03081_;
 wire _03082_;
 wire _03083_;
 wire _03084_;
 wire _03085_;
 wire _03086_;
 wire _03087_;
 wire _03088_;
 wire _03089_;
 wire _03090_;
 wire _03091_;
 wire _03092_;
 wire _03093_;
 wire _03094_;
 wire _03095_;
 wire _03096_;
 wire _03097_;
 wire _03098_;
 wire _03099_;
 wire _03100_;
 wire _03101_;
 wire _03102_;
 wire _03103_;
 wire _03104_;
 wire _03105_;
 wire _03106_;
 wire _03107_;
 wire _03108_;
 wire _03109_;
 wire _03110_;
 wire _03111_;
 wire _03112_;
 wire _03113_;
 wire _03114_;
 wire _03115_;
 wire _03116_;
 wire _03117_;
 wire _03118_;
 wire _03119_;
 wire _03120_;
 wire _03121_;
 wire _03122_;
 wire _03123_;
 wire _03124_;
 wire _03125_;
 wire _03126_;
 wire _03127_;
 wire _03128_;
 wire _03129_;
 wire _03130_;
 wire _03131_;
 wire _03132_;
 wire _03133_;
 wire _03134_;
 wire _03135_;
 wire _03136_;
 wire _03137_;
 wire _03138_;
 wire _03139_;
 wire _03140_;
 wire _03141_;
 wire _03142_;
 wire _03143_;
 wire _03144_;
 wire _03145_;
 wire _03146_;
 wire _03147_;
 wire _03148_;
 wire _03149_;
 wire _03150_;
 wire _03151_;
 wire _03152_;
 wire _03153_;
 wire _03154_;
 wire _03155_;
 wire _03156_;
 wire _03157_;
 wire _03158_;
 wire _03159_;
 wire _03160_;
 wire _03161_;
 wire _03162_;
 wire _03163_;
 wire _03164_;
 wire _03165_;
 wire _03166_;
 wire _03167_;
 wire _03168_;
 wire _03169_;
 wire _03170_;
 wire _03171_;
 wire _03172_;
 wire _03173_;
 wire _03174_;
 wire _03175_;
 wire _03176_;
 wire _03177_;
 wire _03178_;
 wire _03179_;
 wire _03180_;
 wire _03181_;
 wire _03182_;
 wire _03183_;
 wire _03184_;
 wire _03185_;
 wire _03186_;
 wire _03187_;
 wire _03188_;
 wire _03189_;
 wire _03190_;
 wire _03191_;
 wire _03192_;
 wire _03193_;
 wire _03194_;
 wire _03195_;
 wire _03196_;
 wire _03197_;
 wire _03198_;
 wire _03199_;
 wire _03200_;
 wire _03201_;
 wire _03202_;
 wire _03203_;
 wire _03204_;
 wire _03205_;
 wire _03206_;
 wire _03207_;
 wire _03208_;
 wire _03209_;
 wire _03210_;
 wire _03211_;
 wire _03212_;
 wire _03213_;
 wire _03214_;
 wire _03215_;
 wire _03216_;
 wire _03217_;
 wire _03218_;
 wire _03219_;
 wire _03220_;
 wire _03221_;
 wire _03222_;
 wire _03223_;
 wire _03224_;
 wire _03225_;
 wire _03226_;
 wire _03227_;
 wire _03228_;
 wire _03229_;
 wire _03230_;
 wire _03231_;
 wire _03232_;
 wire _03233_;
 wire _03234_;
 wire _03235_;
 wire _03236_;
 wire _03237_;
 wire _03238_;
 wire _03239_;
 wire _03240_;
 wire _03241_;
 wire _03242_;
 wire _03243_;
 wire _03244_;
 wire _03245_;
 wire _03246_;
 wire _03247_;
 wire _03248_;
 wire _03249_;
 wire _03250_;
 wire _03251_;
 wire _03252_;
 wire _03253_;
 wire _03254_;
 wire _03255_;
 wire _03256_;
 wire _03257_;
 wire _03258_;
 wire _03259_;
 wire _03260_;
 wire _03261_;
 wire _03262_;
 wire _03263_;
 wire _03264_;
 wire _03265_;
 wire _03266_;
 wire _03267_;
 wire _03268_;
 wire _03269_;
 wire _03270_;
 wire _03271_;
 wire _03272_;
 wire _03273_;
 wire _03274_;
 wire _03275_;
 wire _03276_;
 wire _03277_;
 wire _03278_;
 wire _03279_;
 wire _03280_;
 wire _03281_;
 wire _03282_;
 wire _03283_;
 wire _03284_;
 wire _03285_;
 wire _03286_;
 wire _03287_;
 wire _03288_;
 wire _03289_;
 wire _03290_;
 wire _03291_;
 wire _03292_;
 wire _03293_;
 wire _03294_;
 wire _03295_;
 wire _03296_;
 wire _03297_;
 wire _03298_;
 wire _03299_;
 wire _03300_;
 wire _03301_;
 wire _03302_;
 wire _03303_;
 wire _03304_;
 wire _03305_;
 wire _03306_;
 wire _03307_;
 wire _03308_;
 wire _03309_;
 wire _03310_;
 wire _03311_;
 wire _03312_;
 wire _03313_;
 wire _03314_;
 wire _03315_;
 wire _03316_;
 wire _03317_;
 wire _03318_;
 wire _03319_;
 wire _03320_;
 wire _03321_;
 wire _03322_;
 wire _03323_;
 wire _03324_;
 wire _03325_;
 wire _03326_;
 wire _03327_;
 wire _03328_;
 wire _03329_;
 wire _03330_;
 wire _03331_;
 wire _03332_;
 wire _03333_;
 wire _03334_;
 wire _03335_;
 wire _03336_;
 wire _03337_;
 wire _03338_;
 wire _03339_;
 wire _03340_;
 wire _03341_;
 wire _03342_;
 wire _03343_;
 wire _03344_;
 wire _03345_;
 wire _03346_;
 wire _03347_;
 wire _03348_;
 wire _03349_;
 wire _03350_;
 wire _03351_;
 wire _03352_;
 wire _03353_;
 wire _03354_;
 wire _03355_;
 wire _03356_;
 wire _03357_;
 wire _03358_;
 wire _03359_;
 wire _03360_;
 wire _03361_;
 wire _03362_;
 wire _03363_;
 wire _03364_;
 wire _03365_;
 wire _03366_;
 wire _03367_;
 wire _03368_;
 wire _03369_;
 wire _03370_;
 wire _03371_;
 wire _03372_;
 wire _03373_;
 wire _03374_;
 wire _03375_;
 wire _03376_;
 wire _03377_;
 wire _03378_;
 wire _03379_;
 wire _03380_;
 wire _03381_;
 wire _03382_;
 wire _03383_;
 wire _03384_;
 wire _03385_;
 wire _03386_;
 wire _03387_;
 wire _03388_;
 wire _03389_;
 wire _03390_;
 wire _03391_;
 wire _03392_;
 wire _03393_;
 wire _03394_;
 wire _03395_;
 wire _03396_;
 wire _03397_;
 wire _03398_;
 wire _03399_;
 wire _03400_;
 wire _03401_;
 wire _03402_;
 wire _03403_;
 wire _03404_;
 wire _03405_;
 wire _03406_;
 wire _03407_;
 wire _03408_;
 wire _03409_;
 wire _03410_;
 wire _03411_;
 wire _03412_;
 wire _03413_;
 wire _03414_;
 wire _03415_;
 wire _03416_;
 wire _03417_;
 wire _03418_;
 wire _03419_;
 wire _03420_;
 wire _03421_;
 wire _03422_;
 wire _03423_;
 wire _03424_;
 wire _03425_;
 wire _03426_;
 wire _03427_;
 wire _03428_;
 wire _03429_;
 wire _03430_;
 wire _03431_;
 wire _03432_;
 wire _03433_;
 wire _03434_;
 wire _03435_;
 wire _03436_;
 wire _03437_;
 wire _03438_;
 wire _03439_;
 wire _03440_;
 wire _03441_;
 wire _03442_;
 wire _03443_;
 wire _03444_;
 wire _03445_;
 wire _03446_;
 wire _03447_;
 wire _03448_;
 wire _03449_;
 wire _03450_;
 wire _03451_;
 wire _03452_;
 wire _03453_;
 wire _03454_;
 wire _03455_;
 wire _03456_;
 wire _03457_;
 wire _03458_;
 wire _03459_;
 wire _03460_;
 wire _03461_;
 wire _03462_;
 wire _03463_;
 wire _03464_;
 wire _03465_;
 wire _03466_;
 wire _03467_;
 wire _03468_;
 wire _03469_;
 wire _03470_;
 wire _03471_;
 wire _03472_;
 wire _03473_;
 wire _03474_;
 wire _03475_;
 wire _03476_;
 wire _03477_;
 wire _03478_;
 wire _03479_;
 wire _03480_;
 wire _03481_;
 wire _03482_;
 wire _03483_;
 wire _03484_;
 wire _03485_;
 wire _03486_;
 wire _03487_;
 wire _03488_;
 wire _03489_;
 wire _03490_;
 wire _03491_;
 wire _03492_;
 wire _03493_;
 wire _03494_;
 wire _03495_;
 wire _03496_;
 wire _03497_;
 wire _03498_;
 wire _03499_;
 wire _03500_;
 wire _03501_;
 wire _03502_;
 wire _03503_;
 wire _03504_;
 wire _03505_;
 wire _03506_;
 wire _03507_;
 wire _03508_;
 wire _03509_;
 wire _03510_;
 wire _03511_;
 wire _03512_;
 wire _03513_;
 wire _03514_;
 wire _03515_;
 wire _03516_;
 wire _03517_;
 wire _03518_;
 wire _03519_;
 wire _03520_;
 wire _03521_;
 wire _03522_;
 wire _03523_;
 wire _03524_;
 wire _03525_;
 wire _03526_;
 wire _03527_;
 wire _03528_;
 wire _03529_;
 wire _03530_;
 wire _03531_;
 wire _03532_;
 wire _03533_;
 wire _03534_;
 wire _03535_;
 wire _03536_;
 wire _03537_;
 wire _03538_;
 wire _03539_;
 wire _03540_;
 wire _03541_;
 wire _03542_;
 wire _03543_;
 wire _03544_;
 wire _03545_;
 wire _03546_;
 wire _03547_;
 wire _03548_;
 wire _03549_;
 wire _03550_;
 wire _03551_;
 wire _03552_;
 wire _03553_;
 wire _03554_;
 wire _03555_;
 wire _03556_;
 wire _03557_;
 wire _03558_;
 wire _03559_;
 wire _03560_;
 wire _03561_;
 wire _03562_;
 wire _03563_;
 wire _03564_;
 wire _03565_;
 wire _03566_;
 wire _03567_;
 wire _03568_;
 wire _03569_;
 wire _03570_;
 wire _03571_;
 wire _03572_;
 wire _03573_;
 wire _03574_;
 wire _03575_;
 wire _03576_;
 wire _03577_;
 wire _03578_;
 wire _03579_;
 wire _03580_;
 wire _03581_;
 wire _03582_;
 wire _03583_;
 wire _03584_;
 wire _03585_;
 wire _03586_;
 wire _03587_;
 wire _03588_;
 wire _03589_;
 wire _03590_;
 wire _03591_;
 wire _03592_;
 wire _03593_;
 wire _03594_;
 wire _03595_;
 wire _03596_;
 wire _03597_;
 wire _03598_;
 wire _03599_;
 wire _03600_;
 wire _03601_;
 wire _03602_;
 wire _03603_;
 wire _03604_;
 wire _03605_;
 wire _03606_;
 wire _03607_;
 wire _03608_;
 wire _03609_;
 wire _03610_;
 wire _03611_;
 wire _03612_;
 wire _03613_;
 wire _03614_;
 wire _03615_;
 wire _03616_;
 wire _03617_;
 wire _03618_;
 wire _03619_;
 wire _03620_;
 wire _03621_;
 wire _03622_;
 wire _03623_;
 wire _03624_;
 wire _03625_;
 wire _03626_;
 wire _03627_;
 wire _03628_;
 wire _03629_;
 wire _03630_;
 wire _03631_;
 wire _03632_;
 wire _03633_;
 wire _03634_;
 wire _03635_;
 wire _03636_;
 wire _03637_;
 wire _03638_;
 wire _03639_;
 wire _03640_;
 wire _03641_;
 wire _03642_;
 wire _03643_;
 wire _03644_;
 wire _03645_;
 wire _03646_;
 wire _03647_;
 wire _03648_;
 wire _03649_;
 wire _03650_;
 wire _03651_;
 wire _03652_;
 wire _03653_;
 wire _03654_;
 wire _03655_;
 wire _03656_;
 wire _03657_;
 wire _03658_;
 wire _03659_;
 wire _03660_;
 wire _03661_;
 wire _03662_;
 wire _03663_;
 wire _03664_;
 wire _03665_;
 wire _03666_;
 wire _03667_;
 wire _03668_;
 wire _03669_;
 wire _03670_;
 wire _03671_;
 wire _03672_;
 wire _03673_;
 wire _03674_;
 wire _03675_;
 wire _03676_;
 wire _03677_;
 wire _03678_;
 wire _03679_;
 wire _03680_;
 wire _03681_;
 wire _03682_;
 wire _03683_;
 wire _03684_;
 wire _03685_;
 wire _03686_;
 wire _03687_;
 wire _03688_;
 wire _03689_;
 wire _03690_;
 wire _03691_;
 wire _03692_;
 wire _03693_;
 wire _03694_;
 wire _03695_;
 wire _03696_;
 wire _03697_;
 wire _03698_;
 wire _03699_;
 wire _03700_;
 wire _03701_;
 wire _03702_;
 wire _03703_;
 wire _03704_;
 wire _03705_;
 wire _03706_;
 wire _03707_;
 wire _03708_;
 wire _03709_;
 wire _03710_;
 wire _03711_;
 wire _03712_;
 wire _03713_;
 wire _03714_;
 wire _03715_;
 wire _03716_;
 wire _03717_;
 wire _03718_;
 wire _03719_;
 wire _03720_;
 wire _03721_;
 wire _03722_;
 wire _03723_;
 wire _03724_;
 wire _03725_;
 wire _03726_;
 wire _03727_;
 wire _03728_;
 wire _03729_;
 wire _03730_;
 wire _03731_;
 wire _03732_;
 wire _03733_;
 wire _03734_;
 wire _03735_;
 wire _03736_;
 wire _03737_;
 wire _03738_;
 wire _03739_;
 wire _03740_;
 wire _03741_;
 wire _03742_;
 wire _03743_;
 wire _03744_;
 wire _03745_;
 wire _03746_;
 wire _03747_;
 wire _03748_;
 wire _03749_;
 wire _03750_;
 wire _03751_;
 wire _03752_;
 wire _03753_;
 wire _03754_;
 wire _03755_;
 wire _03756_;
 wire _03757_;
 wire _03758_;
 wire _03759_;
 wire _03760_;
 wire _03761_;
 wire _03762_;
 wire _03763_;
 wire _03764_;
 wire _03765_;
 wire _03766_;
 wire _03767_;
 wire _03768_;
 wire _03769_;
 wire _03770_;
 wire _03771_;
 wire _03772_;
 wire _03773_;
 wire _03774_;
 wire _03775_;
 wire _03776_;
 wire _03777_;
 wire _03778_;
 wire _03779_;
 wire _03780_;
 wire _03781_;
 wire _03782_;
 wire _03783_;
 wire _03784_;
 wire _03785_;
 wire _03786_;
 wire _03787_;
 wire _03788_;
 wire _03789_;
 wire _03790_;
 wire _03791_;
 wire _03792_;
 wire _03793_;
 wire _03794_;
 wire _03795_;
 wire _03796_;
 wire _03797_;
 wire _03798_;
 wire _03799_;
 wire _03800_;
 wire _03801_;
 wire _03802_;
 wire _03803_;
 wire _03804_;
 wire _03805_;
 wire _03806_;
 wire _03807_;
 wire _03808_;
 wire _03809_;
 wire _03810_;
 wire _03811_;
 wire _03812_;
 wire _03813_;
 wire _03814_;
 wire _03815_;
 wire _03816_;
 wire _03817_;
 wire _03818_;
 wire _03819_;
 wire _03820_;
 wire _03821_;
 wire _03822_;
 wire _03823_;
 wire _03824_;
 wire _03825_;
 wire _03826_;
 wire _03827_;
 wire _03828_;
 wire _03829_;
 wire _03830_;
 wire _03831_;
 wire _03832_;
 wire _03833_;
 wire _03834_;
 wire _03835_;
 wire _03836_;
 wire _03837_;
 wire _03838_;
 wire _03839_;
 wire _03840_;
 wire _03841_;
 wire _03842_;
 wire _03843_;
 wire _03844_;
 wire _03845_;
 wire _03846_;
 wire _03847_;
 wire _03848_;
 wire _03849_;
 wire _03850_;
 wire _03851_;
 wire _03852_;
 wire _03853_;
 wire _03854_;
 wire _03855_;
 wire _03856_;
 wire _03857_;
 wire _03858_;
 wire _03859_;
 wire _03860_;
 wire _03861_;
 wire _03862_;
 wire _03863_;
 wire _03864_;
 wire _03865_;
 wire _03866_;
 wire _03867_;
 wire _03868_;
 wire _03869_;
 wire _03870_;
 wire _03871_;
 wire _03872_;
 wire _03873_;
 wire _03874_;
 wire _03875_;
 wire _03876_;
 wire _03877_;
 wire _03878_;
 wire _03879_;
 wire _03880_;
 wire _03881_;
 wire _03882_;
 wire _03883_;
 wire _03884_;
 wire _03885_;
 wire _03886_;
 wire _03887_;
 wire _03888_;
 wire _03889_;
 wire _03890_;
 wire _03891_;
 wire _03892_;
 wire _03893_;
 wire _03894_;
 wire _03895_;
 wire _03896_;
 wire _03897_;
 wire _03898_;
 wire _03899_;
 wire _03900_;
 wire _03901_;
 wire _03902_;
 wire _03903_;
 wire _03904_;
 wire _03905_;
 wire _03906_;
 wire _03907_;
 wire _03908_;
 wire _03909_;
 wire _03910_;
 wire _03911_;
 wire _03912_;
 wire _03913_;
 wire _03914_;
 wire _03915_;
 wire _03916_;
 wire _03917_;
 wire _03918_;
 wire _03919_;
 wire _03920_;
 wire _03921_;
 wire _03922_;
 wire _03923_;
 wire _03924_;
 wire _03925_;
 wire _03926_;
 wire _03927_;
 wire _03928_;
 wire _03929_;
 wire _03930_;
 wire _03931_;
 wire _03932_;
 wire _03933_;
 wire _03934_;
 wire _03935_;
 wire _03936_;
 wire _03937_;
 wire _03938_;
 wire _03939_;
 wire _03940_;
 wire _03941_;
 wire _03942_;
 wire _03943_;
 wire _03944_;
 wire _03945_;
 wire _03946_;
 wire _03947_;
 wire _03948_;
 wire _03949_;
 wire _03950_;
 wire _03951_;
 wire _03952_;
 wire _03953_;
 wire _03954_;
 wire _03955_;
 wire _03956_;
 wire _03957_;
 wire _03958_;
 wire _03959_;
 wire _03960_;
 wire _03961_;
 wire _03962_;
 wire _03963_;
 wire _03964_;
 wire _03965_;
 wire _03966_;
 wire _03967_;
 wire _03968_;
 wire _03969_;
 wire _03970_;
 wire _03971_;
 wire _03972_;
 wire _03973_;
 wire _03974_;
 wire _03975_;
 wire _03976_;
 wire _03977_;
 wire _03978_;
 wire _03979_;
 wire _03980_;
 wire _03981_;
 wire _03982_;
 wire _03983_;
 wire _03984_;
 wire _03985_;
 wire _03986_;
 wire _03987_;
 wire _03988_;
 wire _03989_;
 wire _03990_;
 wire _03991_;
 wire _03992_;
 wire _03993_;
 wire _03994_;
 wire _03995_;
 wire _03996_;
 wire _03997_;
 wire _03998_;
 wire _03999_;
 wire _04000_;
 wire _04001_;
 wire _04002_;
 wire _04003_;
 wire _04004_;
 wire _04005_;
 wire _04006_;
 wire _04007_;
 wire _04008_;
 wire _04009_;
 wire _04010_;
 wire _04011_;
 wire _04012_;
 wire _04013_;
 wire _04014_;
 wire _04015_;
 wire _04016_;
 wire _04017_;
 wire _04018_;
 wire _04019_;
 wire _04020_;
 wire _04021_;
 wire _04022_;
 wire _04023_;
 wire _04024_;
 wire _04025_;
 wire _04026_;
 wire _04027_;
 wire _04028_;
 wire _04029_;
 wire _04030_;
 wire _04031_;
 wire _04032_;
 wire _04033_;
 wire _04034_;
 wire _04035_;
 wire _04036_;
 wire _04037_;
 wire _04038_;
 wire _04039_;
 wire _04040_;
 wire _04041_;
 wire _04042_;
 wire _04043_;
 wire _04044_;
 wire _04045_;
 wire _04046_;
 wire _04047_;
 wire _04048_;
 wire _04049_;
 wire _04050_;
 wire _04051_;
 wire _04052_;
 wire _04053_;
 wire _04054_;
 wire _04055_;
 wire _04056_;
 wire _04057_;
 wire _04058_;
 wire _04059_;
 wire _04060_;
 wire _04061_;
 wire _04062_;
 wire _04063_;
 wire _04064_;
 wire _04065_;
 wire _04066_;
 wire _04067_;
 wire _04068_;
 wire _04069_;
 wire _04070_;
 wire _04071_;
 wire _04072_;
 wire _04073_;
 wire _04074_;
 wire _04075_;
 wire _04076_;
 wire _04077_;
 wire _04078_;
 wire _04079_;
 wire _04080_;
 wire _04081_;
 wire _04082_;
 wire _04083_;
 wire _04084_;
 wire _04085_;
 wire _04086_;
 wire _04087_;
 wire _04088_;
 wire _04089_;
 wire _04090_;
 wire _04091_;
 wire _04092_;
 wire _04093_;
 wire _04094_;
 wire _04095_;
 wire _04096_;
 wire _04097_;
 wire _04098_;
 wire _04099_;
 wire _04100_;
 wire _04101_;
 wire _04102_;
 wire _04103_;
 wire _04104_;
 wire _04105_;
 wire _04106_;
 wire _04107_;
 wire _04108_;
 wire _04109_;
 wire _04110_;
 wire _04111_;
 wire _04112_;
 wire _04113_;
 wire _04114_;
 wire _04115_;
 wire _04116_;
 wire _04117_;
 wire _04118_;
 wire _04119_;
 wire _04120_;
 wire _04121_;
 wire _04122_;
 wire _04123_;
 wire _04124_;
 wire _04125_;
 wire _04126_;
 wire _04127_;
 wire _04128_;
 wire _04129_;
 wire _04130_;
 wire _04131_;
 wire _04132_;
 wire _04133_;
 wire _04134_;
 wire _04135_;
 wire _04136_;
 wire _04137_;
 wire _04138_;
 wire _04139_;
 wire _04140_;
 wire _04141_;
 wire _04142_;
 wire _04143_;
 wire _04144_;
 wire _04145_;
 wire _04146_;
 wire _04147_;
 wire _04148_;
 wire _04149_;
 wire _04150_;
 wire _04151_;
 wire _04152_;
 wire _04153_;
 wire _04154_;
 wire _04155_;
 wire _04156_;
 wire _04157_;
 wire _04158_;
 wire _04159_;
 wire _04160_;
 wire _04161_;
 wire _04162_;
 wire _04163_;
 wire _04164_;
 wire _04165_;
 wire _04166_;
 wire _04167_;
 wire _04168_;
 wire _04169_;
 wire _04170_;
 wire _04171_;
 wire _04172_;
 wire _04173_;
 wire _04174_;
 wire _04175_;
 wire _04176_;
 wire _04177_;
 wire _04178_;
 wire _04179_;
 wire _04180_;
 wire _04181_;
 wire _04182_;
 wire _04183_;
 wire _04184_;
 wire _04185_;
 wire _04186_;
 wire _04187_;
 wire _04188_;
 wire _04189_;
 wire _04190_;
 wire _04191_;
 wire _04192_;
 wire _04193_;
 wire _04194_;
 wire _04195_;
 wire _04196_;
 wire _04197_;
 wire _04198_;
 wire _04199_;
 wire _04200_;
 wire _04201_;
 wire _04202_;
 wire _04203_;
 wire _04204_;
 wire _04205_;
 wire _04206_;
 wire _04207_;
 wire _04208_;
 wire _04209_;
 wire _04210_;
 wire _04211_;
 wire _04212_;
 wire _04213_;
 wire _04214_;
 wire _04215_;
 wire _04216_;
 wire _04217_;
 wire _04218_;
 wire _04219_;
 wire _04220_;
 wire _04221_;
 wire _04222_;
 wire _04223_;
 wire _04224_;
 wire _04225_;
 wire _04226_;
 wire _04227_;
 wire _04228_;
 wire _04229_;
 wire _04230_;
 wire _04231_;
 wire _04232_;
 wire _04233_;
 wire _04234_;
 wire _04235_;
 wire _04236_;
 wire _04237_;
 wire _04238_;
 wire _04239_;
 wire _04240_;
 wire _04241_;
 wire _04242_;
 wire _04243_;
 wire _04244_;
 wire _04245_;
 wire _04246_;
 wire _04247_;
 wire _04248_;
 wire _04249_;
 wire _04250_;
 wire _04251_;
 wire _04252_;
 wire _04253_;
 wire _04254_;
 wire _04255_;
 wire _04256_;
 wire _04257_;
 wire _04258_;
 wire _04259_;
 wire _04260_;
 wire _04261_;
 wire _04262_;
 wire _04263_;
 wire _04264_;
 wire _04265_;
 wire _04266_;
 wire _04267_;
 wire _04268_;
 wire _04269_;
 wire _04270_;
 wire _04271_;
 wire _04272_;
 wire _04273_;
 wire _04274_;
 wire _04275_;
 wire _04276_;
 wire _04277_;
 wire _04278_;
 wire _04279_;
 wire _04280_;
 wire _04281_;
 wire _04282_;
 wire _04283_;
 wire _04284_;
 wire _04285_;
 wire _04286_;
 wire _04287_;
 wire _04288_;
 wire _04289_;
 wire _04290_;
 wire _04291_;
 wire _04292_;
 wire _04293_;
 wire _04294_;
 wire _04295_;
 wire _04296_;
 wire _04297_;
 wire _04298_;
 wire _04299_;
 wire _04300_;
 wire _04301_;
 wire _04302_;
 wire _04303_;
 wire _04304_;
 wire _04305_;
 wire _04306_;
 wire _04307_;
 wire _04308_;
 wire _04309_;
 wire _04310_;
 wire _04311_;
 wire _04312_;
 wire _04313_;
 wire _04314_;
 wire _04315_;
 wire _04316_;
 wire _04317_;
 wire _04318_;
 wire _04319_;
 wire _04320_;
 wire _04321_;
 wire _04322_;
 wire _04323_;
 wire _04324_;
 wire _04325_;
 wire _04326_;
 wire _04327_;
 wire _04328_;
 wire _04329_;
 wire _04330_;
 wire _04331_;
 wire _04332_;
 wire _04333_;
 wire _04334_;
 wire _04335_;
 wire _04336_;
 wire _04337_;
 wire _04338_;
 wire _04339_;
 wire _04340_;
 wire _04341_;
 wire _04342_;
 wire _04343_;
 wire _04344_;
 wire _04345_;
 wire _04346_;
 wire _04347_;
 wire _04348_;
 wire _04349_;
 wire _04350_;
 wire _04351_;
 wire _04352_;
 wire _04353_;
 wire _04354_;
 wire _04355_;
 wire _04356_;
 wire _04357_;
 wire _04358_;
 wire _04359_;
 wire _04360_;
 wire _04361_;
 wire _04362_;
 wire _04363_;
 wire _04364_;
 wire _04365_;
 wire _04366_;
 wire _04367_;
 wire _04368_;
 wire _04369_;
 wire _04370_;
 wire _04371_;
 wire _04372_;
 wire _04373_;
 wire _04374_;
 wire _04375_;
 wire _04376_;
 wire _04377_;
 wire _04378_;
 wire _04379_;
 wire _04380_;
 wire _04381_;
 wire _04382_;
 wire _04383_;
 wire _04384_;
 wire _04385_;
 wire _04386_;
 wire _04387_;
 wire _04388_;
 wire _04389_;
 wire _04390_;
 wire _04391_;
 wire _04392_;
 wire _04393_;
 wire _04394_;
 wire _04395_;
 wire _04396_;
 wire _04397_;
 wire _04398_;
 wire _04399_;
 wire _04400_;
 wire _04401_;
 wire _04402_;
 wire _04403_;
 wire _04404_;
 wire _04405_;
 wire _04406_;
 wire _04407_;
 wire _04408_;
 wire _04409_;
 wire _04410_;
 wire _04411_;
 wire _04412_;
 wire _04413_;
 wire _04414_;
 wire _04415_;
 wire _04416_;
 wire _04417_;
 wire _04418_;
 wire _04419_;
 wire _04420_;
 wire _04421_;
 wire _04422_;
 wire _04423_;
 wire _04424_;
 wire _04425_;
 wire _04426_;
 wire _04427_;
 wire _04428_;
 wire _04429_;
 wire _04430_;
 wire _04431_;
 wire _04432_;
 wire _04433_;
 wire _04434_;
 wire _04435_;
 wire _04436_;
 wire _04437_;
 wire _04438_;
 wire _04439_;
 wire _04440_;
 wire _04441_;
 wire _04442_;
 wire _04443_;
 wire _04444_;
 wire _04445_;
 wire _04446_;
 wire _04447_;
 wire _04448_;
 wire _04449_;
 wire _04450_;
 wire _04451_;
 wire _04452_;
 wire _04453_;
 wire _04454_;
 wire _04455_;
 wire _04456_;
 wire _04457_;
 wire _04458_;
 wire _04459_;
 wire _04460_;
 wire _04461_;
 wire _04462_;
 wire _04463_;
 wire _04464_;
 wire _04465_;
 wire _04466_;
 wire _04467_;
 wire _04468_;
 wire _04469_;
 wire _04470_;
 wire _04471_;
 wire _04472_;
 wire _04473_;
 wire _04474_;
 wire _04475_;
 wire _04476_;
 wire _04477_;
 wire _04478_;
 wire _04479_;
 wire _04480_;
 wire _04481_;
 wire _04482_;
 wire _04483_;
 wire _04484_;
 wire _04485_;
 wire _04486_;
 wire _04487_;
 wire _04488_;
 wire _04489_;
 wire _04490_;
 wire _04491_;
 wire _04492_;
 wire _04493_;
 wire _04494_;
 wire _04495_;
 wire _04496_;
 wire _04497_;
 wire _04498_;
 wire _04499_;
 wire _04500_;
 wire _04501_;
 wire _04502_;
 wire _04503_;
 wire _04504_;
 wire _04505_;
 wire _04506_;
 wire _04507_;
 wire _04508_;
 wire _04509_;
 wire _04510_;
 wire _04511_;
 wire _04512_;
 wire _04513_;
 wire _04514_;
 wire _04515_;
 wire _04516_;
 wire _04517_;
 wire _04518_;
 wire _04519_;
 wire _04520_;
 wire _04521_;
 wire _04522_;
 wire _04523_;
 wire _04524_;
 wire _04525_;
 wire _04526_;
 wire _04527_;
 wire _04528_;
 wire _04529_;
 wire _04530_;
 wire _04531_;
 wire _04532_;
 wire _04533_;
 wire _04534_;
 wire _04535_;
 wire _04536_;
 wire _04537_;
 wire _04538_;
 wire _04539_;
 wire _04540_;
 wire _04541_;
 wire _04542_;
 wire _04543_;
 wire _04544_;
 wire _04545_;
 wire _04546_;
 wire _04547_;
 wire _04548_;
 wire _04549_;
 wire _04550_;
 wire _04551_;
 wire _04552_;
 wire _04553_;
 wire _04554_;
 wire _04555_;
 wire _04556_;
 wire _04557_;
 wire _04558_;
 wire _04559_;
 wire _04560_;
 wire _04561_;
 wire _04562_;
 wire _04563_;
 wire _04564_;
 wire _04565_;
 wire _04566_;
 wire _04567_;
 wire _04568_;
 wire _04569_;
 wire _04570_;
 wire _04571_;
 wire _04572_;
 wire _04573_;
 wire _04574_;
 wire _04575_;
 wire _04576_;
 wire _04577_;
 wire _04578_;
 wire _04579_;
 wire _04580_;
 wire _04581_;
 wire _04582_;
 wire _04583_;
 wire _04584_;
 wire _04585_;
 wire _04586_;
 wire _04587_;
 wire _04588_;
 wire _04589_;
 wire _04590_;
 wire _04591_;
 wire _04592_;
 wire _04593_;
 wire _04594_;
 wire _04595_;
 wire _04596_;
 wire _04597_;
 wire _04598_;
 wire _04599_;
 wire _04600_;
 wire _04601_;
 wire _04602_;
 wire _04603_;
 wire _04604_;
 wire _04605_;
 wire _04606_;
 wire _04607_;
 wire _04608_;
 wire _04609_;
 wire _04610_;
 wire _04611_;
 wire _04612_;
 wire _04613_;
 wire _04614_;
 wire _04615_;
 wire _04616_;
 wire _04617_;
 wire _04618_;
 wire _04619_;
 wire _04620_;
 wire _04621_;
 wire _04622_;
 wire _04623_;
 wire _04624_;
 wire _04625_;
 wire _04626_;
 wire _04627_;
 wire _04628_;
 wire _04629_;
 wire _04630_;
 wire _04631_;
 wire _04632_;
 wire _04633_;
 wire _04634_;
 wire _04635_;
 wire _04636_;
 wire _04637_;
 wire _04638_;
 wire _04639_;
 wire _04640_;
 wire _04641_;
 wire _04642_;
 wire _04643_;
 wire _04644_;
 wire _04645_;
 wire _04646_;
 wire _04647_;
 wire _04648_;
 wire _04649_;
 wire _04650_;
 wire _04651_;
 wire _04652_;
 wire _04653_;
 wire _04654_;
 wire _04655_;
 wire _04656_;
 wire _04657_;
 wire _04658_;
 wire _04659_;
 wire _04660_;
 wire _04661_;
 wire _04662_;
 wire _04663_;
 wire _04664_;
 wire _04665_;
 wire _04666_;
 wire _04667_;
 wire _04668_;
 wire _04669_;
 wire _04670_;
 wire _04671_;
 wire _04672_;
 wire _04673_;
 wire _04674_;
 wire _04675_;
 wire _04676_;
 wire _04677_;
 wire _04678_;
 wire _04679_;
 wire _04680_;
 wire _04681_;
 wire _04682_;
 wire _04683_;
 wire _04684_;
 wire _04685_;
 wire _04686_;
 wire _04687_;
 wire _04688_;
 wire _04689_;
 wire _04690_;
 wire _04691_;
 wire _04692_;
 wire _04693_;
 wire _04694_;
 wire _04695_;
 wire _04696_;
 wire _04697_;
 wire _04698_;
 wire _04699_;
 wire _04700_;
 wire _04701_;
 wire _04702_;
 wire _04703_;
 wire _04704_;
 wire _04705_;
 wire _04706_;
 wire _04707_;
 wire _04708_;
 wire _04709_;
 wire _04710_;
 wire _04711_;
 wire _04712_;
 wire _04713_;
 wire _04714_;
 wire _04715_;
 wire _04716_;
 wire _04717_;
 wire _04718_;
 wire _04719_;
 wire _04720_;
 wire _04721_;
 wire _04722_;
 wire _04723_;
 wire _04724_;
 wire _04725_;
 wire _04726_;
 wire _04727_;
 wire _04728_;
 wire _04729_;
 wire _04730_;
 wire _04731_;
 wire _04732_;
 wire _04733_;
 wire _04734_;
 wire _04735_;
 wire _04736_;
 wire _04737_;
 wire _04738_;
 wire _04739_;
 wire _04740_;
 wire _04741_;
 wire _04742_;
 wire _04743_;
 wire _04744_;
 wire _04745_;
 wire _04746_;
 wire _04747_;
 wire _04748_;
 wire _04749_;
 wire _04750_;
 wire _04751_;
 wire _04752_;
 wire _04753_;
 wire _04754_;
 wire _04755_;
 wire _04756_;
 wire _04757_;
 wire _04758_;
 wire _04759_;
 wire _04760_;
 wire _04761_;
 wire _04762_;
 wire _04763_;
 wire _04764_;
 wire _04765_;
 wire _04766_;
 wire _04767_;
 wire _04768_;
 wire _04769_;
 wire _04770_;
 wire _04771_;
 wire _04772_;
 wire _04773_;
 wire _04774_;
 wire _04775_;
 wire _04776_;
 wire _04777_;
 wire _04778_;
 wire _04779_;
 wire _04780_;
 wire _04781_;
 wire _04782_;
 wire _04783_;
 wire _04784_;
 wire _04785_;
 wire _04786_;
 wire _04787_;
 wire _04788_;
 wire _04789_;
 wire _04790_;
 wire _04791_;
 wire _04792_;
 wire _04793_;
 wire _04794_;
 wire _04795_;
 wire _04796_;
 wire _04797_;
 wire _04798_;
 wire _04799_;
 wire _04800_;
 wire _04801_;
 wire _04802_;
 wire _04803_;
 wire _04804_;
 wire _04805_;
 wire _04806_;
 wire _04807_;
 wire _04808_;
 wire _04809_;
 wire _04810_;
 wire _04811_;
 wire _04812_;
 wire _04813_;
 wire _04814_;
 wire _04815_;
 wire _04816_;
 wire _04817_;
 wire _04818_;
 wire _04819_;
 wire _04820_;
 wire _04821_;
 wire _04822_;
 wire _04823_;
 wire _04824_;
 wire _04825_;
 wire _04826_;
 wire _04827_;
 wire _04828_;
 wire _04829_;
 wire _04830_;
 wire _04831_;
 wire _04832_;
 wire _04833_;
 wire _04834_;
 wire _04835_;
 wire _04836_;
 wire _04837_;
 wire _04838_;
 wire _04839_;
 wire _04840_;
 wire _04841_;
 wire _04842_;
 wire _04843_;
 wire _04844_;
 wire _04845_;
 wire _04846_;
 wire _04847_;
 wire _04848_;
 wire _04849_;
 wire _04850_;
 wire _04851_;
 wire _04852_;
 wire _04853_;
 wire _04854_;
 wire _04855_;
 wire _04856_;
 wire _04857_;
 wire _04858_;
 wire _04859_;
 wire _04860_;
 wire _04861_;
 wire _04862_;
 wire _04863_;
 wire _04864_;
 wire _04865_;
 wire _04866_;
 wire _04867_;
 wire _04868_;
 wire _04869_;
 wire _04870_;
 wire _04871_;
 wire _04872_;
 wire _04873_;
 wire _04874_;
 wire _04875_;
 wire _04876_;
 wire _04877_;
 wire _04878_;
 wire _04879_;
 wire _04880_;
 wire _04881_;
 wire _04882_;
 wire _04883_;
 wire _04884_;
 wire _04885_;
 wire _04886_;
 wire _04887_;
 wire _04888_;
 wire _04889_;
 wire _04890_;
 wire _04891_;
 wire _04892_;
 wire _04893_;
 wire _04894_;
 wire _04895_;
 wire _04896_;
 wire _04897_;
 wire _04898_;
 wire _04899_;
 wire _04900_;
 wire _04901_;
 wire _04902_;
 wire _04903_;
 wire _04904_;
 wire _04905_;
 wire _04906_;
 wire _04907_;
 wire _04908_;
 wire _04909_;
 wire _04910_;
 wire _04911_;
 wire _04912_;
 wire _04913_;
 wire _04914_;
 wire _04915_;
 wire _04916_;
 wire _04917_;
 wire _04918_;
 wire _04919_;
 wire _04920_;
 wire _04921_;
 wire _04922_;
 wire _04923_;
 wire _04924_;
 wire _04925_;
 wire _04926_;
 wire _04927_;
 wire _04928_;
 wire _04929_;
 wire _04930_;
 wire _04931_;
 wire _04932_;
 wire _04933_;
 wire _04934_;
 wire _04935_;
 wire _04936_;
 wire _04937_;
 wire _04938_;
 wire _04939_;
 wire _04940_;
 wire _04941_;
 wire _04942_;
 wire _04943_;
 wire _04944_;
 wire _04945_;
 wire _04946_;
 wire _04947_;
 wire _04948_;
 wire _04949_;
 wire _04950_;
 wire _04951_;
 wire _04952_;
 wire _04953_;
 wire _04954_;
 wire _04955_;
 wire _04956_;
 wire _04957_;
 wire _04958_;
 wire _04959_;
 wire _04960_;
 wire _04961_;
 wire _04962_;
 wire _04963_;
 wire _04964_;
 wire _04965_;
 wire _04966_;
 wire _04967_;
 wire _04968_;
 wire _04969_;
 wire _04970_;
 wire _04971_;
 wire _04972_;
 wire _04973_;
 wire _04974_;
 wire _04975_;
 wire _04976_;
 wire _04977_;
 wire _04978_;
 wire _04979_;
 wire _04980_;
 wire _04981_;
 wire _04982_;
 wire _04983_;
 wire _04984_;
 wire _04985_;
 wire _04986_;
 wire _04987_;
 wire _04988_;
 wire _04989_;
 wire _04990_;
 wire _04991_;
 wire _04992_;
 wire _04993_;
 wire _04994_;
 wire _04995_;
 wire _04996_;
 wire _04997_;
 wire _04998_;
 wire _04999_;
 wire _05000_;
 wire _05001_;
 wire _05002_;
 wire _05003_;
 wire _05004_;
 wire _05005_;
 wire _05006_;
 wire _05007_;
 wire _05008_;
 wire _05009_;
 wire _05010_;
 wire _05011_;
 wire _05012_;
 wire _05013_;
 wire _05014_;
 wire _05015_;
 wire _05016_;
 wire _05017_;
 wire _05018_;
 wire _05019_;
 wire _05020_;
 wire _05021_;
 wire _05022_;
 wire _05023_;
 wire _05024_;
 wire _05025_;
 wire _05026_;
 wire _05027_;
 wire _05028_;
 wire _05029_;
 wire _05030_;
 wire _05031_;
 wire _05032_;
 wire _05033_;
 wire _05034_;
 wire _05035_;
 wire _05036_;
 wire _05037_;
 wire _05038_;
 wire _05039_;
 wire _05040_;
 wire _05041_;
 wire _05042_;
 wire _05043_;
 wire _05044_;
 wire _05045_;
 wire _05046_;
 wire _05047_;
 wire _05048_;
 wire _05049_;
 wire _05050_;
 wire _05051_;
 wire _05052_;
 wire _05053_;
 wire _05054_;
 wire _05055_;
 wire _05056_;
 wire _05057_;
 wire _05058_;
 wire _05059_;
 wire _05060_;
 wire _05061_;
 wire _05062_;
 wire _05063_;
 wire _05064_;
 wire _05065_;
 wire _05066_;
 wire _05067_;
 wire _05068_;
 wire _05069_;
 wire _05070_;
 wire _05071_;
 wire _05072_;
 wire _05073_;
 wire _05074_;
 wire _05075_;
 wire _05076_;
 wire _05077_;
 wire _05078_;
 wire _05079_;
 wire _05080_;
 wire _05081_;
 wire _05082_;
 wire _05083_;
 wire _05084_;
 wire _05085_;
 wire _05086_;
 wire _05087_;
 wire _05088_;
 wire _05089_;
 wire _05090_;
 wire _05091_;
 wire _05092_;
 wire _05093_;
 wire _05094_;
 wire _05095_;
 wire _05096_;
 wire _05097_;
 wire _05098_;
 wire _05099_;
 wire _05100_;
 wire _05101_;
 wire _05102_;
 wire _05103_;
 wire _05104_;
 wire _05105_;
 wire _05106_;
 wire _05107_;
 wire _05108_;
 wire _05109_;
 wire _05110_;
 wire _05111_;
 wire _05112_;
 wire _05113_;
 wire _05114_;
 wire _05115_;
 wire _05116_;
 wire _05117_;
 wire _05118_;
 wire _05119_;
 wire _05120_;
 wire _05121_;
 wire _05122_;
 wire _05123_;
 wire _05124_;
 wire _05125_;
 wire _05126_;
 wire _05127_;
 wire _05128_;
 wire _05129_;
 wire _05130_;
 wire _05131_;
 wire _05132_;
 wire _05133_;
 wire _05134_;
 wire _05135_;
 wire _05136_;
 wire _05137_;
 wire _05138_;
 wire _05139_;
 wire _05140_;
 wire _05141_;
 wire _05142_;
 wire _05143_;
 wire _05144_;
 wire _05145_;
 wire _05146_;
 wire _05147_;
 wire _05148_;
 wire _05149_;
 wire _05150_;
 wire _05151_;
 wire _05152_;
 wire _05153_;
 wire _05154_;
 wire _05155_;
 wire _05156_;
 wire _05157_;
 wire _05158_;
 wire _05159_;
 wire _05160_;
 wire _05161_;
 wire _05162_;
 wire _05163_;
 wire _05164_;
 wire _05165_;
 wire _05166_;
 wire _05167_;
 wire _05168_;
 wire _05169_;
 wire _05170_;
 wire _05171_;
 wire _05172_;
 wire _05173_;
 wire _05174_;
 wire _05175_;
 wire _05176_;
 wire _05177_;
 wire _05178_;
 wire _05179_;
 wire _05180_;
 wire _05181_;
 wire _05182_;
 wire _05183_;
 wire _05184_;
 wire _05185_;
 wire _05186_;
 wire _05187_;
 wire _05188_;
 wire _05189_;
 wire _05190_;
 wire _05191_;
 wire _05192_;
 wire _05193_;
 wire _05194_;
 wire _05195_;
 wire _05196_;
 wire _05197_;
 wire _05198_;
 wire _05199_;
 wire _05200_;
 wire _05201_;
 wire _05202_;
 wire _05203_;
 wire _05204_;
 wire _05205_;
 wire _05206_;
 wire _05207_;
 wire _05208_;
 wire _05209_;
 wire _05210_;
 wire _05211_;
 wire _05212_;
 wire _05213_;
 wire _05214_;
 wire _05215_;
 wire _05216_;
 wire _05217_;
 wire _05218_;
 wire _05219_;
 wire _05220_;
 wire _05221_;
 wire _05222_;
 wire _05223_;
 wire _05224_;
 wire _05225_;
 wire _05226_;
 wire _05227_;
 wire _05228_;
 wire _05229_;
 wire _05230_;
 wire _05231_;
 wire _05232_;
 wire _05233_;
 wire _05234_;
 wire _05235_;
 wire _05236_;
 wire _05237_;
 wire _05238_;
 wire _05239_;
 wire _05240_;
 wire _05241_;
 wire _05242_;
 wire _05243_;
 wire _05244_;
 wire _05245_;
 wire _05246_;
 wire _05247_;
 wire _05248_;
 wire _05249_;
 wire _05250_;
 wire _05251_;
 wire _05252_;
 wire _05253_;
 wire _05254_;
 wire _05255_;
 wire _05256_;
 wire _05257_;
 wire _05258_;
 wire _05259_;
 wire _05260_;
 wire _05261_;
 wire _05262_;
 wire _05263_;
 wire _05264_;
 wire _05265_;
 wire _05266_;
 wire _05267_;
 wire _05268_;
 wire _05269_;
 wire _05270_;
 wire _05271_;
 wire _05272_;
 wire _05273_;
 wire _05274_;
 wire _05275_;
 wire _05276_;
 wire _05277_;
 wire _05278_;
 wire _05279_;
 wire _05280_;
 wire _05281_;
 wire _05282_;
 wire _05283_;
 wire _05284_;
 wire _05285_;
 wire _05286_;
 wire _05287_;
 wire _05288_;
 wire _05289_;
 wire _05290_;
 wire _05291_;
 wire _05292_;
 wire _05293_;
 wire _05294_;
 wire _05295_;
 wire _05296_;
 wire _05297_;
 wire _05298_;
 wire _05299_;
 wire _05300_;
 wire _05301_;
 wire _05302_;
 wire _05303_;
 wire _05304_;
 wire _05305_;
 wire _05306_;
 wire _05307_;
 wire _05308_;
 wire _05309_;
 wire _05310_;
 wire _05311_;
 wire _05312_;
 wire _05313_;
 wire _05314_;
 wire _05315_;
 wire _05316_;
 wire _05317_;
 wire _05318_;
 wire _05319_;
 wire _05320_;
 wire _05321_;
 wire _05322_;
 wire _05323_;
 wire _05324_;
 wire _05325_;
 wire _05326_;
 wire _05327_;
 wire _05328_;
 wire _05329_;
 wire _05330_;
 wire _05331_;
 wire _05332_;
 wire _05333_;
 wire _05334_;
 wire _05335_;
 wire _05336_;
 wire _05337_;
 wire _05338_;
 wire _05339_;
 wire _05340_;
 wire _05341_;
 wire _05342_;
 wire _05343_;
 wire _05344_;
 wire _05345_;
 wire _05346_;
 wire _05347_;
 wire _05348_;
 wire _05349_;
 wire _05350_;
 wire _05351_;
 wire _05352_;
 wire _05353_;
 wire _05354_;
 wire _05355_;
 wire _05356_;
 wire _05357_;
 wire _05358_;
 wire _05359_;
 wire _05360_;
 wire _05361_;
 wire _05362_;
 wire _05363_;
 wire _05364_;
 wire _05365_;
 wire _05366_;
 wire _05367_;
 wire _05368_;
 wire _05369_;
 wire _05370_;
 wire _05371_;
 wire _05372_;
 wire _05373_;
 wire _05374_;
 wire _05375_;
 wire _05376_;
 wire _05377_;
 wire _05378_;
 wire _05379_;
 wire _05380_;
 wire _05381_;
 wire _05382_;
 wire _05383_;
 wire _05384_;
 wire _05385_;
 wire _05386_;
 wire _05387_;
 wire _05388_;
 wire _05389_;
 wire _05390_;
 wire _05391_;
 wire _05392_;
 wire _05393_;
 wire _05394_;
 wire _05395_;
 wire _05396_;
 wire _05397_;
 wire _05398_;
 wire _05399_;
 wire _05400_;
 wire _05401_;
 wire _05402_;
 wire _05403_;
 wire _05404_;
 wire _05405_;
 wire _05406_;
 wire _05407_;
 wire _05408_;
 wire _05409_;
 wire _05410_;
 wire _05411_;
 wire _05412_;
 wire _05413_;
 wire _05414_;
 wire _05415_;
 wire _05416_;
 wire _05417_;
 wire _05418_;
 wire _05419_;
 wire _05420_;
 wire _05421_;
 wire _05422_;
 wire _05423_;
 wire _05424_;
 wire _05425_;
 wire _05426_;
 wire _05427_;
 wire _05428_;
 wire _05429_;
 wire _05430_;
 wire _05431_;
 wire _05432_;
 wire _05433_;
 wire _05434_;
 wire _05435_;
 wire _05436_;
 wire _05437_;
 wire _05438_;
 wire _05439_;
 wire _05440_;
 wire _05441_;
 wire _05442_;
 wire _05443_;
 wire _05444_;
 wire _05445_;
 wire _05446_;
 wire _05447_;
 wire _05448_;
 wire _05449_;
 wire _05450_;
 wire _05451_;
 wire _05452_;
 wire _05453_;
 wire _05454_;
 wire _05455_;
 wire _05456_;
 wire _05457_;
 wire _05458_;
 wire _05459_;
 wire _05460_;
 wire _05461_;
 wire _05462_;
 wire _05463_;
 wire _05464_;
 wire _05465_;
 wire _05466_;
 wire _05467_;
 wire _05468_;
 wire _05469_;
 wire _05470_;
 wire _05471_;
 wire _05472_;
 wire _05473_;
 wire _05474_;
 wire _05475_;
 wire _05476_;
 wire _05477_;
 wire _05478_;
 wire _05479_;
 wire _05480_;
 wire _05481_;
 wire _05482_;
 wire _05483_;
 wire _05484_;
 wire _05485_;
 wire _05486_;
 wire _05487_;
 wire _05488_;
 wire _05489_;
 wire _05490_;
 wire _05491_;
 wire _05492_;
 wire _05493_;
 wire _05494_;
 wire _05495_;
 wire _05496_;
 wire _05497_;
 wire _05498_;
 wire _05499_;
 wire _05500_;
 wire _05501_;
 wire _05502_;
 wire _05503_;
 wire _05504_;
 wire _05505_;
 wire _05506_;
 wire _05507_;
 wire _05508_;
 wire _05509_;
 wire _05510_;
 wire _05511_;
 wire _05512_;
 wire _05513_;
 wire _05514_;
 wire _05515_;
 wire _05516_;
 wire _05517_;
 wire _05518_;
 wire _05519_;
 wire _05520_;
 wire _05521_;
 wire _05522_;
 wire _05523_;
 wire _05524_;
 wire _05525_;
 wire _05526_;
 wire _05527_;
 wire _05528_;
 wire _05529_;
 wire _05530_;
 wire _05531_;
 wire _05532_;
 wire _05533_;
 wire _05534_;
 wire _05535_;
 wire _05536_;
 wire _05537_;
 wire _05538_;
 wire _05539_;
 wire _05540_;
 wire _05541_;
 wire _05542_;
 wire _05543_;
 wire _05544_;
 wire _05545_;
 wire _05546_;
 wire _05547_;
 wire _05548_;
 wire _05549_;
 wire _05550_;
 wire _05551_;
 wire _05552_;
 wire _05553_;
 wire _05554_;
 wire _05555_;
 wire _05556_;
 wire _05557_;
 wire _05558_;
 wire _05559_;
 wire _05560_;
 wire _05561_;
 wire _05562_;
 wire _05563_;
 wire _05564_;
 wire _05565_;
 wire _05566_;
 wire _05567_;
 wire _05568_;
 wire _05569_;
 wire _05570_;
 wire _05571_;
 wire _05572_;
 wire _05573_;
 wire _05574_;
 wire _05575_;
 wire _05576_;
 wire _05577_;
 wire _05578_;
 wire _05579_;
 wire _05580_;
 wire _05581_;
 wire _05582_;
 wire _05583_;
 wire _05584_;
 wire _05585_;
 wire _05586_;
 wire _05587_;
 wire _05588_;
 wire _05589_;
 wire _05590_;
 wire _05591_;
 wire _05592_;
 wire _05593_;
 wire _05594_;
 wire _05595_;
 wire _05596_;
 wire _05597_;
 wire _05598_;
 wire _05599_;
 wire _05600_;
 wire _05601_;
 wire _05602_;
 wire _05603_;
 wire _05604_;
 wire _05605_;
 wire _05606_;
 wire _05607_;
 wire _05608_;
 wire _05609_;
 wire _05610_;
 wire _05611_;
 wire _05612_;
 wire _05613_;
 wire _05614_;
 wire _05615_;
 wire _05616_;
 wire _05617_;
 wire _05618_;
 wire _05619_;
 wire _05620_;
 wire _05621_;
 wire _05622_;
 wire _05623_;
 wire _05624_;
 wire _05625_;
 wire _05626_;
 wire _05627_;
 wire _05628_;
 wire _05629_;
 wire _05630_;
 wire _05631_;
 wire _05632_;
 wire _05633_;
 wire _05634_;
 wire _05635_;
 wire _05636_;
 wire _05637_;
 wire _05638_;
 wire _05639_;
 wire _05640_;
 wire _05641_;
 wire _05642_;
 wire _05643_;
 wire _05644_;
 wire _05645_;
 wire _05646_;
 wire _05647_;
 wire _05648_;
 wire _05649_;
 wire _05650_;
 wire _05651_;
 wire _05652_;
 wire _05653_;
 wire _05654_;
 wire _05655_;
 wire _05656_;
 wire _05657_;
 wire _05658_;
 wire _05659_;
 wire _05660_;
 wire _05661_;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire clknet_leaf_0_clk;
 wire \byte_counter[0] ;
 wire \byte_counter[1] ;
 wire \byte_counter[2] ;
 wire \byte_counter[3] ;
 wire \cmd_reg[0] ;
 wire \cmd_reg[1] ;
 wire \cmd_reg[2] ;
 wire \cmd_reg[3] ;
 wire \cmd_reg[4] ;
 wire \cmd_reg[5] ;
 wire \cmd_reg[6] ;
 wire \cmd_reg[7] ;
 wire \cordic_atan2_result[0] ;
 wire \cordic_atan2_result[10] ;
 wire \cordic_atan2_result[11] ;
 wire \cordic_atan2_result[12] ;
 wire \cordic_atan2_result[13] ;
 wire \cordic_atan2_result[14] ;
 wire \cordic_atan2_result[15] ;
 wire \cordic_atan2_result[16] ;
 wire \cordic_atan2_result[17] ;
 wire \cordic_atan2_result[18] ;
 wire \cordic_atan2_result[19] ;
 wire \cordic_atan2_result[1] ;
 wire \cordic_atan2_result[20] ;
 wire \cordic_atan2_result[21] ;
 wire \cordic_atan2_result[22] ;
 wire \cordic_atan2_result[23] ;
 wire \cordic_atan2_result[2] ;
 wire \cordic_atan2_result[3] ;
 wire \cordic_atan2_result[4] ;
 wire \cordic_atan2_result[5] ;
 wire \cordic_atan2_result[6] ;
 wire \cordic_atan2_result[7] ;
 wire \cordic_atan2_result[8] ;
 wire \cordic_atan2_result[9] ;
 wire cordic_busy;
 wire cordic_en_atan2;
 wire cordic_en_get_atan2;
 wire cordic_en_get_normalize;
 wire cordic_en_get_sin_cos;
 wire cordic_en_get_sqrt;
 wire cordic_en_normalize;
 wire cordic_en_sin_cos;
 wire cordic_en_sqrt;
 wire \cordic_inst.CASE_cordic_state_BITS_7_TO_3_0_262144_1_13107_ETC__q2[19] ;
 wire \cordic_inst.CASE_cordic_state_BITS_7_TO_3_0_3217_1_1901_2__ETC__q3[0] ;
 wire \cordic_inst.CASE_cordic_state_BITS_7_TO_3_0_3217_1_1901_2__ETC__q3[10] ;
 wire \cordic_inst.CASE_cordic_state_BITS_7_TO_3_0_3217_1_1901_2__ETC__q3[11] ;
 wire \cordic_inst.CASE_cordic_state_BITS_7_TO_3_0_3217_1_1901_2__ETC__q3[1] ;
 wire \cordic_inst.CASE_cordic_state_BITS_7_TO_3_0_3217_1_1901_2__ETC__q3[2] ;
 wire \cordic_inst.CASE_cordic_state_BITS_7_TO_3_0_3217_1_1901_2__ETC__q3[3] ;
 wire \cordic_inst.CASE_cordic_state_BITS_7_TO_3_0_3217_1_1901_2__ETC__q3[4] ;
 wire \cordic_inst.CASE_cordic_state_BITS_7_TO_3_0_3217_1_1901_2__ETC__q3[5] ;
 wire \cordic_inst.CASE_cordic_state_BITS_7_TO_3_0_3217_1_1901_2__ETC__q3[6] ;
 wire \cordic_inst.CASE_cordic_state_BITS_7_TO_3_0_3217_1_1901_2__ETC__q3[7] ;
 wire \cordic_inst.CASE_cordic_state_BITS_7_TO_3_0_3217_1_1901_2__ETC__q3[8] ;
 wire \cordic_inst.CASE_cordic_state_BITS_7_TO_3_0_3217_1_1901_2__ETC__q3[9] ;
 wire \cordic_inst.IF_IF_cordic_state_BITS_2_TO_1_EQ_1_THEN_NOT_c_ETC___d36[1] ;
 wire \cordic_inst.MUX_cordic_state$write_1__VAL_1[32] ;
 wire \cordic_inst.MUX_cordic_state$write_1__VAL_1[33] ;
 wire \cordic_inst.MUX_cordic_state$write_1__VAL_1[34] ;
 wire \cordic_inst.MUX_cordic_state$write_1__VAL_1[35] ;
 wire \cordic_inst.MUX_cordic_state$write_1__VAL_1[36] ;
 wire \cordic_inst.MUX_cordic_state$write_1__VAL_1[37] ;
 wire \cordic_inst.MUX_cordic_state$write_1__VAL_1[38] ;
 wire \cordic_inst.MUX_cordic_state$write_1__VAL_1[39] ;
 wire \cordic_inst.MUX_cordic_state$write_1__VAL_1[40] ;
 wire \cordic_inst.MUX_cordic_state$write_1__VAL_1[41] ;
 wire \cordic_inst.MUX_cordic_state$write_1__VAL_1[42] ;
 wire \cordic_inst.MUX_cordic_state$write_1__VAL_1[43] ;
 wire \cordic_inst.MUX_cordic_state$write_1__VAL_1[44] ;
 wire \cordic_inst.MUX_cordic_state$write_1__VAL_1[45] ;
 wire \cordic_inst.MUX_cordic_state$write_1__VAL_1[46] ;
 wire \cordic_inst.MUX_cordic_state$write_1__VAL_1[47] ;
 wire \cordic_inst.MUX_cordic_state$write_1__VAL_1[48] ;
 wire \cordic_inst.MUX_cordic_state$write_1__VAL_1[49] ;
 wire \cordic_inst.MUX_cordic_state$write_1__VAL_1[50] ;
 wire \cordic_inst.MUX_cordic_state$write_1__VAL_1[51] ;
 wire \cordic_inst.MUX_cordic_state$write_1__VAL_1[52] ;
 wire \cordic_inst.MUX_cordic_state$write_1__VAL_1[53] ;
 wire \cordic_inst.MUX_cordic_state$write_1__VAL_1[54] ;
 wire \cordic_inst.MUX_cordic_state$write_1__VAL_1[55] ;
 wire \cordic_inst.MUX_cordic_state$write_1__VAL_1[56] ;
 wire \cordic_inst.MUX_cordic_state$write_1__VAL_1[57] ;
 wire \cordic_inst.MUX_cordic_state$write_1__VAL_1[58] ;
 wire \cordic_inst.MUX_cordic_state$write_1__VAL_1[59] ;
 wire \cordic_inst.MUX_cordic_state$write_1__VAL_1[60] ;
 wire \cordic_inst.MUX_cordic_state$write_1__VAL_1[61] ;
 wire \cordic_inst.MUX_cordic_state$write_1__VAL_1[62] ;
 wire \cordic_inst.MUX_cordic_state$write_1__VAL_1[63] ;
 wire \cordic_inst.MUX_cordic_state$write_1__VAL_1[64] ;
 wire \cordic_inst.MUX_cordic_state$write_1__VAL_1[65] ;
 wire \cordic_inst.MUX_cordic_state$write_1__VAL_1[66] ;
 wire \cordic_inst.MUX_cordic_state$write_1__VAL_1[67] ;
 wire \cordic_inst.MUX_cordic_state$write_1__VAL_1[68] ;
 wire \cordic_inst.MUX_cordic_state$write_1__VAL_1[69] ;
 wire \cordic_inst.MUX_cordic_state$write_1__VAL_1[70] ;
 wire \cordic_inst.MUX_cordic_state$write_1__VAL_1[71] ;
 wire \cordic_inst.MUX_cordic_state$write_1__VAL_1[72] ;
 wire \cordic_inst.MUX_cordic_state$write_1__VAL_1[73] ;
 wire \cordic_inst.MUX_cordic_state$write_1__VAL_1[74] ;
 wire \cordic_inst.MUX_cordic_state$write_1__VAL_1[75] ;
 wire \cordic_inst.MUX_cordic_state$write_1__VAL_1[76] ;
 wire \cordic_inst.MUX_cordic_state$write_1__VAL_1[77] ;
 wire \cordic_inst.MUX_cordic_state$write_1__VAL_1[78] ;
 wire \cordic_inst.MUX_cordic_state$write_1__VAL_1[79] ;
 wire \cordic_inst.cordic_state[0] ;
 wire \cordic_inst.cordic_state[32] ;
 wire \cordic_inst.cordic_state[33] ;
 wire \cordic_inst.cordic_state[34] ;
 wire \cordic_inst.cordic_state[35] ;
 wire \cordic_inst.cordic_state[36] ;
 wire \cordic_inst.cordic_state[37] ;
 wire \cordic_inst.cordic_state[38] ;
 wire \cordic_inst.cordic_state[39] ;
 wire \cordic_inst.cordic_state[3] ;
 wire \cordic_inst.cordic_state[40] ;
 wire \cordic_inst.cordic_state[41] ;
 wire \cordic_inst.cordic_state[42] ;
 wire \cordic_inst.cordic_state[43] ;
 wire \cordic_inst.cordic_state[44] ;
 wire \cordic_inst.cordic_state[45] ;
 wire \cordic_inst.cordic_state[46] ;
 wire \cordic_inst.cordic_state[47] ;
 wire \cordic_inst.cordic_state[48] ;
 wire \cordic_inst.cordic_state[49] ;
 wire \cordic_inst.cordic_state[4] ;
 wire \cordic_inst.cordic_state[50] ;
 wire \cordic_inst.cordic_state[51] ;
 wire \cordic_inst.cordic_state[52] ;
 wire \cordic_inst.cordic_state[53] ;
 wire \cordic_inst.cordic_state[54] ;
 wire \cordic_inst.cordic_state[55] ;
 wire \cordic_inst.cordic_state[56] ;
 wire \cordic_inst.cordic_state[57] ;
 wire \cordic_inst.cordic_state[58] ;
 wire \cordic_inst.cordic_state[59] ;
 wire \cordic_inst.cordic_state[5] ;
 wire \cordic_inst.cordic_state[60] ;
 wire \cordic_inst.cordic_state[61] ;
 wire \cordic_inst.cordic_state[62] ;
 wire \cordic_inst.cordic_state[63] ;
 wire \cordic_inst.cordic_state[64] ;
 wire \cordic_inst.cordic_state[65] ;
 wire \cordic_inst.cordic_state[66] ;
 wire \cordic_inst.cordic_state[67] ;
 wire \cordic_inst.cordic_state[68] ;
 wire \cordic_inst.cordic_state[69] ;
 wire \cordic_inst.cordic_state[6] ;
 wire \cordic_inst.cordic_state[70] ;
 wire \cordic_inst.cordic_state[71] ;
 wire \cordic_inst.cordic_state[72] ;
 wire \cordic_inst.cordic_state[73] ;
 wire \cordic_inst.cordic_state[74] ;
 wire \cordic_inst.cordic_state[75] ;
 wire \cordic_inst.cordic_state[76] ;
 wire \cordic_inst.cordic_state[77] ;
 wire \cordic_inst.cordic_state[78] ;
 wire \cordic_inst.cordic_state[79] ;
 wire \cordic_inst.cordic_state[7] ;
 wire \cordic_inst.current_op[0] ;
 wire \cordic_inst.current_op[1] ;
 wire \cordic_inst.current_op[2] ;
 wire \cordic_inst.current_op[3] ;
 wire \cordic_inst.get_normalize[24] ;
 wire \cordic_inst.get_normalize[25] ;
 wire \cordic_inst.get_normalize[26] ;
 wire \cordic_inst.get_normalize[27] ;
 wire \cordic_inst.get_normalize[28] ;
 wire \cordic_inst.get_normalize[29] ;
 wire \cordic_inst.get_normalize[30] ;
 wire \cordic_inst.get_normalize[31] ;
 wire \cordic_inst.get_normalize[32] ;
 wire \cordic_inst.get_normalize[33] ;
 wire \cordic_inst.get_normalize[34] ;
 wire \cordic_inst.get_normalize[35] ;
 wire \cordic_inst.get_normalize[36] ;
 wire \cordic_inst.get_normalize[37] ;
 wire \cordic_inst.get_normalize[38] ;
 wire \cordic_inst.get_normalize[39] ;
 wire \cordic_inst.get_normalize[40] ;
 wire \cordic_inst.get_normalize[41] ;
 wire \cordic_inst.get_normalize[42] ;
 wire \cordic_inst.get_normalize[43] ;
 wire \cordic_inst.get_normalize[44] ;
 wire \cordic_inst.get_normalize[45] ;
 wire \cordic_inst.get_normalize[46] ;
 wire \cordic_inst.get_normalize[47] ;
 wire \cordic_inst.get_normalize[48] ;
 wire \cordic_inst.get_normalize[49] ;
 wire \cordic_inst.get_normalize[50] ;
 wire \cordic_inst.get_normalize[51] ;
 wire \cordic_inst.get_normalize[52] ;
 wire \cordic_inst.get_normalize[53] ;
 wire \cordic_inst.get_normalize[54] ;
 wire \cordic_inst.get_normalize[55] ;
 wire \cordic_inst.get_normalize[56] ;
 wire \cordic_inst.get_normalize[57] ;
 wire \cordic_inst.get_normalize[58] ;
 wire \cordic_inst.get_normalize[59] ;
 wire \cordic_inst.get_normalize[60] ;
 wire \cordic_inst.get_normalize[61] ;
 wire \cordic_inst.get_normalize[62] ;
 wire \cordic_inst.get_normalize[63] ;
 wire \cordic_inst.get_normalize[64] ;
 wire \cordic_inst.get_normalize[65] ;
 wire \cordic_inst.get_normalize[66] ;
 wire \cordic_inst.get_normalize[67] ;
 wire \cordic_inst.get_normalize[68] ;
 wire \cordic_inst.get_normalize[69] ;
 wire \cordic_inst.get_normalize[70] ;
 wire \cordic_inst.get_normalize[71] ;
 wire \cordic_inst.operation_pending ;
 wire \cordic_inst.operation_started ;
 wire \cordic_inst.result_ready ;
 wire \exec_phase[1] ;
 wire \exec_phase[2] ;
 wire mac_en_clear;
 wire mac_en_get_mac;
 wire mac_en_get_msu;
 wire mac_en_get_multiply;
 wire mac_en_mac;
 wire mac_en_msu;
 wire mac_en_multiply;
 wire \mac_inst.RDY_get_mac ;
 wire \mac_inst.RDY_get_msu ;
 wire \mac_inst.RDY_get_multiply ;
 wire \mac_inst.accumulator[0] ;
 wire \mac_inst.accumulator[10] ;
 wire \mac_inst.accumulator[11] ;
 wire \mac_inst.accumulator[12] ;
 wire \mac_inst.accumulator[13] ;
 wire \mac_inst.accumulator[14] ;
 wire \mac_inst.accumulator[15] ;
 wire \mac_inst.accumulator[16] ;
 wire \mac_inst.accumulator[17] ;
 wire \mac_inst.accumulator[18] ;
 wire \mac_inst.accumulator[19] ;
 wire \mac_inst.accumulator[1] ;
 wire \mac_inst.accumulator[20] ;
 wire \mac_inst.accumulator[21] ;
 wire \mac_inst.accumulator[22] ;
 wire \mac_inst.accumulator[23] ;
 wire \mac_inst.accumulator[2] ;
 wire \mac_inst.accumulator[3] ;
 wire \mac_inst.accumulator[4] ;
 wire \mac_inst.accumulator[5] ;
 wire \mac_inst.accumulator[6] ;
 wire \mac_inst.accumulator[7] ;
 wire \mac_inst.accumulator[8] ;
 wire \mac_inst.accumulator[9] ;
 wire \mac_inst.get_mac[0] ;
 wire \mac_inst.get_mac[10] ;
 wire \mac_inst.get_mac[11] ;
 wire \mac_inst.get_mac[12] ;
 wire \mac_inst.get_mac[13] ;
 wire \mac_inst.get_mac[14] ;
 wire \mac_inst.get_mac[15] ;
 wire \mac_inst.get_mac[16] ;
 wire \mac_inst.get_mac[17] ;
 wire \mac_inst.get_mac[18] ;
 wire \mac_inst.get_mac[19] ;
 wire \mac_inst.get_mac[1] ;
 wire \mac_inst.get_mac[20] ;
 wire \mac_inst.get_mac[21] ;
 wire \mac_inst.get_mac[22] ;
 wire \mac_inst.get_mac[23] ;
 wire \mac_inst.get_mac[2] ;
 wire \mac_inst.get_mac[3] ;
 wire \mac_inst.get_mac[4] ;
 wire \mac_inst.get_mac[5] ;
 wire \mac_inst.get_mac[6] ;
 wire \mac_inst.get_mac[7] ;
 wire \mac_inst.get_mac[8] ;
 wire \mac_inst.get_mac[9] ;
 wire \mac_inst.get_msu[0] ;
 wire \mac_inst.get_msu[10] ;
 wire \mac_inst.get_msu[11] ;
 wire \mac_inst.get_msu[12] ;
 wire \mac_inst.get_msu[13] ;
 wire \mac_inst.get_msu[14] ;
 wire \mac_inst.get_msu[15] ;
 wire \mac_inst.get_msu[16] ;
 wire \mac_inst.get_msu[17] ;
 wire \mac_inst.get_msu[18] ;
 wire \mac_inst.get_msu[19] ;
 wire \mac_inst.get_msu[1] ;
 wire \mac_inst.get_msu[20] ;
 wire \mac_inst.get_msu[21] ;
 wire \mac_inst.get_msu[22] ;
 wire \mac_inst.get_msu[23] ;
 wire \mac_inst.get_msu[2] ;
 wire \mac_inst.get_msu[3] ;
 wire \mac_inst.get_msu[4] ;
 wire \mac_inst.get_msu[5] ;
 wire \mac_inst.get_msu[6] ;
 wire \mac_inst.get_msu[7] ;
 wire \mac_inst.get_msu[8] ;
 wire \mac_inst.get_msu[9] ;
 wire \mac_inst.get_multiply[0] ;
 wire \mac_inst.get_multiply[10] ;
 wire \mac_inst.get_multiply[11] ;
 wire \mac_inst.get_multiply[12] ;
 wire \mac_inst.get_multiply[13] ;
 wire \mac_inst.get_multiply[14] ;
 wire \mac_inst.get_multiply[15] ;
 wire \mac_inst.get_multiply[16] ;
 wire \mac_inst.get_multiply[17] ;
 wire \mac_inst.get_multiply[18] ;
 wire \mac_inst.get_multiply[19] ;
 wire \mac_inst.get_multiply[1] ;
 wire \mac_inst.get_multiply[20] ;
 wire \mac_inst.get_multiply[21] ;
 wire \mac_inst.get_multiply[22] ;
 wire \mac_inst.get_multiply[23] ;
 wire \mac_inst.get_multiply[2] ;
 wire \mac_inst.get_multiply[3] ;
 wire \mac_inst.get_multiply[4] ;
 wire \mac_inst.get_multiply[5] ;
 wire \mac_inst.get_multiply[6] ;
 wire \mac_inst.get_multiply[7] ;
 wire \mac_inst.get_multiply[8] ;
 wire \mac_inst.get_multiply[9] ;
 wire rd_prev;
 wire \result_reg[0] ;
 wire \result_reg[10] ;
 wire \result_reg[11] ;
 wire \result_reg[12] ;
 wire \result_reg[13] ;
 wire \result_reg[14] ;
 wire \result_reg[15] ;
 wire \result_reg[16] ;
 wire \result_reg[17] ;
 wire \result_reg[18] ;
 wire \result_reg[19] ;
 wire \result_reg[1] ;
 wire \result_reg[20] ;
 wire \result_reg[21] ;
 wire \result_reg[22] ;
 wire \result_reg[23] ;
 wire \result_reg[24] ;
 wire \result_reg[25] ;
 wire \result_reg[26] ;
 wire \result_reg[27] ;
 wire \result_reg[28] ;
 wire \result_reg[29] ;
 wire \result_reg[2] ;
 wire \result_reg[30] ;
 wire \result_reg[31] ;
 wire \result_reg[32] ;
 wire \result_reg[33] ;
 wire \result_reg[34] ;
 wire \result_reg[35] ;
 wire \result_reg[36] ;
 wire \result_reg[37] ;
 wire \result_reg[38] ;
 wire \result_reg[39] ;
 wire \result_reg[3] ;
 wire \result_reg[40] ;
 wire \result_reg[41] ;
 wire \result_reg[42] ;
 wire \result_reg[43] ;
 wire \result_reg[44] ;
 wire \result_reg[45] ;
 wire \result_reg[46] ;
 wire \result_reg[47] ;
 wire \result_reg[48] ;
 wire \result_reg[49] ;
 wire \result_reg[4] ;
 wire \result_reg[50] ;
 wire \result_reg[51] ;
 wire \result_reg[52] ;
 wire \result_reg[53] ;
 wire \result_reg[54] ;
 wire \result_reg[55] ;
 wire \result_reg[56] ;
 wire \result_reg[57] ;
 wire \result_reg[58] ;
 wire \result_reg[59] ;
 wire \result_reg[5] ;
 wire \result_reg[60] ;
 wire \result_reg[61] ;
 wire \result_reg[62] ;
 wire \result_reg[63] ;
 wire \result_reg[64] ;
 wire \result_reg[65] ;
 wire \result_reg[66] ;
 wire \result_reg[67] ;
 wire \result_reg[68] ;
 wire \result_reg[69] ;
 wire \result_reg[6] ;
 wire \result_reg[70] ;
 wire \result_reg[71] ;
 wire \result_reg[7] ;
 wire \result_reg[8] ;
 wire \result_reg[9] ;
 wire \state[0] ;
 wire \state[1] ;
 wire \state[2] ;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire wr_prev;
 wire net1200;
 wire net1201;
 wire net1202;
 wire net1203;
 wire net1204;
 wire net1205;
 wire net1206;
 wire net1207;
 wire net1208;
 wire net1209;
 wire net1210;
 wire net1211;
 wire net1212;
 wire net1213;
 wire net1214;
 wire net1215;
 wire net1216;
 wire net1217;
 wire net1218;
 wire net1219;
 wire net1220;
 wire net1221;
 wire net1222;
 wire net1223;
 wire net1224;
 wire net1225;
 wire net1226;
 wire net1227;
 wire net1228;
 wire net1229;
 wire net1230;
 wire net1231;
 wire net1232;
 wire net1233;
 wire net1234;
 wire net1235;
 wire net1236;
 wire net1237;
 wire net1238;
 wire net1239;
 wire net1240;
 wire net1241;
 wire net1242;
 wire net1243;
 wire net1244;
 wire net1245;
 wire net1246;
 wire net1247;
 wire net1248;
 wire net1249;
 wire net1250;
 wire net1251;
 wire net1252;
 wire net1253;
 wire net1254;
 wire net1255;
 wire net1256;
 wire net1257;
 wire net1258;
 wire net1259;
 wire net1260;
 wire net1261;
 wire net1262;
 wire net1263;
 wire net1264;
 wire net1265;
 wire net1266;
 wire net1267;
 wire net1268;
 wire net1269;
 wire net1270;
 wire net1271;
 wire net1272;
 wire net1273;
 wire net1274;
 wire net1275;
 wire net1276;
 wire net1277;
 wire net1278;
 wire net1279;
 wire net1280;
 wire net1281;
 wire net1282;
 wire net1283;
 wire net1284;
 wire net1285;
 wire net1286;
 wire net1287;
 wire net1288;
 wire net1289;
 wire net1290;
 wire net1291;
 wire net1292;
 wire net1293;
 wire net1294;
 wire net1295;
 wire net1296;
 wire net1297;
 wire net1298;
 wire net1299;
 wire net1300;
 wire net1301;
 wire net1302;
 wire net1303;
 wire net1304;
 wire net1305;
 wire net1306;
 wire net1307;
 wire net1308;
 wire net1309;
 wire net1310;
 wire net1311;
 wire net1312;
 wire net1313;
 wire net1314;
 wire net1315;
 wire net1316;
 wire net1317;
 wire net1318;
 wire net1319;
 wire net1320;
 wire net1321;
 wire net1322;
 wire net1323;
 wire net1324;
 wire net1325;
 wire net1326;
 wire net1327;
 wire net1328;
 wire net1329;
 wire net1330;
 wire net1331;
 wire net1332;
 wire net1333;
 wire net1334;
 wire net1335;
 wire net1336;
 wire net1337;
 wire net1338;
 wire net1339;
 wire net1340;
 wire net1341;
 wire net1342;
 wire net1343;
 wire net1344;
 wire net1345;
 wire net1346;
 wire net1347;
 wire net1348;
 wire net1349;
 wire net1350;
 wire net1351;
 wire net1352;
 wire net1353;
 wire net1354;
 wire net1355;
 wire net1356;
 wire net1357;
 wire net1358;
 wire net1359;
 wire net1360;
 wire net1361;
 wire net1362;
 wire net1363;
 wire net1364;
 wire net1365;
 wire net1366;
 wire net1367;
 wire net1368;
 wire net1369;
 wire net1370;
 wire net1371;
 wire net1372;
 wire net1373;
 wire net1374;
 wire net1375;
 wire net1376;
 wire net1377;
 wire net1378;
 wire net1379;
 wire net1380;
 wire net1381;
 wire net1382;
 wire net1383;
 wire net1384;
 wire net1385;
 wire net1386;
 wire net1387;
 wire net1388;
 wire net1389;
 wire net1390;
 wire net1391;
 wire net1392;
 wire net1393;
 wire net1394;
 wire net1395;
 wire net1396;
 wire net1397;
 wire net1398;
 wire net1399;
 wire net1400;
 wire net1401;
 wire net1402;
 wire net1403;
 wire net1404;
 wire net1405;
 wire net1406;
 wire net1407;
 wire net1408;
 wire net1409;
 wire net1410;
 wire net1411;
 wire net1412;
 wire net1413;
 wire net1414;
 wire net1415;
 wire net1416;
 wire net1417;
 wire net1418;
 wire net1419;
 wire net1420;
 wire net1421;
 wire net1422;
 wire net1423;
 wire net1424;
 wire net1425;
 wire net1426;
 wire net1427;
 wire net1428;
 wire net1429;
 wire net1430;
 wire net1431;
 wire net1432;
 wire net1433;
 wire net1434;
 wire net1435;
 wire net1436;
 wire net1437;
 wire net1438;
 wire net1439;
 wire net1440;
 wire net1441;
 wire net1442;
 wire net1443;
 wire net1444;
 wire net1445;
 wire net1446;
 wire net1447;
 wire net1448;
 wire net1449;
 wire net1450;
 wire net1451;
 wire net1452;
 wire net1453;
 wire net1454;
 wire net1455;
 wire net1456;
 wire net1457;
 wire net1458;
 wire net1459;
 wire net1460;
 wire net1461;
 wire net1462;
 wire net1463;
 wire net1464;
 wire net1465;
 wire net1466;
 wire net1467;
 wire net1468;
 wire net1469;
 wire net1470;
 wire net1471;
 wire net1472;
 wire net1473;
 wire net1474;
 wire net1475;
 wire net1476;
 wire net1477;
 wire net1478;
 wire net1479;
 wire net1480;
 wire net1481;
 wire net1482;
 wire net1483;
 wire net1484;
 wire net1485;
 wire net1486;
 wire net1487;
 wire net1488;
 wire net1489;
 wire net1490;
 wire net1491;
 wire net1492;
 wire net1493;
 wire net1494;
 wire net1495;
 wire net1496;
 wire net1497;
 wire net1498;
 wire net1499;
 wire net1500;
 wire net1501;
 wire net1502;
 wire net1503;
 wire net1504;
 wire net1505;
 wire net1506;
 wire net1507;
 wire net1508;
 wire net1509;
 wire net1510;
 wire net1511;
 wire net1512;
 wire net1513;
 wire net1514;
 wire net1515;
 wire net1516;
 wire net1517;
 wire net1518;
 wire net1519;
 wire net1520;
 wire net1521;
 wire net1522;
 wire net1523;
 wire net1524;
 wire net1525;
 wire net1526;
 wire net1527;
 wire net1528;
 wire net1529;
 wire net1530;
 wire net1531;
 wire net1532;
 wire net1533;
 wire net1534;
 wire net1535;
 wire net1536;
 wire net1537;
 wire net1538;
 wire net1539;
 wire net1540;
 wire net1541;
 wire net1542;
 wire net1543;
 wire net1544;
 wire net1545;
 wire net1546;
 wire net1547;
 wire net1548;
 wire net1549;
 wire net1550;
 wire net1551;
 wire net1552;
 wire net1553;
 wire net1554;
 wire net1555;
 wire net1556;
 wire net1557;
 wire net1558;
 wire net1559;
 wire net1560;
 wire net1561;
 wire net1562;
 wire net1563;
 wire net1564;
 wire net1565;
 wire net1566;
 wire net1567;
 wire net1568;
 wire net1569;
 wire net1570;
 wire net1571;
 wire net1572;
 wire net1573;
 wire net1574;
 wire net1575;
 wire net1576;
 wire net1577;
 wire net1578;
 wire net1579;
 wire net1580;
 wire net1581;
 wire net1582;
 wire net1583;
 wire net1584;
 wire net1585;
 wire net1586;
 wire net1587;
 wire net1588;
 wire net1589;
 wire net1590;
 wire net1591;
 wire net1592;
 wire net1593;
 wire net1594;
 wire net1595;
 wire net1596;
 wire net1597;
 wire net1598;
 wire net1599;
 wire net1600;
 wire net1601;
 wire net1602;
 wire net1603;
 wire net1604;
 wire net1605;
 wire net1606;
 wire net1607;
 wire net1608;
 wire net1609;
 wire net1610;
 wire net1611;
 wire net1612;
 wire net1613;
 wire net1614;
 wire net1615;
 wire net1616;
 wire net1617;
 wire net1618;
 wire net1619;
 wire net1620;
 wire net1621;
 wire net1622;
 wire net1623;
 wire net1624;
 wire net1625;
 wire net1626;
 wire net1627;
 wire net1628;
 wire net1629;
 wire net1630;
 wire net1631;
 wire net1632;
 wire net1633;
 wire net1634;
 wire net1635;
 wire net1636;
 wire net1637;
 wire net1638;
 wire net1639;
 wire net1640;
 wire net1641;
 wire net1642;
 wire net1643;
 wire net1644;
 wire net1645;
 wire net1646;
 wire net1647;
 wire net1648;
 wire net1649;
 wire net1650;
 wire net1651;
 wire net1652;
 wire net1653;
 wire net1654;
 wire net1655;
 wire net1656;
 wire net1657;
 wire net1658;
 wire net1659;
 wire net1660;
 wire net1661;
 wire net1662;
 wire net1663;
 wire net1664;
 wire net1665;
 wire net1666;
 wire net1667;
 wire net1668;
 wire net1669;
 wire net1670;
 wire net1671;
 wire net1672;
 wire net1673;
 wire net1674;
 wire net1675;
 wire net1676;
 wire net1677;
 wire net1678;
 wire net1679;
 wire net1680;
 wire net1681;
 wire net1682;
 wire net1683;
 wire net1684;
 wire net1685;
 wire net1686;
 wire net1687;
 wire net1688;
 wire net1689;
 wire net1690;
 wire net1691;
 wire net1692;
 wire net1693;
 wire net1694;
 wire net1695;
 wire net1696;
 wire net1697;
 wire net1698;
 wire net1699;
 wire net1700;
 wire net1701;
 wire net1702;
 wire net1703;
 wire net1704;
 wire net1705;
 wire net1706;
 wire net1707;
 wire net1708;
 wire net1709;
 wire net1710;
 wire net1711;
 wire net1712;
 wire net1713;
 wire net1714;
 wire net1715;
 wire net1716;
 wire net1717;
 wire net1718;
 wire net1719;
 wire net1720;
 wire net1721;
 wire net1722;
 wire net1723;
 wire net1724;
 wire net1725;
 wire net1726;
 wire net1727;
 wire net1728;
 wire net1729;
 wire net1730;
 wire net1731;
 wire net1732;
 wire net1733;
 wire net1734;
 wire net1735;
 wire net1736;
 wire net1737;
 wire net1738;
 wire net1739;
 wire net1740;
 wire net1741;
 wire net1742;
 wire net1743;
 wire net1744;
 wire net1745;
 wire net1746;
 wire net1747;
 wire net1748;
 wire net1749;
 wire net1750;
 wire net1751;
 wire net1752;
 wire net1753;
 wire net1754;
 wire net1755;
 wire net1756;
 wire net1757;
 wire net1758;
 wire net1759;
 wire net1760;
 wire net1761;
 wire net1762;
 wire net1763;
 wire net1764;
 wire net1765;
 wire net1766;
 wire net1767;
 wire net1768;
 wire net1769;
 wire net1770;
 wire net1771;
 wire net1772;
 wire net1773;
 wire net1774;
 wire net1775;
 wire net1776;
 wire net1777;
 wire net1778;
 wire net1779;
 wire net1780;
 wire net1781;
 wire net1782;
 wire net1783;
 wire net1784;
 wire net1785;
 wire net1786;
 wire net1787;
 wire net1788;
 wire net1789;
 wire net1790;
 wire net1791;
 wire net1792;
 wire net1793;
 wire net1794;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_28_clk;
 wire clknet_leaf_29_clk;
 wire clknet_leaf_30_clk;
 wire clknet_leaf_31_clk;
 wire clknet_leaf_32_clk;
 wire clknet_leaf_33_clk;
 wire clknet_leaf_34_clk;
 wire clknet_leaf_35_clk;
 wire clknet_leaf_36_clk;
 wire clknet_leaf_37_clk;
 wire clknet_leaf_38_clk;
 wire clknet_leaf_39_clk;
 wire clknet_leaf_40_clk;
 wire clknet_leaf_41_clk;
 wire clknet_leaf_42_clk;
 wire clknet_leaf_43_clk;
 wire clknet_leaf_44_clk;
 wire clknet_leaf_45_clk;
 wire clknet_leaf_46_clk;
 wire clknet_leaf_47_clk;
 wire clknet_leaf_48_clk;
 wire clknet_leaf_49_clk;
 wire clknet_leaf_50_clk;
 wire clknet_leaf_51_clk;
 wire clknet_leaf_52_clk;
 wire clknet_leaf_53_clk;
 wire clknet_leaf_54_clk;
 wire clknet_leaf_55_clk;
 wire clknet_leaf_56_clk;
 wire clknet_leaf_57_clk;
 wire clknet_leaf_58_clk;
 wire clknet_leaf_59_clk;
 wire clknet_leaf_60_clk;
 wire clknet_leaf_61_clk;
 wire clknet_leaf_62_clk;
 wire clknet_leaf_63_clk;
 wire clknet_leaf_64_clk;
 wire clknet_leaf_65_clk;
 wire clknet_leaf_67_clk;
 wire clknet_leaf_68_clk;
 wire clknet_0_clk;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net860;
 wire net861;

 sg13g2_inv_1 _05909_ (.Y(_05531_),
    .A(net684));
 sg13g2_inv_1 _05910_ (.Y(_05532_),
    .A(\mac_inst.accumulator[18] ));
 sg13g2_inv_1 _05911_ (.Y(_05533_),
    .A(\mac_inst.accumulator[12] ));
 sg13g2_inv_1 _05912_ (.Y(_05534_),
    .A(\mac_inst.accumulator[11] ));
 sg13g2_inv_1 _05913_ (.Y(_05535_),
    .A(\mac_inst.accumulator[9] ));
 sg13g2_inv_1 _05914_ (.Y(_05536_),
    .A(\mac_inst.accumulator[5] ));
 sg13g2_inv_1 _05915_ (.Y(_05537_),
    .A(\mac_inst.accumulator[4] ));
 sg13g2_inv_1 _05916_ (.Y(_05538_),
    .A(\mac_inst.accumulator[3] ));
 sg13g2_inv_1 _05917_ (.Y(_05539_),
    .A(net1472));
 sg13g2_inv_1 _05918_ (.Y(_05540_),
    .A(net527));
 sg13g2_inv_1 _05919_ (.Y(_05541_),
    .A(net427));
 sg13g2_inv_1 _05920_ (.Y(_05542_),
    .A(net501));
 sg13g2_inv_1 _05921_ (.Y(_05543_),
    .A(net468));
 sg13g2_inv_1 _05922_ (.Y(_05544_),
    .A(net362));
 sg13g2_inv_1 _05923_ (.Y(_05545_),
    .A(net424));
 sg13g2_inv_1 _05924_ (.Y(_05546_),
    .A(net404));
 sg13g2_inv_1 _05925_ (.Y(_05547_),
    .A(net374));
 sg13g2_inv_1 _05926_ (.Y(_05548_),
    .A(net368));
 sg13g2_inv_1 _05927_ (.Y(_05549_),
    .A(net354));
 sg13g2_inv_1 _05928_ (.Y(_05550_),
    .A(net370));
 sg13g2_inv_1 _05929_ (.Y(_05551_),
    .A(net355));
 sg13g2_inv_4 _05930_ (.A(net1492),
    .Y(_05552_));
 sg13g2_inv_2 _05931_ (.Y(_05553_),
    .A(net1496));
 sg13g2_inv_1 _05932_ (.Y(_05554_),
    .A(net1513));
 sg13g2_inv_2 _05933_ (.Y(_05555_),
    .A(net1569));
 sg13g2_inv_2 _05934_ (.Y(_05556_),
    .A(net1606));
 sg13g2_inv_2 _05935_ (.Y(_05557_),
    .A(net1616));
 sg13g2_inv_4 _05936_ (.A(net1629),
    .Y(_05558_));
 sg13g2_inv_2 _05937_ (.Y(_05559_),
    .A(net1645));
 sg13g2_inv_1 _05938_ (.Y(_05560_),
    .A(net1656));
 sg13g2_inv_1 _05939_ (.Y(_05561_),
    .A(net1662));
 sg13g2_inv_1 _05940_ (.Y(_05562_),
    .A(net1670));
 sg13g2_inv_1 _05941_ (.Y(_05563_),
    .A(net1679));
 sg13g2_inv_2 _05942_ (.Y(_05564_),
    .A(net1684));
 sg13g2_inv_1 _05943_ (.Y(_05565_),
    .A(net1693));
 sg13g2_inv_1 _05944_ (.Y(_05566_),
    .A(net1703));
 sg13g2_inv_1 _05945_ (.Y(_05567_),
    .A(net1709));
 sg13g2_inv_1 _05946_ (.Y(_05568_),
    .A(net1714));
 sg13g2_inv_4 _05947_ (.A(net1727),
    .Y(_05569_));
 sg13g2_inv_4 _05948_ (.A(net1515),
    .Y(_05570_));
 sg13g2_inv_4 _05949_ (.A(net1526),
    .Y(_05571_));
 sg13g2_inv_1 _05950_ (.Y(_05572_),
    .A(net1542));
 sg13g2_inv_4 _05951_ (.A(net1546),
    .Y(_05573_));
 sg13g2_inv_4 _05952_ (.A(net1550),
    .Y(_05574_));
 sg13g2_inv_1 _05953_ (.Y(_05575_),
    .A(net499));
 sg13g2_inv_2 _05954_ (.Y(_05576_),
    .A(net1403));
 sg13g2_inv_1 _05955_ (.Y(_05577_),
    .A(\cordic_inst.cordic_state[77] ));
 sg13g2_inv_2 _05956_ (.Y(_05578_),
    .A(\cordic_inst.cordic_state[75] ));
 sg13g2_inv_1 _05957_ (.Y(_05579_),
    .A(net768));
 sg13g2_inv_1 _05958_ (.Y(_05580_),
    .A(net678));
 sg13g2_inv_1 _05959_ (.Y(_05581_),
    .A(\cordic_inst.cordic_state[57] ));
 sg13g2_inv_2 _05960_ (.Y(_05582_),
    .A(\cordic_inst.cordic_state[51] ));
 sg13g2_inv_2 _05961_ (.Y(_05583_),
    .A(net771));
 sg13g2_inv_2 _05962_ (.Y(_05584_),
    .A(net689));
 sg13g2_inv_1 _05963_ (.Y(_05585_),
    .A(\cordic_atan2_result[19] ));
 sg13g2_inv_1 _05964_ (.Y(_05586_),
    .A(\cordic_atan2_result[10] ));
 sg13g2_inv_1 _05965_ (.Y(_05587_),
    .A(net672));
 sg13g2_inv_1 _05966_ (.Y(_05588_),
    .A(net1427));
 sg13g2_inv_2 _05967_ (.Y(_05589_),
    .A(net1438));
 sg13g2_inv_2 _05968_ (.Y(_05590_),
    .A(net1443));
 sg13g2_inv_1 _05969_ (.Y(_05591_),
    .A(net1446));
 sg13g2_inv_1 _05970_ (.Y(_05592_),
    .A(net716));
 sg13g2_inv_1 _05971_ (.Y(_05593_),
    .A(net1753));
 sg13g2_inv_1 _05972_ (.Y(_05594_),
    .A(net1561));
 sg13g2_inv_2 _05973_ (.Y(_05595_),
    .A(net772));
 sg13g2_inv_1 _05974_ (.Y(_05596_),
    .A(\exec_phase[2] ));
 sg13g2_inv_1 _05975_ (.Y(_05597_),
    .A(net1467));
 sg13g2_inv_2 _05976_ (.Y(_05598_),
    .A(net574));
 sg13g2_nor2_1 _05977_ (.A(\state[0] ),
    .B(\state[1] ),
    .Y(_05599_));
 sg13g2_and2_1 _05978_ (.A(net1561),
    .B(_05599_),
    .X(_05600_));
 sg13g2_nand2_2 _05979_ (.Y(_05601_),
    .A(net1561),
    .B(_05599_));
 sg13g2_nor2_1 _05980_ (.A(\cmd_reg[7] ),
    .B(net789),
    .Y(_05602_));
 sg13g2_nand3b_1 _05981_ (.B(_05602_),
    .C(net619),
    .Y(_05603_),
    .A_N(net625));
 sg13g2_nor2_1 _05982_ (.A(net691),
    .B(net718),
    .Y(_05604_));
 sg13g2_nor4_2 _05983_ (.A(net1560),
    .B(net715),
    .C(net691),
    .Y(_05605_),
    .D(net718));
 sg13g2_nor2b_1 _05984_ (.A(_05603_),
    .B_N(_05605_),
    .Y(_05606_));
 sg13g2_nand2b_2 _05985_ (.Y(_05607_),
    .B(_05605_),
    .A_N(_05603_));
 sg13g2_nand2_2 _05986_ (.Y(_05608_),
    .A(net715),
    .B(_05604_));
 sg13g2_nor2_1 _05987_ (.A(_05603_),
    .B(_05608_),
    .Y(_05609_));
 sg13g2_or2_1 _05988_ (.X(_05610_),
    .B(_05608_),
    .A(_05603_));
 sg13g2_nand2_1 _05989_ (.Y(_05611_),
    .A(_05607_),
    .B(_05610_));
 sg13g2_a21oi_1 _05990_ (.A1(_05607_),
    .A2(_05610_),
    .Y(_05612_),
    .B1(_05601_));
 sg13g2_nand3b_1 _05991_ (.B(net625),
    .C(_05602_),
    .Y(_05613_),
    .A_N(net824));
 sg13g2_inv_1 _05992_ (.Y(_05614_),
    .A(_05613_));
 sg13g2_nor4_2 _05993_ (.A(net691),
    .B(net718),
    .C(_05601_),
    .Y(_05615_),
    .D(_05613_));
 sg13g2_nor2_2 _05994_ (.A(_05612_),
    .B(_05615_),
    .Y(_05616_));
 sg13g2_o21ai_1 _05995_ (.B1(_05616_),
    .Y(_05617_),
    .A1(net1561),
    .A2(_05599_));
 sg13g2_nor2b_2 _05996_ (.A(net810),
    .B_N(net724),
    .Y(_05618_));
 sg13g2_nand2_2 _05997_ (.Y(_05619_),
    .A(_05594_),
    .B(_05618_));
 sg13g2_nand3b_1 _05998_ (.B(_05604_),
    .C(net693),
    .Y(_05620_),
    .A_N(net715));
 sg13g2_or2_1 _05999_ (.X(_05621_),
    .B(_05620_),
    .A(_05603_));
 sg13g2_nor2b_2 _06000_ (.A(_05619_),
    .B_N(_05621_),
    .Y(_05622_));
 sg13g2_nor2b_2 _06001_ (.A(net1561),
    .B_N(net810),
    .Y(_05623_));
 sg13g2_nor2b_2 _06002_ (.A(net806),
    .B_N(net9),
    .Y(_05624_));
 sg13g2_nand2b_1 _06003_ (.Y(_05625_),
    .B(net9),
    .A_N(wr_prev));
 sg13g2_nand2b_2 _06004_ (.Y(_05626_),
    .B(net774),
    .A_N(net1465));
 sg13g2_nor3_1 _06005_ (.A(net1464),
    .B(\byte_counter[3] ),
    .C(_05626_),
    .Y(_05627_));
 sg13g2_nand2_1 _06006_ (.Y(_05628_),
    .A(_05624_),
    .B(net1326));
 sg13g2_nor2_2 _06007_ (.A(net790),
    .B(_05598_),
    .Y(_05629_));
 sg13g2_nand2_1 _06008_ (.Y(_05630_),
    .A(_05596_),
    .B(_00028_));
 sg13g2_and2_1 _06009_ (.A(net663),
    .B(_05629_),
    .X(_05631_));
 sg13g2_nand2b_1 _06010_ (.Y(_05632_),
    .B(net1318),
    .A_N(\mac_inst.RDY_get_multiply ));
 sg13g2_nor2_1 _06011_ (.A(net1560),
    .B(_05610_),
    .Y(_05633_));
 sg13g2_inv_1 _06012_ (.Y(_05634_),
    .A(net1276));
 sg13g2_o21ai_1 _06013_ (.B1(_05632_),
    .Y(_05635_),
    .A1(\mac_inst.RDY_get_mac ),
    .A2(_05634_));
 sg13g2_and2_1 _06014_ (.A(net1560),
    .B(_05609_),
    .X(_05636_));
 sg13g2_nand2_2 _06015_ (.Y(_05637_),
    .A(net1560),
    .B(_05609_));
 sg13g2_nor2_2 _06016_ (.A(_05608_),
    .B(_05613_),
    .Y(_05638_));
 sg13g2_nor3_1 _06017_ (.A(net1560),
    .B(_05608_),
    .C(_05613_),
    .Y(_05639_));
 sg13g2_nand2b_2 _06018_ (.Y(_05640_),
    .B(_05638_),
    .A_N(net1560));
 sg13g2_nand3_1 _06019_ (.B(\cordic_inst.cordic_state[0] ),
    .C(\cordic_inst.current_op[3] ),
    .A(\cordic_inst.result_ready ),
    .Y(_05641_));
 sg13g2_nand2_1 _06020_ (.Y(_05642_),
    .A(net1313),
    .B(_05641_));
 sg13g2_o21ai_1 _06021_ (.B1(_05642_),
    .Y(_05643_),
    .A1(\mac_inst.RDY_get_msu ),
    .A2(_05637_));
 sg13g2_o21ai_1 _06022_ (.B1(_05631_),
    .Y(_05644_),
    .A1(_05635_),
    .A2(_05643_));
 sg13g2_nand2_2 _06023_ (.Y(_05645_),
    .A(_05605_),
    .B(_05614_));
 sg13g2_inv_1 _06024_ (.Y(_05646_),
    .A(_05645_));
 sg13g2_nand2_1 _06025_ (.Y(_05647_),
    .A(_05640_),
    .B(_05645_));
 sg13g2_nand3_1 _06026_ (.B(_00028_),
    .C(_05647_),
    .A(\exec_phase[2] ),
    .Y(_05648_));
 sg13g2_nor2_1 _06027_ (.A(\exec_phase[1] ),
    .B(_05630_),
    .Y(_05649_));
 sg13g2_nand2b_2 _06028_ (.Y(_05650_),
    .B(_05629_),
    .A_N(\exec_phase[1] ));
 sg13g2_o21ai_1 _06029_ (.B1(_05649_),
    .Y(_05651_),
    .A1(net1318),
    .A2(net1276));
 sg13g2_nand3_1 _06030_ (.B(_05648_),
    .C(_05651_),
    .A(_05644_),
    .Y(_05652_));
 sg13g2_nand2_1 _06031_ (.Y(_05653_),
    .A(_05600_),
    .B(_05652_));
 sg13g2_nand3_1 _06032_ (.B(\cordic_inst.cordic_state[0] ),
    .C(\cordic_inst.current_op[0] ),
    .A(\cordic_inst.result_ready ),
    .Y(_05654_));
 sg13g2_nand3_1 _06033_ (.B(_05646_),
    .C(_05654_),
    .A(_05631_),
    .Y(_05655_));
 sg13g2_a22oi_1 _06034_ (.Y(_05656_),
    .B1(_05650_),
    .B2(_05655_),
    .A2(_05645_),
    .A1(_05637_));
 sg13g2_nor2_1 _06035_ (.A(_05601_),
    .B(_05629_),
    .Y(_05657_));
 sg13g2_a22oi_1 _06036_ (.Y(_05658_),
    .B1(_05657_),
    .B2(net1276),
    .A2(_05656_),
    .A1(_05600_));
 sg13g2_o21ai_1 _06037_ (.B1(_05625_),
    .Y(_05659_),
    .A1(_05622_),
    .A2(net1382));
 sg13g2_o21ai_1 _06038_ (.B1(_05657_),
    .Y(_05660_),
    .A1(net1318),
    .A2(net1271));
 sg13g2_nand2_2 _06039_ (.Y(_05661_),
    .A(_05598_),
    .B(_05600_));
 sg13g2_nor2_1 _06040_ (.A(_05645_),
    .B(_05661_),
    .Y(_00013_));
 sg13g2_and2_1 _06041_ (.A(net1560),
    .B(_05638_),
    .X(_00411_));
 sg13g2_nand2_1 _06042_ (.Y(_00412_),
    .A(net1560),
    .B(_05638_));
 sg13g2_nor2_1 _06043_ (.A(_05661_),
    .B(net1254),
    .Y(_00012_));
 sg13g2_nand3_1 _06044_ (.B(net1313),
    .C(_05649_),
    .A(_05600_),
    .Y(_00413_));
 sg13g2_nand2_1 _06045_ (.Y(_00414_),
    .A(_05660_),
    .B(_00413_));
 sg13g2_nor3_1 _06046_ (.A(_00013_),
    .B(_00012_),
    .C(_00414_),
    .Y(_00415_));
 sg13g2_nand4_1 _06047_ (.B(_05658_),
    .C(_05659_),
    .A(_05653_),
    .Y(_00416_),
    .D(_00415_));
 sg13g2_nand2_1 _06048_ (.Y(_00417_),
    .A(net1561),
    .B(_05618_));
 sg13g2_nor2b_1 _06049_ (.A(rd_prev),
    .B_N(net10),
    .Y(_00418_));
 sg13g2_nor2b_2 _06050_ (.A(_00417_),
    .B_N(_00418_),
    .Y(_00419_));
 sg13g2_nor2_1 _06051_ (.A(_05646_),
    .B(net1260),
    .Y(_00420_));
 sg13g2_nor4_2 _06052_ (.A(\byte_counter[1] ),
    .B(net1465),
    .C(net1464),
    .Y(_00421_),
    .D(_05595_));
 sg13g2_nand2b_2 _06053_ (.Y(_00422_),
    .B(net1465),
    .A_N(\byte_counter[1] ));
 sg13g2_nand2_2 _06054_ (.Y(_00423_),
    .A(net1464),
    .B(_05595_));
 sg13g2_nor2_2 _06055_ (.A(_00422_),
    .B(_00423_),
    .Y(_00424_));
 sg13g2_nor2b_1 _06056_ (.A(_05645_),
    .B_N(net1306),
    .Y(_00425_));
 sg13g2_a221oi_1 _06057_ (.B2(net1260),
    .C1(_00425_),
    .B1(net1325),
    .A1(net1326),
    .Y(_00426_),
    .A2(_00420_));
 sg13g2_inv_1 _06058_ (.Y(_00427_),
    .A(_00426_));
 sg13g2_nor2_1 _06059_ (.A(_05637_),
    .B(_05661_),
    .Y(_00020_));
 sg13g2_nor3_1 _06060_ (.A(_05598_),
    .B(_05601_),
    .C(_05621_),
    .Y(_00428_));
 sg13g2_or2_1 _06061_ (.X(_00429_),
    .B(_05620_),
    .A(_05613_));
 sg13g2_inv_1 _06062_ (.Y(_00430_),
    .A(_00429_));
 sg13g2_and4_1 _06063_ (.A(\cordic_inst.result_ready ),
    .B(\cordic_inst.cordic_state[0] ),
    .C(\cordic_inst.current_op[1] ),
    .D(_05631_),
    .X(_00431_));
 sg13g2_nor3_1 _06064_ (.A(_05601_),
    .B(_00429_),
    .C(_00431_),
    .Y(_00432_));
 sg13g2_or3_1 _06065_ (.A(\mac_inst.RDY_get_mac ),
    .B(\mac_inst.RDY_get_msu ),
    .C(\mac_inst.RDY_get_multiply ),
    .X(_00433_));
 sg13g2_nor2_2 _06066_ (.A(_05621_),
    .B(_05661_),
    .Y(_00015_));
 sg13g2_nand2_1 _06067_ (.Y(_00434_),
    .A(_00433_),
    .B(_00015_));
 sg13g2_nand3_1 _06068_ (.B(\cordic_inst.cordic_state[0] ),
    .C(\cordic_inst.current_op[2] ),
    .A(\cordic_inst.result_ready ),
    .Y(_00435_));
 sg13g2_a22oi_1 _06069_ (.Y(_00436_),
    .B1(_05631_),
    .B2(_00435_),
    .A2(_00028_),
    .A1(\exec_phase[2] ));
 sg13g2_nand2_1 _06070_ (.Y(_00437_),
    .A(_05600_),
    .B(net1258));
 sg13g2_nand2_2 _06071_ (.Y(_00438_),
    .A(_05600_),
    .B(_05631_));
 sg13g2_a21oi_1 _06072_ (.A1(_05650_),
    .A2(_00436_),
    .Y(_00439_),
    .B1(_00437_));
 sg13g2_nor2_1 _06073_ (.A(_05640_),
    .B(_05661_),
    .Y(_00007_));
 sg13g2_nor3_2 _06074_ (.A(net1561),
    .B(net724),
    .C(\state[1] ),
    .Y(_00440_));
 sg13g2_nand2_1 _06075_ (.Y(_00441_),
    .A(_05625_),
    .B(_00440_));
 sg13g2_nand2_1 _06076_ (.Y(_00442_),
    .A(net1382),
    .B(_05624_));
 sg13g2_o21ai_1 _06077_ (.B1(_00441_),
    .Y(_00443_),
    .A1(net1326),
    .A2(_00442_));
 sg13g2_nor2_1 _06078_ (.A(_00417_),
    .B(_00418_),
    .Y(_00444_));
 sg13g2_nor3_1 _06079_ (.A(_00007_),
    .B(_00443_),
    .C(_00444_),
    .Y(_00445_));
 sg13g2_nor4_1 _06080_ (.A(_00020_),
    .B(_00428_),
    .C(_00432_),
    .D(_00439_),
    .Y(_00446_));
 sg13g2_nand4_1 _06081_ (.B(_00434_),
    .C(_00445_),
    .A(_00413_),
    .Y(_00447_),
    .D(_00446_));
 sg13g2_a21oi_1 _06082_ (.A1(net1307),
    .A2(_00426_),
    .Y(_00448_),
    .B1(_00447_));
 sg13g2_nand2b_2 _06083_ (.Y(_00449_),
    .B(_00448_),
    .A_N(_00416_));
 sg13g2_nand2_1 _06084_ (.Y(_00450_),
    .A(net1382),
    .B(_05628_));
 sg13g2_inv_1 _06085_ (.Y(_00451_),
    .A(_00450_));
 sg13g2_nor4_1 _06086_ (.A(net1318),
    .B(net1276),
    .C(_05638_),
    .D(_00430_),
    .Y(_00452_));
 sg13g2_nor2_1 _06087_ (.A(net724),
    .B(_00442_),
    .Y(_00453_));
 sg13g2_nand2_2 _06088_ (.Y(_00454_),
    .A(net1326),
    .B(_00453_));
 sg13g2_o21ai_1 _06089_ (.B1(_05617_),
    .Y(_00455_),
    .A1(_00452_),
    .A2(_00454_));
 sg13g2_nor3_2 _06090_ (.A(_05622_),
    .B(_00451_),
    .C(_00455_),
    .Y(_00456_));
 sg13g2_and2_1 _06091_ (.A(_05616_),
    .B(_00456_),
    .X(_00457_));
 sg13g2_o21ai_1 _06092_ (.B1(_05616_),
    .Y(_00029_),
    .A1(_05598_),
    .A2(_00456_));
 sg13g2_and2_1 _06093_ (.A(cordic_en_normalize),
    .B(net1767),
    .X(_00458_));
 sg13g2_nor2_2 _06094_ (.A(cordic_en_normalize),
    .B(cordic_en_sqrt),
    .Y(_00459_));
 sg13g2_or2_1 _06095_ (.X(_00460_),
    .B(cordic_en_sqrt),
    .A(cordic_en_normalize));
 sg13g2_nor2_2 _06096_ (.A(net1474),
    .B(net1360),
    .Y(_00461_));
 sg13g2_nor2_2 _06097_ (.A(net1484),
    .B(net1478),
    .Y(_00462_));
 sg13g2_and2_1 _06098_ (.A(net1371),
    .B(net1359),
    .X(_00463_));
 sg13g2_nand2_2 _06099_ (.Y(_00464_),
    .A(net1372),
    .B(net1359));
 sg13g2_nor2_1 _06100_ (.A(net1746),
    .B(net1323),
    .Y(_00465_));
 sg13g2_nand2_1 _06101_ (.Y(_00466_),
    .A(net1770),
    .B(_00463_));
 sg13g2_a21o_1 _06102_ (.A2(_00465_),
    .A1(net545),
    .B1(net1373),
    .X(_00024_));
 sg13g2_nor2_1 _06103_ (.A(cordic_busy),
    .B(_05596_),
    .Y(_00467_));
 sg13g2_a21oi_1 _06104_ (.A1(_05615_),
    .A2(_00467_),
    .Y(_00468_),
    .B1(net663));
 sg13g2_nor2_1 _06105_ (.A(_05596_),
    .B(_00433_),
    .Y(_00469_));
 sg13g2_nand2_1 _06106_ (.Y(_00470_),
    .A(_05612_),
    .B(_00469_));
 sg13g2_o21ai_1 _06107_ (.B1(_00470_),
    .Y(_00026_),
    .A1(_00457_),
    .A2(net664));
 sg13g2_nor2_1 _06108_ (.A(_05661_),
    .B(_00429_),
    .Y(_00014_));
 sg13g2_nor2_1 _06109_ (.A(_05607_),
    .B(_05661_),
    .Y(_00021_));
 sg13g2_nor2_1 _06110_ (.A(_05634_),
    .B(_05661_),
    .Y(_00019_));
 sg13g2_a22oi_1 _06111_ (.Y(_00471_),
    .B1(_00433_),
    .B2(_05612_),
    .A2(_05615_),
    .A1(cordic_busy));
 sg13g2_a21o_1 _06112_ (.A2(_00471_),
    .A1(_00456_),
    .B1(_05596_),
    .X(_00472_));
 sg13g2_o21ai_1 _06113_ (.B1(_00472_),
    .Y(_00027_),
    .A1(net574),
    .A2(_05616_));
 sg13g2_o21ai_1 _06114_ (.B1(_00461_),
    .Y(_00473_),
    .A1(cordic_en_sin_cos),
    .A2(net661));
 sg13g2_nand2_1 _06115_ (.Y(_00022_),
    .A(net1768),
    .B(net662));
 sg13g2_nor2_1 _06116_ (.A(cordic_en_normalize),
    .B(net1747),
    .Y(_00474_));
 sg13g2_a22oi_1 _06117_ (.Y(_00475_),
    .B1(net1350),
    .B2(cordic_en_sqrt),
    .A2(_00465_),
    .A1(net564));
 sg13g2_inv_1 _06118_ (.Y(_00023_),
    .A(net565));
 sg13g2_and2_1 _06119_ (.A(net1477),
    .B(net1371),
    .X(_00476_));
 sg13g2_a21oi_1 _06120_ (.A1(net523),
    .A2(_00463_),
    .Y(_00477_),
    .B1(net1322));
 sg13g2_nor2_1 _06121_ (.A(net1746),
    .B(_00477_),
    .Y(_00025_));
 sg13g2_nor2b_2 _06122_ (.A(\cordic_inst.cordic_state[0] ),
    .B_N(cordic_busy),
    .Y(_00478_));
 sg13g2_nand2_2 _06123_ (.Y(_00479_),
    .A(_05592_),
    .B(cordic_busy));
 sg13g2_nor2_1 _06124_ (.A(net1323),
    .B(net1348),
    .Y(_00480_));
 sg13g2_nand2_1 _06125_ (.Y(_00481_),
    .A(_00463_),
    .B(_00479_));
 sg13g2_nor2_2 _06126_ (.A(net1480),
    .B(_00479_),
    .Y(_00482_));
 sg13g2_nand2b_2 _06127_ (.Y(_00483_),
    .B(net1349),
    .A_N(net1484));
 sg13g2_nor2_2 _06128_ (.A(net1475),
    .B(_00483_),
    .Y(_00484_));
 sg13g2_nand2_2 _06129_ (.Y(_00485_),
    .A(net1359),
    .B(net1348));
 sg13g2_nor2_2 _06130_ (.A(net1360),
    .B(_00485_),
    .Y(_00486_));
 sg13g2_and2_1 _06131_ (.A(net1446),
    .B(net1456),
    .X(_00487_));
 sg13g2_nand3_1 _06132_ (.B(net1446),
    .C(net1458),
    .A(net1443),
    .Y(_00488_));
 sg13g2_or2_1 _06133_ (.X(_00489_),
    .B(_00488_),
    .A(net1391));
 sg13g2_nand2_1 _06134_ (.Y(_00490_),
    .A(_00486_),
    .B(_00489_));
 sg13g2_inv_1 _06135_ (.Y(_00491_),
    .A(_00490_));
 sg13g2_o21ai_1 _06136_ (.B1(net1427),
    .Y(_00492_),
    .A1(net1293),
    .A2(_00491_));
 sg13g2_nand3b_1 _06137_ (.B(net1397),
    .C(_00486_),
    .Y(_00493_),
    .A_N(_00489_));
 sg13g2_and3_2 _06138_ (.X(_00494_),
    .A(net1754),
    .B(_00492_),
    .C(_00493_));
 sg13g2_inv_1 _06139_ (.Y(_00188_),
    .A(_00494_));
 sg13g2_or2_1 _06140_ (.X(_00495_),
    .B(_00487_),
    .A(net1443));
 sg13g2_nand3_1 _06141_ (.B(_00488_),
    .C(_00495_),
    .A(_00486_),
    .Y(_00496_));
 sg13g2_nand2_1 _06142_ (.Y(_00497_),
    .A(net1443),
    .B(net1293));
 sg13g2_and3_2 _06143_ (.X(_00498_),
    .A(net1754),
    .B(_00496_),
    .C(_00497_));
 sg13g2_inv_2 _06144_ (.Y(_00186_),
    .A(_00498_));
 sg13g2_nand2_2 _06145_ (.Y(_00499_),
    .A(net1391),
    .B(_00488_));
 sg13g2_o21ai_1 _06146_ (.B1(_00499_),
    .Y(_00500_),
    .A1(net1438),
    .A2(_00486_));
 sg13g2_a21oi_2 _06147_ (.B1(_00500_),
    .Y(_00501_),
    .A2(_00490_),
    .A1(net1285));
 sg13g2_a22oi_1 _06148_ (.Y(_00502_),
    .B1(_00491_),
    .B2(_00499_),
    .A2(net1294),
    .A1(net1438));
 sg13g2_nor2_2 _06149_ (.A(_00186_),
    .B(_00501_),
    .Y(_00503_));
 sg13g2_or2_1 _06150_ (.X(_00504_),
    .B(_00503_),
    .A(_00494_));
 sg13g2_inv_1 _06151_ (.Y(_00030_),
    .A(_00504_));
 sg13g2_nand2_1 _06152_ (.Y(_00505_),
    .A(_00494_),
    .B(_00498_));
 sg13g2_nor2_2 _06153_ (.A(net1446),
    .B(net1456),
    .Y(_00506_));
 sg13g2_or2_1 _06154_ (.X(_00507_),
    .B(net1456),
    .A(net1446));
 sg13g2_nor2_1 _06155_ (.A(_00487_),
    .B(_00506_),
    .Y(_00508_));
 sg13g2_a22oi_1 _06156_ (.Y(_00509_),
    .B1(_00486_),
    .B2(_00508_),
    .A2(net1294),
    .A1(net1446));
 sg13g2_nor2_2 _06157_ (.A(net1736),
    .B(_00509_),
    .Y(_00185_));
 sg13g2_nand2b_1 _06158_ (.Y(_00510_),
    .B(_00486_),
    .A_N(net1458));
 sg13g2_nand2_1 _06159_ (.Y(_00511_),
    .A(net1458),
    .B(net1294));
 sg13g2_nand3_1 _06160_ (.B(_00510_),
    .C(_00511_),
    .A(net1754),
    .Y(_00184_));
 sg13g2_o21ai_1 _06161_ (.B1(_00185_),
    .Y(_00512_),
    .A1(_00502_),
    .A2(_00184_));
 sg13g2_o21ai_1 _06162_ (.B1(_00504_),
    .Y(_00001_),
    .A1(_00505_),
    .A2(_00512_));
 sg13g2_nand2_1 _06163_ (.Y(_00513_),
    .A(_00498_),
    .B(_00184_));
 sg13g2_nand2_1 _06164_ (.Y(_00514_),
    .A(net1754),
    .B(_00501_));
 sg13g2_inv_1 _06165_ (.Y(_00187_),
    .A(_00514_));
 sg13g2_nand2_1 _06166_ (.Y(_00515_),
    .A(_00509_),
    .B(_00187_));
 sg13g2_o21ai_1 _06167_ (.B1(_00504_),
    .Y(_00006_),
    .A1(_00513_),
    .A2(_00515_));
 sg13g2_nand4_1 _06168_ (.B(_00509_),
    .C(_00510_),
    .A(net1754),
    .Y(_00516_),
    .D(_00511_));
 sg13g2_a21oi_1 _06169_ (.A1(_00503_),
    .A2(_00516_),
    .Y(_00517_),
    .B1(_00006_));
 sg13g2_a21oi_1 _06170_ (.A1(_00188_),
    .A2(_00503_),
    .Y(_00002_),
    .B1(_00517_));
 sg13g2_nand2_2 _06171_ (.Y(_00518_),
    .A(_00494_),
    .B(_00502_));
 sg13g2_nand2_2 _06172_ (.Y(_00519_),
    .A(_00494_),
    .B(_00503_));
 sg13g2_nor2b_1 _06173_ (.A(_00519_),
    .B_N(_00516_),
    .Y(_00520_));
 sg13g2_nand3_1 _06174_ (.B(_00503_),
    .C(_00516_),
    .A(_00494_),
    .Y(_00521_));
 sg13g2_nand2_1 _06175_ (.Y(_00522_),
    .A(_00185_),
    .B(_00184_));
 sg13g2_inv_1 _06176_ (.Y(_00523_),
    .A(_00522_));
 sg13g2_o21ai_1 _06177_ (.B1(_00504_),
    .Y(_00524_),
    .A1(_00518_),
    .A2(_00522_));
 sg13g2_nand2b_1 _06178_ (.Y(_00003_),
    .B(_00521_),
    .A_N(_00524_));
 sg13g2_o21ai_1 _06179_ (.B1(_00184_),
    .Y(_00525_),
    .A1(net1736),
    .A2(_00509_));
 sg13g2_xnor2_1 _06180_ (.Y(_00526_),
    .A(_00186_),
    .B(_00525_));
 sg13g2_o21ai_1 _06181_ (.B1(_00504_),
    .Y(_00004_),
    .A1(_00518_),
    .A2(_00526_));
 sg13g2_o21ai_1 _06182_ (.B1(_00504_),
    .Y(_00005_),
    .A1(_00521_),
    .A2(_00523_));
 sg13g2_or2_1 _06183_ (.X(_00527_),
    .B(_00516_),
    .A(_00505_));
 sg13g2_o21ai_1 _06184_ (.B1(_00504_),
    .Y(_00000_),
    .A1(_00516_),
    .A2(_00519_));
 sg13g2_nand2_1 _06185_ (.Y(_00528_),
    .A(_00498_),
    .B(_00501_));
 sg13g2_nor2_1 _06186_ (.A(_00185_),
    .B(_00519_),
    .Y(_00116_));
 sg13g2_nor2_1 _06187_ (.A(_05637_),
    .B(_00438_),
    .Y(_00017_));
 sg13g2_nor2_1 _06188_ (.A(_05634_),
    .B(_00438_),
    .Y(_00016_));
 sg13g2_nor2_1 _06189_ (.A(_05607_),
    .B(_00438_),
    .Y(_00018_));
 sg13g2_nor2_1 _06190_ (.A(net1254),
    .B(_00438_),
    .Y(_00009_));
 sg13g2_nor2_1 _06191_ (.A(_00429_),
    .B(_00438_),
    .Y(_00011_));
 sg13g2_nor2_1 _06192_ (.A(_05640_),
    .B(_00438_),
    .Y(_00008_));
 sg13g2_nor2_1 _06193_ (.A(_05645_),
    .B(_00438_),
    .Y(_00010_));
 sg13g2_or2_1 _06194_ (.X(_00529_),
    .B(_00184_),
    .A(_00509_));
 sg13g2_or2_1 _06195_ (.X(_00530_),
    .B(_00529_),
    .A(_00505_));
 sg13g2_nor3_2 _06196_ (.A(net1464),
    .B(\byte_counter[3] ),
    .C(_00422_),
    .Y(_00531_));
 sg13g2_nand2_1 _06197_ (.Y(_00532_),
    .A(_00453_),
    .B(net1320));
 sg13g2_mux2_1 _06198_ (.A0(net1),
    .A1(net1733),
    .S(net1250),
    .X(_00031_));
 sg13g2_nor2_1 _06199_ (.A(net2),
    .B(net1249),
    .Y(_00533_));
 sg13g2_a21oi_1 _06200_ (.A1(_05569_),
    .A2(net1250),
    .Y(_00032_),
    .B1(_00533_));
 sg13g2_mux2_1 _06201_ (.A0(net3),
    .A1(net1720),
    .S(net1250),
    .X(_00033_));
 sg13g2_nor2_1 _06202_ (.A(net4),
    .B(net1249),
    .Y(_00534_));
 sg13g2_a21oi_1 _06203_ (.A1(_05568_),
    .A2(net1249),
    .Y(_00034_),
    .B1(_00534_));
 sg13g2_nor2_1 _06204_ (.A(net5),
    .B(net1249),
    .Y(_00535_));
 sg13g2_a21oi_1 _06205_ (.A1(_05567_),
    .A2(net1249),
    .Y(_00035_),
    .B1(_00535_));
 sg13g2_nor2_1 _06206_ (.A(net6),
    .B(net1249),
    .Y(_00536_));
 sg13g2_a21oi_1 _06207_ (.A1(_05566_),
    .A2(net1249),
    .Y(_00036_),
    .B1(_00536_));
 sg13g2_mux2_1 _06208_ (.A0(net7),
    .A1(net1698),
    .S(net1250),
    .X(_00037_));
 sg13g2_nor2_1 _06209_ (.A(net8),
    .B(net1249),
    .Y(_00537_));
 sg13g2_a21oi_1 _06210_ (.A1(_05565_),
    .A2(net1250),
    .Y(_00038_),
    .B1(_00537_));
 sg13g2_nor2_1 _06211_ (.A(net1),
    .B(net1252),
    .Y(_00538_));
 sg13g2_a21oi_1 _06212_ (.A1(_05564_),
    .A2(net1252),
    .Y(_00039_),
    .B1(_00538_));
 sg13g2_nor2_1 _06213_ (.A(net2),
    .B(net1251),
    .Y(_00539_));
 sg13g2_a21oi_1 _06214_ (.A1(_05563_),
    .A2(net1251),
    .Y(_00040_),
    .B1(_00539_));
 sg13g2_mux2_1 _06215_ (.A0(net3),
    .A1(net1674),
    .S(_00454_),
    .X(_00041_));
 sg13g2_nor2_1 _06216_ (.A(net4),
    .B(net1251),
    .Y(_00540_));
 sg13g2_a21oi_1 _06217_ (.A1(_05562_),
    .A2(net1251),
    .Y(_00042_),
    .B1(_00540_));
 sg13g2_mux2_1 _06218_ (.A0(net5),
    .A1(net1666),
    .S(net1252),
    .X(_00043_));
 sg13g2_nor2_1 _06219_ (.A(net6),
    .B(net1251),
    .Y(_00541_));
 sg13g2_a21oi_1 _06220_ (.A1(_05561_),
    .A2(net1251),
    .Y(_00044_),
    .B1(_00541_));
 sg13g2_mux2_1 _06221_ (.A0(net7),
    .A1(net1658),
    .S(net1252),
    .X(_00045_));
 sg13g2_nor2_1 _06222_ (.A(net8),
    .B(net1251),
    .Y(_00542_));
 sg13g2_a21oi_1 _06223_ (.A1(_05560_),
    .A2(net1251),
    .Y(_00046_),
    .B1(_00542_));
 sg13g2_nand2_1 _06224_ (.Y(_00543_),
    .A(net724),
    .B(net1382));
 sg13g2_nand3_1 _06225_ (.B(net1382),
    .C(_05624_),
    .A(net761),
    .Y(_00544_));
 sg13g2_nor4_2 _06226_ (.A(\byte_counter[1] ),
    .B(net1465),
    .C(net1464),
    .Y(_00545_),
    .D(\byte_counter[3] ));
 sg13g2_nor2b_2 _06227_ (.A(_00544_),
    .B_N(net1347),
    .Y(_00546_));
 sg13g2_nand2_1 _06228_ (.Y(_00547_),
    .A(net1),
    .B(net1278));
 sg13g2_o21ai_1 _06229_ (.B1(_00547_),
    .Y(_00047_),
    .A1(_05559_),
    .A2(net1278));
 sg13g2_mux2_1 _06230_ (.A0(net1633),
    .A1(net2),
    .S(net1279),
    .X(_00048_));
 sg13g2_nand2_1 _06231_ (.Y(_00548_),
    .A(net3),
    .B(net1278));
 sg13g2_o21ai_1 _06232_ (.B1(_00548_),
    .Y(_00049_),
    .A1(_05558_),
    .A2(net1278));
 sg13g2_mux2_1 _06233_ (.A0(net1627),
    .A1(net4),
    .S(net1279),
    .X(_00050_));
 sg13g2_nand2_1 _06234_ (.Y(_00549_),
    .A(net5),
    .B(net1278));
 sg13g2_o21ai_1 _06235_ (.B1(_00549_),
    .Y(_00051_),
    .A1(_05557_),
    .A2(net1278));
 sg13g2_mux2_1 _06236_ (.A0(net1615),
    .A1(net6),
    .S(net1279),
    .X(_00052_));
 sg13g2_mux2_1 _06237_ (.A0(net1611),
    .A1(net7),
    .S(net1279),
    .X(_00053_));
 sg13g2_nand2_1 _06238_ (.Y(_00550_),
    .A(net8),
    .B(net1278));
 sg13g2_o21ai_1 _06239_ (.B1(_00550_),
    .Y(_00054_),
    .A1(_05556_),
    .A2(net1278));
 sg13g2_nor4_2 _06240_ (.A(net1464),
    .B(net772),
    .C(_00422_),
    .Y(_00551_),
    .D(_00544_));
 sg13g2_mux2_1 _06241_ (.A0(net1601),
    .A1(net1),
    .S(net1277),
    .X(_00055_));
 sg13g2_mux2_1 _06242_ (.A0(net1596),
    .A1(net2),
    .S(net1277),
    .X(_00056_));
 sg13g2_mux2_1 _06243_ (.A0(net1589),
    .A1(net3),
    .S(net1277),
    .X(_00057_));
 sg13g2_mux2_1 _06244_ (.A0(net1582),
    .A1(net4),
    .S(net1277),
    .X(_00058_));
 sg13g2_mux2_1 _06245_ (.A0(net1576),
    .A1(net5),
    .S(net1277),
    .X(_00059_));
 sg13g2_mux2_1 _06246_ (.A0(net1572),
    .A1(net6),
    .S(net1277),
    .X(_00060_));
 sg13g2_nand2_1 _06247_ (.Y(_00552_),
    .A(net7),
    .B(net1277));
 sg13g2_o21ai_1 _06248_ (.B1(_00552_),
    .Y(_00061_),
    .A1(_05555_),
    .A2(net1277));
 sg13g2_mux2_1 _06249_ (.A0(net1564),
    .A1(net8),
    .S(_00551_),
    .X(_00062_));
 sg13g2_and2_1 _06250_ (.A(\cordic_inst.cordic_state[32] ),
    .B(net1255),
    .X(_00553_));
 sg13g2_a21oi_1 _06251_ (.A1(\cordic_inst.get_normalize[24] ),
    .A2(net1261),
    .Y(_00554_),
    .B1(_00553_));
 sg13g2_a21oi_1 _06252_ (.A1(_00028_),
    .A2(_00436_),
    .Y(_00555_),
    .B1(net1254));
 sg13g2_nand2b_1 _06253_ (.Y(_00556_),
    .B(_05600_),
    .A_N(_00555_));
 sg13g2_nor2_1 _06254_ (.A(_05629_),
    .B(_05645_),
    .Y(_00557_));
 sg13g2_o21ai_1 _06255_ (.B1(_05658_),
    .Y(_00558_),
    .A1(_05650_),
    .A2(net1254));
 sg13g2_or4_1 _06256_ (.A(_00420_),
    .B(_00556_),
    .C(_00557_),
    .D(_00558_),
    .X(_00559_));
 sg13g2_nand2_1 _06257_ (.Y(_00560_),
    .A(net350),
    .B(net1218));
 sg13g2_o21ai_1 _06258_ (.B1(_00560_),
    .Y(_00063_),
    .A1(_00554_),
    .A2(net1218));
 sg13g2_and2_1 _06259_ (.A(\cordic_inst.cordic_state[33] ),
    .B(net1256),
    .X(_00561_));
 sg13g2_a21oi_1 _06260_ (.A1(\cordic_inst.get_normalize[25] ),
    .A2(net1262),
    .Y(_00562_),
    .B1(_00561_));
 sg13g2_nand2_1 _06261_ (.Y(_00563_),
    .A(net340),
    .B(net1220));
 sg13g2_o21ai_1 _06262_ (.B1(_00563_),
    .Y(_00064_),
    .A1(net1220),
    .A2(_00562_));
 sg13g2_and2_1 _06263_ (.A(\cordic_inst.cordic_state[34] ),
    .B(net1255),
    .X(_00564_));
 sg13g2_a21oi_1 _06264_ (.A1(\cordic_inst.get_normalize[26] ),
    .A2(net1265),
    .Y(_00565_),
    .B1(_00564_));
 sg13g2_nand2_1 _06265_ (.Y(_00566_),
    .A(net292),
    .B(net1216));
 sg13g2_o21ai_1 _06266_ (.B1(_00566_),
    .Y(_00065_),
    .A1(net1217),
    .A2(_00565_));
 sg13g2_nor2_1 _06267_ (.A(_05584_),
    .B(net1259),
    .Y(_00567_));
 sg13g2_a21oi_1 _06268_ (.A1(\cordic_inst.get_normalize[27] ),
    .A2(net1259),
    .Y(_00568_),
    .B1(_00567_));
 sg13g2_nand2_1 _06269_ (.Y(_00569_),
    .A(net300),
    .B(net1214));
 sg13g2_o21ai_1 _06270_ (.B1(_00569_),
    .Y(_00066_),
    .A1(net1214),
    .A2(_00568_));
 sg13g2_and2_1 _06271_ (.A(\cordic_inst.cordic_state[36] ),
    .B(net1255),
    .X(_00570_));
 sg13g2_a21oi_1 _06272_ (.A1(\cordic_inst.get_normalize[28] ),
    .A2(net1262),
    .Y(_00571_),
    .B1(_00570_));
 sg13g2_nand2_1 _06273_ (.Y(_00572_),
    .A(net302),
    .B(net1220));
 sg13g2_o21ai_1 _06274_ (.B1(_00572_),
    .Y(_00067_),
    .A1(net1220),
    .A2(_00571_));
 sg13g2_and2_1 _06275_ (.A(net1426),
    .B(net1253),
    .X(_00573_));
 sg13g2_a21oi_1 _06276_ (.A1(\cordic_inst.get_normalize[29] ),
    .A2(net1259),
    .Y(_00574_),
    .B1(_00573_));
 sg13g2_nand2_1 _06277_ (.Y(_00575_),
    .A(net282),
    .B(net1213));
 sg13g2_o21ai_1 _06278_ (.B1(_00575_),
    .Y(_00068_),
    .A1(net1213),
    .A2(_00574_));
 sg13g2_and2_1 _06279_ (.A(net1425),
    .B(net1254),
    .X(_00576_));
 sg13g2_a21oi_1 _06280_ (.A1(\cordic_inst.get_normalize[30] ),
    .A2(net1259),
    .Y(_00577_),
    .B1(_00576_));
 sg13g2_nand2_1 _06281_ (.Y(_00578_),
    .A(net324),
    .B(net1220));
 sg13g2_o21ai_1 _06282_ (.B1(_00578_),
    .Y(_00069_),
    .A1(net1218),
    .A2(_00577_));
 sg13g2_and2_1 _06283_ (.A(\cordic_inst.cordic_state[39] ),
    .B(net1255),
    .X(_00579_));
 sg13g2_a21oi_1 _06284_ (.A1(\cordic_inst.get_normalize[31] ),
    .A2(net1261),
    .Y(_00580_),
    .B1(_00579_));
 sg13g2_nand2_1 _06285_ (.Y(_00581_),
    .A(net410),
    .B(net1218));
 sg13g2_o21ai_1 _06286_ (.B1(_00581_),
    .Y(_00070_),
    .A1(net1218),
    .A2(_00580_));
 sg13g2_and2_1 _06287_ (.A(net1423),
    .B(net1253),
    .X(_00582_));
 sg13g2_a21oi_1 _06288_ (.A1(net414),
    .A2(net1257),
    .Y(_00583_),
    .B1(_00582_));
 sg13g2_nand2_1 _06289_ (.Y(_00584_),
    .A(net524),
    .B(net1211));
 sg13g2_o21ai_1 _06290_ (.B1(_00584_),
    .Y(_00071_),
    .A1(net1211),
    .A2(_00583_));
 sg13g2_and2_1 _06291_ (.A(net1422),
    .B(net1254),
    .X(_00585_));
 sg13g2_a21oi_1 _06292_ (.A1(\cordic_inst.get_normalize[33] ),
    .A2(net1257),
    .Y(_00586_),
    .B1(_00585_));
 sg13g2_nand2_1 _06293_ (.Y(_00587_),
    .A(net478),
    .B(net1211));
 sg13g2_o21ai_1 _06294_ (.B1(_00587_),
    .Y(_00072_),
    .A1(net1211),
    .A2(_00586_));
 sg13g2_and2_1 _06295_ (.A(net1421),
    .B(net1253),
    .X(_00588_));
 sg13g2_a21oi_1 _06296_ (.A1(net449),
    .A2(net1257),
    .Y(_00589_),
    .B1(_00588_));
 sg13g2_nand2_1 _06297_ (.Y(_00590_),
    .A(net532),
    .B(net1210));
 sg13g2_o21ai_1 _06298_ (.B1(_00590_),
    .Y(_00073_),
    .A1(net1210),
    .A2(_00589_));
 sg13g2_and2_1 _06299_ (.A(\cordic_inst.cordic_state[43] ),
    .B(net1253),
    .X(_00591_));
 sg13g2_a21oi_1 _06300_ (.A1(\cordic_inst.get_normalize[35] ),
    .A2(net1258),
    .Y(_00592_),
    .B1(_00591_));
 sg13g2_nand2_1 _06301_ (.Y(_00593_),
    .A(net402),
    .B(net1215));
 sg13g2_o21ai_1 _06302_ (.B1(_00593_),
    .Y(_00074_),
    .A1(net1215),
    .A2(_00592_));
 sg13g2_and2_1 _06303_ (.A(\cordic_inst.cordic_state[44] ),
    .B(net1253),
    .X(_00594_));
 sg13g2_a21oi_1 _06304_ (.A1(net464),
    .A2(net1257),
    .Y(_00595_),
    .B1(_00594_));
 sg13g2_nand2_1 _06305_ (.Y(_00596_),
    .A(net504),
    .B(net1210));
 sg13g2_o21ai_1 _06306_ (.B1(_00596_),
    .Y(_00075_),
    .A1(net1210),
    .A2(_00595_));
 sg13g2_and2_1 _06307_ (.A(\cordic_inst.cordic_state[45] ),
    .B(net1256),
    .X(_00597_));
 sg13g2_a21oi_1 _06308_ (.A1(\cordic_inst.get_normalize[37] ),
    .A2(net1257),
    .Y(_00598_),
    .B1(_00597_));
 sg13g2_nand2_1 _06309_ (.Y(_00599_),
    .A(net431),
    .B(net1210));
 sg13g2_o21ai_1 _06310_ (.B1(_00599_),
    .Y(_00076_),
    .A1(net1210),
    .A2(_00598_));
 sg13g2_and2_1 _06311_ (.A(\cordic_inst.cordic_state[46] ),
    .B(net1253),
    .X(_00600_));
 sg13g2_a21oi_1 _06312_ (.A1(net391),
    .A2(net1258),
    .Y(_00601_),
    .B1(_00600_));
 sg13g2_nand2_1 _06313_ (.Y(_00602_),
    .A(net451),
    .B(net1210));
 sg13g2_o21ai_1 _06314_ (.B1(_00602_),
    .Y(_00077_),
    .A1(net1210),
    .A2(_00601_));
 sg13g2_and2_1 _06315_ (.A(net1416),
    .B(net1253),
    .X(_00603_));
 sg13g2_a21oi_1 _06316_ (.A1(\cordic_inst.get_normalize[39] ),
    .A2(net1259),
    .Y(_00604_),
    .B1(_00603_));
 sg13g2_nand2_1 _06317_ (.Y(_00605_),
    .A(net389),
    .B(net1214));
 sg13g2_o21ai_1 _06318_ (.B1(_00605_),
    .Y(_00078_),
    .A1(net1214),
    .A2(_00604_));
 sg13g2_and2_1 _06319_ (.A(net1415),
    .B(net1253),
    .X(_00606_));
 sg13g2_a21oi_1 _06320_ (.A1(net513),
    .A2(net1258),
    .Y(_00607_),
    .B1(_00606_));
 sg13g2_nand2_1 _06321_ (.Y(_00608_),
    .A(net530),
    .B(net1212));
 sg13g2_o21ai_1 _06322_ (.B1(_00608_),
    .Y(_00079_),
    .A1(net1211),
    .A2(_00607_));
 sg13g2_nor2_2 _06323_ (.A(_05583_),
    .B(net1258),
    .Y(_00609_));
 sg13g2_a21oi_1 _06324_ (.A1(\cordic_inst.get_normalize[41] ),
    .A2(net1261),
    .Y(_00610_),
    .B1(_00609_));
 sg13g2_nand2_1 _06325_ (.Y(_00611_),
    .A(net316),
    .B(net1224));
 sg13g2_o21ai_1 _06326_ (.B1(_00611_),
    .Y(_00080_),
    .A1(net1216),
    .A2(_00610_));
 sg13g2_and2_1 _06327_ (.A(net1414),
    .B(net1254),
    .X(_00612_));
 sg13g2_a21oi_1 _06328_ (.A1(\cordic_inst.get_normalize[42] ),
    .A2(net1257),
    .Y(_00613_),
    .B1(_00612_));
 sg13g2_nand2_1 _06329_ (.Y(_00614_),
    .A(net320),
    .B(net1212));
 sg13g2_o21ai_1 _06330_ (.B1(_00614_),
    .Y(_00081_),
    .A1(net1212),
    .A2(_00613_));
 sg13g2_nor2_1 _06331_ (.A(_05582_),
    .B(net1259),
    .Y(_00615_));
 sg13g2_a21oi_1 _06332_ (.A1(\cordic_inst.get_normalize[43] ),
    .A2(net1259),
    .Y(_00616_),
    .B1(_00615_));
 sg13g2_nand2_1 _06333_ (.Y(_00617_),
    .A(net344),
    .B(net1214));
 sg13g2_o21ai_1 _06334_ (.B1(_00617_),
    .Y(_00082_),
    .A1(net1214),
    .A2(_00616_));
 sg13g2_and2_1 _06335_ (.A(net1413),
    .B(net1255),
    .X(_00618_));
 sg13g2_a21oi_1 _06336_ (.A1(\cordic_inst.get_normalize[44] ),
    .A2(net1263),
    .Y(_00619_),
    .B1(_00618_));
 sg13g2_nand2_1 _06337_ (.Y(_00620_),
    .A(net381),
    .B(net1221));
 sg13g2_o21ai_1 _06338_ (.B1(_00620_),
    .Y(_00083_),
    .A1(net1221),
    .A2(_00619_));
 sg13g2_and2_1 _06339_ (.A(net1412),
    .B(net1255),
    .X(_00621_));
 sg13g2_a21oi_1 _06340_ (.A1(net470),
    .A2(net1263),
    .Y(_00622_),
    .B1(_00621_));
 sg13g2_nand2_1 _06341_ (.Y(_00623_),
    .A(net480),
    .B(net1219));
 sg13g2_o21ai_1 _06342_ (.B1(_00623_),
    .Y(_00084_),
    .A1(net1219),
    .A2(_00622_));
 sg13g2_and2_1 _06343_ (.A(\cordic_inst.cordic_state[54] ),
    .B(net1255),
    .X(_00624_));
 sg13g2_a21oi_1 _06344_ (.A1(\cordic_inst.get_normalize[46] ),
    .A2(net1262),
    .Y(_00625_),
    .B1(_00624_));
 sg13g2_nand2_1 _06345_ (.Y(_00626_),
    .A(net332),
    .B(net1219));
 sg13g2_o21ai_1 _06346_ (.B1(_00626_),
    .Y(_00085_),
    .A1(net1219),
    .A2(_00625_));
 sg13g2_and2_1 _06347_ (.A(net1410),
    .B(net1255),
    .X(_00627_));
 sg13g2_a21oi_1 _06348_ (.A1(\cordic_inst.get_normalize[47] ),
    .A2(net1262),
    .Y(_00628_),
    .B1(_00627_));
 sg13g2_nand2_1 _06349_ (.Y(_00629_),
    .A(net360),
    .B(net1219));
 sg13g2_o21ai_1 _06350_ (.B1(_00629_),
    .Y(_00086_),
    .A1(net1219),
    .A2(_00628_));
 sg13g2_nand2_1 _06351_ (.Y(_00630_),
    .A(net418),
    .B(net1261));
 sg13g2_nand2_1 _06352_ (.Y(_00631_),
    .A(\result_reg[48] ),
    .B(net1217));
 sg13g2_o21ai_1 _06353_ (.B1(_00631_),
    .Y(_00087_),
    .A1(net1217),
    .A2(_00630_));
 sg13g2_nand2_1 _06354_ (.Y(_00632_),
    .A(\cordic_inst.get_normalize[49] ),
    .B(net1264));
 sg13g2_nand2_1 _06355_ (.Y(_00633_),
    .A(net395),
    .B(net1224));
 sg13g2_o21ai_1 _06356_ (.B1(_00633_),
    .Y(_00088_),
    .A1(net1224),
    .A2(_00632_));
 sg13g2_nand2_1 _06357_ (.Y(_00634_),
    .A(net290),
    .B(net1216));
 sg13g2_nand2_1 _06358_ (.Y(_00635_),
    .A(\cordic_inst.get_normalize[50] ),
    .B(net1261));
 sg13g2_o21ai_1 _06359_ (.B1(_00634_),
    .Y(_00089_),
    .A1(net1216),
    .A2(_00635_));
 sg13g2_nand2_1 _06360_ (.Y(_00636_),
    .A(\result_reg[51] ),
    .B(net1217));
 sg13g2_nand2_1 _06361_ (.Y(_00637_),
    .A(net466),
    .B(net1261));
 sg13g2_o21ai_1 _06362_ (.B1(_00636_),
    .Y(_00090_),
    .A1(net1217),
    .A2(_00637_));
 sg13g2_nand2_1 _06363_ (.Y(_00638_),
    .A(net434),
    .B(net1264));
 sg13g2_nand2_1 _06364_ (.Y(_00639_),
    .A(net498),
    .B(net1225));
 sg13g2_o21ai_1 _06365_ (.B1(_00639_),
    .Y(_00091_),
    .A1(net1225),
    .A2(_00638_));
 sg13g2_nand2_1 _06366_ (.Y(_00640_),
    .A(net288),
    .B(net1213));
 sg13g2_nand2_1 _06367_ (.Y(_00641_),
    .A(\cordic_inst.get_normalize[53] ),
    .B(net1260));
 sg13g2_o21ai_1 _06368_ (.B1(_00640_),
    .Y(_00092_),
    .A1(net1213),
    .A2(_00641_));
 sg13g2_nand2_1 _06369_ (.Y(_00642_),
    .A(\cordic_inst.get_normalize[54] ),
    .B(net1260));
 sg13g2_nand2_1 _06370_ (.Y(_00643_),
    .A(net330),
    .B(net1213));
 sg13g2_o21ai_1 _06371_ (.B1(_00643_),
    .Y(_00093_),
    .A1(net1212),
    .A2(_00642_));
 sg13g2_nand2_1 _06372_ (.Y(_00644_),
    .A(\cordic_inst.get_normalize[55] ),
    .B(net1264));
 sg13g2_nand2_1 _06373_ (.Y(_00645_),
    .A(net322),
    .B(net1224));
 sg13g2_o21ai_1 _06374_ (.B1(_00645_),
    .Y(_00094_),
    .A1(net1224),
    .A2(_00644_));
 sg13g2_nand2_1 _06375_ (.Y(_00646_),
    .A(net453),
    .B(net1257));
 sg13g2_nand2_1 _06376_ (.Y(_00647_),
    .A(net491),
    .B(net1212));
 sg13g2_o21ai_1 _06377_ (.B1(_00647_),
    .Y(_00095_),
    .A1(net1212),
    .A2(_00646_));
 sg13g2_nand2_1 _06378_ (.Y(_00648_),
    .A(\result_reg[57] ),
    .B(net1216));
 sg13g2_nand2_1 _06379_ (.Y(_00649_),
    .A(net383),
    .B(net1261));
 sg13g2_o21ai_1 _06380_ (.B1(_00648_),
    .Y(_00096_),
    .A1(net1216),
    .A2(_00649_));
 sg13g2_nand2_1 _06381_ (.Y(_00650_),
    .A(net459),
    .B(net1261));
 sg13g2_nand2_1 _06382_ (.Y(_00651_),
    .A(net509),
    .B(net1216));
 sg13g2_o21ai_1 _06383_ (.B1(_00651_),
    .Y(_00097_),
    .A1(net1216),
    .A2(_00650_));
 sg13g2_nand2_1 _06384_ (.Y(_00652_),
    .A(net348),
    .B(net1212));
 sg13g2_nand2_1 _06385_ (.Y(_00653_),
    .A(\cordic_inst.get_normalize[59] ),
    .B(net1257));
 sg13g2_o21ai_1 _06386_ (.B1(_00652_),
    .Y(_00098_),
    .A1(net1212),
    .A2(_00653_));
 sg13g2_nand2_1 _06387_ (.Y(_00654_),
    .A(\cordic_inst.get_normalize[60] ),
    .B(net1260));
 sg13g2_nand2_1 _06388_ (.Y(_00655_),
    .A(net308),
    .B(net1213));
 sg13g2_o21ai_1 _06389_ (.B1(_00655_),
    .Y(_00099_),
    .A1(net1213),
    .A2(_00654_));
 sg13g2_nand2_1 _06390_ (.Y(_00656_),
    .A(\cordic_inst.get_normalize[61] ),
    .B(net1264));
 sg13g2_nand2_1 _06391_ (.Y(_00657_),
    .A(net346),
    .B(net1224));
 sg13g2_o21ai_1 _06392_ (.B1(_00657_),
    .Y(_00100_),
    .A1(net1225),
    .A2(_00656_));
 sg13g2_nand2_1 _06393_ (.Y(_00658_),
    .A(net540),
    .B(net1225));
 sg13g2_nand2_1 _06394_ (.Y(_00659_),
    .A(net358),
    .B(net1264));
 sg13g2_o21ai_1 _06395_ (.B1(_00658_),
    .Y(_00101_),
    .A1(net1225),
    .A2(_00659_));
 sg13g2_nand2_1 _06396_ (.Y(_00660_),
    .A(\result_reg[63] ),
    .B(net1225));
 sg13g2_nand2_1 _06397_ (.Y(_00661_),
    .A(net363),
    .B(net1264));
 sg13g2_o21ai_1 _06398_ (.B1(_00660_),
    .Y(_00102_),
    .A1(net1225),
    .A2(_00661_));
 sg13g2_nand2_1 _06399_ (.Y(_00662_),
    .A(net393),
    .B(net1224));
 sg13g2_nand2_1 _06400_ (.Y(_00663_),
    .A(\cordic_inst.get_normalize[64] ),
    .B(net1265));
 sg13g2_o21ai_1 _06401_ (.B1(_00662_),
    .Y(_00103_),
    .A1(net1224),
    .A2(_00663_));
 sg13g2_nand2_1 _06402_ (.Y(_00664_),
    .A(\cordic_inst.get_normalize[65] ),
    .B(net1263));
 sg13g2_nand2_1 _06403_ (.Y(_00665_),
    .A(net440),
    .B(net1222));
 sg13g2_o21ai_1 _06404_ (.B1(_00665_),
    .Y(_00104_),
    .A1(net1222),
    .A2(_00664_));
 sg13g2_nand2_1 _06405_ (.Y(_00666_),
    .A(net486),
    .B(net1222));
 sg13g2_nand2_1 _06406_ (.Y(_00667_),
    .A(net399),
    .B(net1263));
 sg13g2_o21ai_1 _06407_ (.B1(_00666_),
    .Y(_00105_),
    .A1(net1222),
    .A2(_00667_));
 sg13g2_nand2_1 _06408_ (.Y(_00668_),
    .A(net284),
    .B(net1214));
 sg13g2_nand2_1 _06409_ (.Y(_00669_),
    .A(\cordic_inst.get_normalize[67] ),
    .B(net1259));
 sg13g2_o21ai_1 _06410_ (.B1(_00668_),
    .Y(_00106_),
    .A1(net1214),
    .A2(_00669_));
 sg13g2_nand2_1 _06411_ (.Y(_00670_),
    .A(net326),
    .B(net1219));
 sg13g2_nand2_1 _06412_ (.Y(_00671_),
    .A(\cordic_inst.get_normalize[68] ),
    .B(net1262));
 sg13g2_o21ai_1 _06413_ (.B1(_00670_),
    .Y(_00107_),
    .A1(net1219),
    .A2(_00671_));
 sg13g2_nand2_1 _06414_ (.Y(_00672_),
    .A(net474),
    .B(net1262));
 sg13g2_nand2_1 _06415_ (.Y(_00673_),
    .A(\result_reg[69] ),
    .B(net1221));
 sg13g2_o21ai_1 _06416_ (.B1(_00673_),
    .Y(_00108_),
    .A1(net1221),
    .A2(_00672_));
 sg13g2_nand2_1 _06417_ (.Y(_00674_),
    .A(net507),
    .B(net1262));
 sg13g2_nand2_1 _06418_ (.Y(_00675_),
    .A(net526),
    .B(net1221));
 sg13g2_o21ai_1 _06419_ (.B1(_00675_),
    .Y(_00109_),
    .A1(net1221),
    .A2(_00674_));
 sg13g2_nand2_1 _06420_ (.Y(_00676_),
    .A(net379),
    .B(net1262));
 sg13g2_nand2_1 _06421_ (.Y(_00677_),
    .A(\result_reg[71] ),
    .B(net1221));
 sg13g2_o21ai_1 _06422_ (.B1(_00677_),
    .Y(_00110_),
    .A1(net1221),
    .A2(_00676_));
 sg13g2_a21oi_1 _06423_ (.A1(_00513_),
    .A2(_00529_),
    .Y(_00111_),
    .B1(_00518_));
 sg13g2_nor3_1 _06424_ (.A(_00498_),
    .B(_00516_),
    .C(_00518_),
    .Y(_00117_));
 sg13g2_or2_1 _06425_ (.X(_00112_),
    .B(_00117_),
    .A(_00520_));
 sg13g2_nand3_1 _06426_ (.B(_00528_),
    .C(_00529_),
    .A(_00494_),
    .Y(_00678_));
 sg13g2_a21oi_1 _06427_ (.A1(_00186_),
    .A2(_00515_),
    .Y(_00113_),
    .B1(_00678_));
 sg13g2_nand2_1 _06428_ (.Y(_00114_),
    .A(_00521_),
    .B(_00530_));
 sg13g2_o21ai_1 _06429_ (.B1(_00527_),
    .Y(_00115_),
    .A1(_00519_),
    .A2(_00522_));
 sg13g2_nor2_2 _06430_ (.A(_05618_),
    .B(_00440_),
    .Y(_00679_));
 sg13g2_nand2_1 _06431_ (.Y(_00680_),
    .A(\byte_counter[1] ),
    .B(net1465));
 sg13g2_nor3_2 _06432_ (.A(net1464),
    .B(\byte_counter[3] ),
    .C(_00680_),
    .Y(_00681_));
 sg13g2_and2_1 _06433_ (.A(net342),
    .B(net1320),
    .X(_00682_));
 sg13g2_a22oi_1 _06434_ (.Y(_00683_),
    .B1(net1347),
    .B2(net328),
    .A2(net1325),
    .A1(net393));
 sg13g2_nand3_1 _06435_ (.B(net1465),
    .C(net1464),
    .A(\byte_counter[1] ),
    .Y(_00684_));
 sg13g2_nor2_2 _06436_ (.A(\byte_counter[3] ),
    .B(_00684_),
    .Y(_00685_));
 sg13g2_nor2_2 _06437_ (.A(_05626_),
    .B(_00423_),
    .Y(_00686_));
 sg13g2_nor3_2 _06438_ (.A(\byte_counter[1] ),
    .B(net1465),
    .C(_00423_),
    .Y(_00687_));
 sg13g2_a221oi_1 _06439_ (.B2(\result_reg[48] ),
    .C1(_00682_),
    .B1(_00686_),
    .A1(net605),
    .Y(_00688_),
    .A2(net1326));
 sg13g2_a22oi_1 _06440_ (.Y(_00689_),
    .B1(_00687_),
    .B2(net524),
    .A2(_00681_),
    .A1(net350));
 sg13g2_a22oi_1 _06441_ (.Y(_00690_),
    .B1(_00685_),
    .B2(net491),
    .A2(net1306),
    .A1(net530));
 sg13g2_nand4_1 _06442_ (.B(_00688_),
    .C(_00689_),
    .A(_00683_),
    .Y(_00691_),
    .D(_00690_));
 sg13g2_a22oi_1 _06443_ (.Y(_00692_),
    .B1(_00691_),
    .B2(net1307),
    .A2(_00679_),
    .A1(net631));
 sg13g2_inv_1 _06444_ (.Y(_00118_),
    .A(net632));
 sg13g2_a22oi_1 _06445_ (.Y(_00693_),
    .B1(net1347),
    .B2(net334),
    .A2(net1325),
    .A1(net440));
 sg13g2_nand2_1 _06446_ (.Y(_00694_),
    .A(net340),
    .B(_00681_));
 sg13g2_a22oi_1 _06447_ (.Y(_00695_),
    .B1(_00687_),
    .B2(\result_reg[33] ),
    .A2(net1326),
    .A1(\result_reg[17] ));
 sg13g2_a22oi_1 _06448_ (.Y(_00696_),
    .B1(_00686_),
    .B2(net395),
    .A2(net1306),
    .A1(net316));
 sg13g2_a22oi_1 _06449_ (.Y(_00697_),
    .B1(_00685_),
    .B2(\result_reg[57] ),
    .A2(net1320),
    .A1(\result_reg[9] ));
 sg13g2_and2_1 _06450_ (.A(_00695_),
    .B(_00697_),
    .X(_00698_));
 sg13g2_nand4_1 _06451_ (.B(_00694_),
    .C(_00696_),
    .A(_00693_),
    .Y(_00699_),
    .D(_00698_));
 sg13g2_a22oi_1 _06452_ (.Y(_00700_),
    .B1(_00699_),
    .B2(net1307),
    .A2(_00679_),
    .A1(net644));
 sg13g2_inv_1 _06453_ (.Y(_00119_),
    .A(net645));
 sg13g2_a22oi_1 _06454_ (.Y(_00701_),
    .B1(_00687_),
    .B2(net532),
    .A2(net1306),
    .A1(net320));
 sg13g2_a22oi_1 _06455_ (.Y(_00702_),
    .B1(_00686_),
    .B2(net290),
    .A2(_00681_),
    .A1(net292));
 sg13g2_nand2_1 _06456_ (.Y(_00703_),
    .A(net486),
    .B(net1325));
 sg13g2_a22oi_1 _06457_ (.Y(_00704_),
    .B1(net1320),
    .B2(net294),
    .A2(net1327),
    .A1(net298));
 sg13g2_nand2_1 _06458_ (.Y(_00705_),
    .A(_00703_),
    .B(_00704_));
 sg13g2_a221oi_1 _06459_ (.B2(net509),
    .C1(_00705_),
    .B1(_00685_),
    .A1(net385),
    .Y(_00706_),
    .A2(net1347));
 sg13g2_nand3_1 _06460_ (.B(_00702_),
    .C(_00706_),
    .A(_00701_),
    .Y(_00707_));
 sg13g2_a22oi_1 _06461_ (.Y(_00708_),
    .B1(_00707_),
    .B2(net1307),
    .A2(_00679_),
    .A1(net647));
 sg13g2_inv_1 _06462_ (.Y(_00120_),
    .A(net648));
 sg13g2_a22oi_1 _06463_ (.Y(_00709_),
    .B1(_00686_),
    .B2(\result_reg[51] ),
    .A2(net1320),
    .A1(net296));
 sg13g2_a22oi_1 _06464_ (.Y(_00710_),
    .B1(_00687_),
    .B2(\result_reg[35] ),
    .A2(_00681_),
    .A1(\result_reg[27] ));
 sg13g2_and2_1 _06465_ (.A(_00709_),
    .B(_00710_),
    .X(_00711_));
 sg13g2_a22oi_1 _06466_ (.Y(_00712_),
    .B1(net1347),
    .B2(net312),
    .A2(net1325),
    .A1(net284));
 sg13g2_nand2_1 _06467_ (.Y(_00713_),
    .A(net348),
    .B(_00685_));
 sg13g2_a22oi_1 _06468_ (.Y(_00714_),
    .B1(net1306),
    .B2(net344),
    .A2(net1326),
    .A1(net338));
 sg13g2_nand4_1 _06469_ (.B(_00712_),
    .C(_00713_),
    .A(_00711_),
    .Y(_00715_),
    .D(_00714_));
 sg13g2_a22oi_1 _06470_ (.Y(_00716_),
    .B1(_00715_),
    .B2(net1307),
    .A2(_00679_),
    .A1(net649));
 sg13g2_inv_1 _06471_ (.Y(_00121_),
    .A(net650));
 sg13g2_a22oi_1 _06472_ (.Y(_00717_),
    .B1(_00686_),
    .B2(\result_reg[52] ),
    .A2(net1327),
    .A1(\result_reg[20] ));
 sg13g2_a22oi_1 _06473_ (.Y(_00718_),
    .B1(_00681_),
    .B2(net302),
    .A2(net1306),
    .A1(\result_reg[44] ));
 sg13g2_and2_1 _06474_ (.A(_00717_),
    .B(_00718_),
    .X(_00719_));
 sg13g2_a22oi_1 _06475_ (.Y(_00720_),
    .B1(net1347),
    .B2(net304),
    .A2(net1325),
    .A1(net326));
 sg13g2_nand2_1 _06476_ (.Y(_00721_),
    .A(net308),
    .B(_00685_));
 sg13g2_a22oi_1 _06477_ (.Y(_00722_),
    .B1(_00687_),
    .B2(net504),
    .A2(net1320),
    .A1(net576));
 sg13g2_nand4_1 _06478_ (.B(_00720_),
    .C(_00721_),
    .A(_00719_),
    .Y(_00723_),
    .D(_00722_));
 sg13g2_a22oi_1 _06479_ (.Y(_00724_),
    .B1(_00723_),
    .B2(_00419_),
    .A2(_00679_),
    .A1(net655));
 sg13g2_inv_1 _06480_ (.Y(_00122_),
    .A(net656));
 sg13g2_nand2_1 _06481_ (.Y(_00725_),
    .A(net282),
    .B(_00681_));
 sg13g2_a22oi_1 _06482_ (.Y(_00726_),
    .B1(_00687_),
    .B2(net431),
    .A2(_00686_),
    .A1(net288));
 sg13g2_a22oi_1 _06483_ (.Y(_00727_),
    .B1(_00531_),
    .B2(net286),
    .A2(net1306),
    .A1(\result_reg[45] ));
 sg13g2_a22oi_1 _06484_ (.Y(_00728_),
    .B1(_00685_),
    .B2(\result_reg[61] ),
    .A2(net1327),
    .A1(\result_reg[21] ));
 sg13g2_nand2_1 _06485_ (.Y(_00729_),
    .A(_00727_),
    .B(_00728_));
 sg13g2_a221oi_1 _06486_ (.B2(net318),
    .C1(_00729_),
    .B1(net1347),
    .A1(\result_reg[69] ),
    .Y(_00730_),
    .A2(net1325));
 sg13g2_nand3_1 _06487_ (.B(_00726_),
    .C(_00730_),
    .A(_00725_),
    .Y(_00731_));
 sg13g2_a22oi_1 _06488_ (.Y(_00732_),
    .B1(_00731_),
    .B2(net1307),
    .A2(_00679_),
    .A1(net636));
 sg13g2_inv_1 _06489_ (.Y(_00123_),
    .A(net637));
 sg13g2_a22oi_1 _06490_ (.Y(_00733_),
    .B1(net1347),
    .B2(net280),
    .A2(net1325),
    .A1(net526));
 sg13g2_nand2_1 _06491_ (.Y(_00734_),
    .A(net566),
    .B(net1320));
 sg13g2_a22oi_1 _06492_ (.Y(_00735_),
    .B1(_00681_),
    .B2(\result_reg[30] ),
    .A2(net1306),
    .A1(\result_reg[46] ));
 sg13g2_a22oi_1 _06493_ (.Y(_00736_),
    .B1(_00687_),
    .B2(net451),
    .A2(_00686_),
    .A1(net330));
 sg13g2_a22oi_1 _06494_ (.Y(_00737_),
    .B1(_00685_),
    .B2(\result_reg[62] ),
    .A2(net1327),
    .A1(\result_reg[22] ));
 sg13g2_and2_1 _06495_ (.A(_00735_),
    .B(_00737_),
    .X(_00738_));
 sg13g2_nand4_1 _06496_ (.B(_00734_),
    .C(_00736_),
    .A(_00733_),
    .Y(_00739_),
    .D(_00738_));
 sg13g2_a22oi_1 _06497_ (.Y(_00740_),
    .B1(_00739_),
    .B2(net1307),
    .A2(_00679_),
    .A1(net641));
 sg13g2_inv_1 _06498_ (.Y(_00124_),
    .A(net642));
 sg13g2_a22oi_1 _06499_ (.Y(_00741_),
    .B1(_00687_),
    .B2(\result_reg[39] ),
    .A2(_00681_),
    .A1(\result_reg[31] ));
 sg13g2_a22oi_1 _06500_ (.Y(_00742_),
    .B1(_00686_),
    .B2(\result_reg[55] ),
    .A2(net1327),
    .A1(\result_reg[23] ));
 sg13g2_and2_1 _06501_ (.A(_00741_),
    .B(_00742_),
    .X(_00743_));
 sg13g2_a22oi_1 _06502_ (.Y(_00744_),
    .B1(net1320),
    .B2(net571),
    .A2(_00424_),
    .A1(net360));
 sg13g2_nand2_1 _06503_ (.Y(_00745_),
    .A(\result_reg[63] ),
    .B(_00685_));
 sg13g2_a22oi_1 _06504_ (.Y(_00746_),
    .B1(_00545_),
    .B2(net306),
    .A2(_00421_),
    .A1(\result_reg[71] ));
 sg13g2_nand4_1 _06505_ (.B(_00744_),
    .C(_00745_),
    .A(_00743_),
    .Y(_00747_),
    .D(_00746_));
 sg13g2_a22oi_1 _06506_ (.Y(_00748_),
    .B1(_00747_),
    .B2(_00419_),
    .A2(_00679_),
    .A1(net754));
 sg13g2_nand2_1 _06507_ (.Y(_00125_),
    .A(_05619_),
    .B(net755));
 sg13g2_nor2_1 _06508_ (.A(net724),
    .B(_00452_),
    .Y(_00749_));
 sg13g2_a21oi_1 _06509_ (.A1(net1382),
    .A2(_00749_),
    .Y(_00750_),
    .B1(_00440_));
 sg13g2_a21oi_1 _06510_ (.A1(_05616_),
    .A2(_00750_),
    .Y(_00751_),
    .B1(_00449_));
 sg13g2_a21o_1 _06511_ (.A2(_00449_),
    .A1(net724),
    .B1(_00751_),
    .X(_00126_));
 sg13g2_a21oi_1 _06512_ (.A1(net1382),
    .A2(_00749_),
    .Y(_00752_),
    .B1(_05622_));
 sg13g2_o21ai_1 _06513_ (.B1(_00450_),
    .Y(_00127_),
    .A1(_00449_),
    .A2(_00752_));
 sg13g2_nor2b_1 _06514_ (.A(_00749_),
    .B_N(net1382),
    .Y(_00753_));
 sg13g2_o21ai_1 _06515_ (.B1(_05616_),
    .Y(_00754_),
    .A1(_05619_),
    .A2(_05621_));
 sg13g2_nor3_1 _06516_ (.A(_00449_),
    .B(_00753_),
    .C(_00754_),
    .Y(_00755_));
 sg13g2_a21oi_1 _06517_ (.A1(_05594_),
    .A2(_00449_),
    .Y(_00128_),
    .B1(_00755_));
 sg13g2_nand2_2 _06518_ (.Y(_00756_),
    .A(_05624_),
    .B(_00440_));
 sg13g2_mux2_1 _06519_ (.A0(net1),
    .A1(net715),
    .S(_00756_),
    .X(_00129_));
 sg13g2_mux2_1 _06520_ (.A0(net2),
    .A1(net693),
    .S(_00756_),
    .X(_00130_));
 sg13g2_mux2_1 _06521_ (.A0(net3),
    .A1(net718),
    .S(_00756_),
    .X(_00131_));
 sg13g2_mux2_1 _06522_ (.A0(net4),
    .A1(net691),
    .S(_00756_),
    .X(_00132_));
 sg13g2_mux2_1 _06523_ (.A0(net5),
    .A1(net625),
    .S(_00756_),
    .X(_00133_));
 sg13g2_mux2_1 _06524_ (.A0(net6),
    .A1(net619),
    .S(_00756_),
    .X(_00134_));
 sg13g2_mux2_1 _06525_ (.A0(net7),
    .A1(net582),
    .S(_00756_),
    .X(_00135_));
 sg13g2_mux2_1 _06526_ (.A0(net8),
    .A1(net568),
    .S(_00756_),
    .X(_00136_));
 sg13g2_nand2_2 _06527_ (.Y(_00757_),
    .A(_05622_),
    .B(_05624_));
 sg13g2_mux2_1 _06528_ (.A0(net1),
    .A1(net1557),
    .S(net1232),
    .X(_00137_));
 sg13g2_nor2_1 _06529_ (.A(net2),
    .B(net1231),
    .Y(_00758_));
 sg13g2_a21oi_1 _06530_ (.A1(_05574_),
    .A2(net1231),
    .Y(_00138_),
    .B1(_00758_));
 sg13g2_nor2_1 _06531_ (.A(net3),
    .B(net1232),
    .Y(_00759_));
 sg13g2_a21oi_1 _06532_ (.A1(_05573_),
    .A2(net1232),
    .Y(_00139_),
    .B1(_00759_));
 sg13g2_nor2_1 _06533_ (.A(net4),
    .B(net1231),
    .Y(_00760_));
 sg13g2_a21oi_1 _06534_ (.A1(_05572_),
    .A2(net1231),
    .Y(_00140_),
    .B1(_00760_));
 sg13g2_mux2_1 _06535_ (.A0(net5),
    .A1(net1531),
    .S(net1232),
    .X(_00141_));
 sg13g2_nor2_1 _06536_ (.A(net6),
    .B(net1231),
    .Y(_00761_));
 sg13g2_a21oi_1 _06537_ (.A1(_05571_),
    .A2(net1231),
    .Y(_00142_),
    .B1(_00761_));
 sg13g2_mux2_1 _06538_ (.A0(net7),
    .A1(net1525),
    .S(net1232),
    .X(_00143_));
 sg13g2_nor2_1 _06539_ (.A(net8),
    .B(net1231),
    .Y(_00762_));
 sg13g2_a21oi_1 _06540_ (.A1(_05570_),
    .A2(net1231),
    .Y(_00144_),
    .B1(_00762_));
 sg13g2_nor2_2 _06541_ (.A(_05628_),
    .B(_00543_),
    .Y(_00763_));
 sg13g2_nand2_1 _06542_ (.Y(_00764_),
    .A(net1),
    .B(net1248));
 sg13g2_o21ai_1 _06543_ (.B1(_00764_),
    .Y(_00145_),
    .A1(_05554_),
    .A2(net1248));
 sg13g2_mux2_1 _06544_ (.A0(net1507),
    .A1(net2),
    .S(net1247),
    .X(_00146_));
 sg13g2_mux2_1 _06545_ (.A0(net1505),
    .A1(net3),
    .S(net1247),
    .X(_00147_));
 sg13g2_mux2_1 _06546_ (.A0(net1501),
    .A1(net4),
    .S(net1247),
    .X(_00148_));
 sg13g2_mux2_1 _06547_ (.A0(net1497),
    .A1(net5),
    .S(net1247),
    .X(_00149_));
 sg13g2_nand2_1 _06548_ (.Y(_00765_),
    .A(net6),
    .B(net1247));
 sg13g2_o21ai_1 _06549_ (.B1(_00765_),
    .Y(_00150_),
    .A1(_05553_),
    .A2(net1247));
 sg13g2_nand2_1 _06550_ (.Y(_00766_),
    .A(net7),
    .B(net1247));
 sg13g2_o21ai_1 _06551_ (.B1(_00766_),
    .Y(_00151_),
    .A1(_05552_),
    .A2(net1247));
 sg13g2_mux2_1 _06552_ (.A0(net1489),
    .A1(net8),
    .S(net1248),
    .X(_00152_));
 sg13g2_or3_1 _06553_ (.A(_00432_),
    .B(_00439_),
    .C(_00007_),
    .X(_00767_));
 sg13g2_and3_1 _06554_ (.X(_00768_),
    .A(_05637_),
    .B(_05645_),
    .C(_00452_));
 sg13g2_a22oi_1 _06555_ (.Y(_00769_),
    .B1(_05647_),
    .B2(_05598_),
    .A2(_05630_),
    .A1(_05611_));
 sg13g2_a21oi_1 _06556_ (.A1(_05640_),
    .A2(_00429_),
    .Y(_00770_),
    .B1(_05650_));
 sg13g2_nor4_1 _06557_ (.A(_05652_),
    .B(_00556_),
    .C(_00768_),
    .D(_00770_),
    .Y(_00771_));
 sg13g2_nor2_1 _06558_ (.A(_05656_),
    .B(_00767_),
    .Y(_00772_));
 sg13g2_nand3_1 _06559_ (.B(_00771_),
    .C(_00772_),
    .A(_00769_),
    .Y(_00773_));
 sg13g2_nand2_1 _06560_ (.Y(_00774_),
    .A(net328),
    .B(net1207));
 sg13g2_nor2_1 _06561_ (.A(_05611_),
    .B(net1313),
    .Y(_00775_));
 sg13g2_a22oi_1 _06562_ (.Y(_00776_),
    .B1(net1269),
    .B2(\mac_inst.get_msu[0] ),
    .A2(net1316),
    .A1(\mac_inst.get_multiply[0] ));
 sg13g2_a22oi_1 _06563_ (.Y(_00777_),
    .B1(net1309),
    .B2(\cordic_atan2_result[0] ),
    .A2(net1273),
    .A1(\mac_inst.get_mac[0] ));
 sg13g2_nand2_1 _06564_ (.Y(_00778_),
    .A(_00776_),
    .B(_00777_));
 sg13g2_a21oi_1 _06565_ (.A1(\cordic_inst.cordic_state[56] ),
    .A2(net1228),
    .Y(_00779_),
    .B1(_00778_));
 sg13g2_o21ai_1 _06566_ (.B1(_00774_),
    .Y(_00153_),
    .A1(net1208),
    .A2(_00779_));
 sg13g2_nand2_1 _06567_ (.Y(_00780_),
    .A(net334),
    .B(net1207));
 sg13g2_a22oi_1 _06568_ (.Y(_00781_),
    .B1(net1310),
    .B2(\cordic_atan2_result[1] ),
    .A2(net1274),
    .A1(\mac_inst.get_mac[1] ));
 sg13g2_a22oi_1 _06569_ (.Y(_00782_),
    .B1(net1269),
    .B2(\mac_inst.get_msu[1] ),
    .A2(net1316),
    .A1(\mac_inst.get_multiply[1] ));
 sg13g2_nand2_1 _06570_ (.Y(_00783_),
    .A(_00781_),
    .B(_00782_));
 sg13g2_a21oi_1 _06571_ (.A1(\cordic_inst.cordic_state[57] ),
    .A2(net1229),
    .Y(_00784_),
    .B1(_00783_));
 sg13g2_o21ai_1 _06572_ (.B1(_00780_),
    .Y(_00154_),
    .A1(net1207),
    .A2(_00784_));
 sg13g2_nand2_1 _06573_ (.Y(_00785_),
    .A(net385),
    .B(net1205));
 sg13g2_a22oi_1 _06574_ (.Y(_00786_),
    .B1(net1269),
    .B2(\mac_inst.get_msu[2] ),
    .A2(net1316),
    .A1(net370));
 sg13g2_a22oi_1 _06575_ (.Y(_00787_),
    .B1(net1310),
    .B2(\cordic_atan2_result[2] ),
    .A2(net1274),
    .A1(\mac_inst.get_mac[2] ));
 sg13g2_nand2_1 _06576_ (.Y(_00788_),
    .A(_00786_),
    .B(_00787_));
 sg13g2_a21oi_1 _06577_ (.A1(\cordic_inst.cordic_state[58] ),
    .A2(net1229),
    .Y(_00789_),
    .B1(_00788_));
 sg13g2_o21ai_1 _06578_ (.B1(_00785_),
    .Y(_00155_),
    .A1(net1205),
    .A2(_00789_));
 sg13g2_nand2_1 _06579_ (.Y(_00790_),
    .A(net312),
    .B(net1203));
 sg13g2_a22oi_1 _06580_ (.Y(_00791_),
    .B1(net1274),
    .B2(\mac_inst.get_mac[3] ),
    .A2(net1314),
    .A1(\mac_inst.get_multiply[3] ));
 sg13g2_a22oi_1 _06581_ (.Y(_00792_),
    .B1(net1308),
    .B2(\cordic_atan2_result[3] ),
    .A2(net1268),
    .A1(\mac_inst.get_msu[3] ));
 sg13g2_nand2_1 _06582_ (.Y(_00793_),
    .A(_00791_),
    .B(_00792_));
 sg13g2_a21oi_1 _06583_ (.A1(\cordic_inst.cordic_state[59] ),
    .A2(net1227),
    .Y(_00794_),
    .B1(_00793_));
 sg13g2_o21ai_1 _06584_ (.B1(_00790_),
    .Y(_00156_),
    .A1(net1203),
    .A2(_00794_));
 sg13g2_nand2_1 _06585_ (.Y(_00795_),
    .A(net304),
    .B(net1205));
 sg13g2_a22oi_1 _06586_ (.Y(_00796_),
    .B1(net1268),
    .B2(\mac_inst.get_msu[4] ),
    .A2(net1315),
    .A1(\mac_inst.get_multiply[4] ));
 sg13g2_a22oi_1 _06587_ (.Y(_00797_),
    .B1(net1308),
    .B2(\cordic_atan2_result[4] ),
    .A2(net1272),
    .A1(\mac_inst.get_mac[4] ));
 sg13g2_nand2_1 _06588_ (.Y(_00798_),
    .A(_00796_),
    .B(_00797_));
 sg13g2_a21oi_1 _06589_ (.A1(\cordic_inst.cordic_state[60] ),
    .A2(net1230),
    .Y(_00799_),
    .B1(_00798_));
 sg13g2_o21ai_1 _06590_ (.B1(_00795_),
    .Y(_00157_),
    .A1(net1203),
    .A2(_00799_));
 sg13g2_nand2_1 _06591_ (.Y(_00800_),
    .A(net318),
    .B(net1209));
 sg13g2_a22oi_1 _06592_ (.Y(_00801_),
    .B1(net1267),
    .B2(\mac_inst.get_msu[5] ),
    .A2(net1314),
    .A1(\mac_inst.get_multiply[5] ));
 sg13g2_a22oi_1 _06593_ (.Y(_00802_),
    .B1(net1308),
    .B2(\cordic_atan2_result[5] ),
    .A2(net1272),
    .A1(\mac_inst.get_mac[5] ));
 sg13g2_nand2_1 _06594_ (.Y(_00803_),
    .A(_00801_),
    .B(_00802_));
 sg13g2_a21oi_1 _06595_ (.A1(\cordic_inst.cordic_state[61] ),
    .A2(net1229),
    .Y(_00804_),
    .B1(_00803_));
 sg13g2_o21ai_1 _06596_ (.B1(_00800_),
    .Y(_00158_),
    .A1(net1205),
    .A2(_00804_));
 sg13g2_nand2_1 _06597_ (.Y(_00805_),
    .A(net280),
    .B(net1203));
 sg13g2_a22oi_1 _06598_ (.Y(_00806_),
    .B1(net1268),
    .B2(\mac_inst.get_msu[6] ),
    .A2(net1314),
    .A1(\mac_inst.get_multiply[6] ));
 sg13g2_a22oi_1 _06599_ (.Y(_00807_),
    .B1(net1308),
    .B2(\cordic_atan2_result[6] ),
    .A2(net1272),
    .A1(\mac_inst.get_mac[6] ));
 sg13g2_nand2_1 _06600_ (.Y(_00808_),
    .A(_00806_),
    .B(_00807_));
 sg13g2_a21oi_1 _06601_ (.A1(\cordic_inst.cordic_state[62] ),
    .A2(net1230),
    .Y(_00809_),
    .B1(_00808_));
 sg13g2_o21ai_1 _06602_ (.B1(_00805_),
    .Y(_00159_),
    .A1(net1203),
    .A2(_00809_));
 sg13g2_nand2_1 _06603_ (.Y(_00810_),
    .A(net306),
    .B(net1209));
 sg13g2_a22oi_1 _06604_ (.Y(_00811_),
    .B1(net1267),
    .B2(\mac_inst.get_msu[7] ),
    .A2(net1314),
    .A1(\mac_inst.get_multiply[7] ));
 sg13g2_a22oi_1 _06605_ (.Y(_00812_),
    .B1(net1308),
    .B2(\cordic_atan2_result[7] ),
    .A2(net1272),
    .A1(\mac_inst.get_mac[7] ));
 sg13g2_nand2_1 _06606_ (.Y(_00813_),
    .A(_00811_),
    .B(_00812_));
 sg13g2_a21oi_1 _06607_ (.A1(\cordic_inst.cordic_state[63] ),
    .A2(net1229),
    .Y(_00814_),
    .B1(_00813_));
 sg13g2_o21ai_1 _06608_ (.B1(_00810_),
    .Y(_00160_),
    .A1(net1209),
    .A2(_00814_));
 sg13g2_nand2_1 _06609_ (.Y(_00815_),
    .A(net342),
    .B(net1203));
 sg13g2_a22oi_1 _06610_ (.Y(_00816_),
    .B1(net1272),
    .B2(\mac_inst.get_mac[8] ),
    .A2(net1314),
    .A1(\mac_inst.get_multiply[8] ));
 sg13g2_a22oi_1 _06611_ (.Y(_00817_),
    .B1(net1308),
    .B2(\cordic_atan2_result[8] ),
    .A2(net1267),
    .A1(\mac_inst.get_msu[8] ));
 sg13g2_nand2_2 _06612_ (.Y(_00818_),
    .A(_00816_),
    .B(_00817_));
 sg13g2_a21oi_2 _06613_ (.B1(_00818_),
    .Y(_00819_),
    .A2(net1227),
    .A1(\cordic_inst.cordic_state[64] ));
 sg13g2_o21ai_1 _06614_ (.B1(_00815_),
    .Y(_00161_),
    .A1(net1203),
    .A2(_00819_));
 sg13g2_nand2_1 _06615_ (.Y(_00820_),
    .A(net356),
    .B(net1204));
 sg13g2_a22oi_1 _06616_ (.Y(_00821_),
    .B1(net1272),
    .B2(\mac_inst.get_mac[9] ),
    .A2(net1314),
    .A1(\mac_inst.get_multiply[9] ));
 sg13g2_a22oi_1 _06617_ (.Y(_00822_),
    .B1(net1308),
    .B2(\cordic_atan2_result[9] ),
    .A2(net1267),
    .A1(\mac_inst.get_msu[9] ));
 sg13g2_nand2_2 _06618_ (.Y(_00823_),
    .A(_00821_),
    .B(_00822_));
 sg13g2_a21oi_2 _06619_ (.B1(_00823_),
    .Y(_00824_),
    .A2(net1227),
    .A1(\cordic_inst.cordic_state[65] ));
 sg13g2_o21ai_1 _06620_ (.B1(_00820_),
    .Y(_00162_),
    .A1(net1204),
    .A2(_00824_));
 sg13g2_nand2_1 _06621_ (.Y(_00825_),
    .A(net294),
    .B(net1205));
 sg13g2_a22oi_1 _06622_ (.Y(_00826_),
    .B1(net1267),
    .B2(\mac_inst.get_msu[10] ),
    .A2(net1314),
    .A1(\mac_inst.get_multiply[10] ));
 sg13g2_a22oi_1 _06623_ (.Y(_00827_),
    .B1(net1308),
    .B2(\cordic_atan2_result[10] ),
    .A2(net1272),
    .A1(\mac_inst.get_mac[10] ));
 sg13g2_nand2_1 _06624_ (.Y(_00828_),
    .A(_00826_),
    .B(_00827_));
 sg13g2_a21oi_2 _06625_ (.B1(_00828_),
    .Y(_00829_),
    .A2(net1227),
    .A1(\cordic_inst.cordic_state[66] ));
 sg13g2_o21ai_1 _06626_ (.B1(_00825_),
    .Y(_00163_),
    .A1(net1205),
    .A2(_00829_));
 sg13g2_nand2_1 _06627_ (.Y(_00830_),
    .A(net296),
    .B(net1204));
 sg13g2_a22oi_1 _06628_ (.Y(_00831_),
    .B1(net1267),
    .B2(\mac_inst.get_msu[11] ),
    .A2(net1314),
    .A1(\mac_inst.get_multiply[11] ));
 sg13g2_a22oi_1 _06629_ (.Y(_00832_),
    .B1(net1312),
    .B2(\cordic_atan2_result[11] ),
    .A2(net1272),
    .A1(\mac_inst.get_mac[11] ));
 sg13g2_nand2_1 _06630_ (.Y(_00833_),
    .A(_00831_),
    .B(_00832_));
 sg13g2_a21oi_2 _06631_ (.B1(_00833_),
    .Y(_00834_),
    .A2(net1227),
    .A1(\cordic_inst.cordic_state[67] ));
 sg13g2_o21ai_1 _06632_ (.B1(_00830_),
    .Y(_00164_),
    .A1(net1204),
    .A2(_00834_));
 sg13g2_nand2_1 _06633_ (.Y(_00835_),
    .A(\cordic_inst.cordic_state[68] ),
    .B(net1227));
 sg13g2_a22oi_1 _06634_ (.Y(_00836_),
    .B1(net1268),
    .B2(net433),
    .A2(net1315),
    .A1(\mac_inst.get_multiply[12] ));
 sg13g2_a22oi_1 _06635_ (.Y(_00837_),
    .B1(net1312),
    .B2(\cordic_atan2_result[12] ),
    .A2(net1276),
    .A1(net563));
 sg13g2_nand3_1 _06636_ (.B(_00836_),
    .C(_00837_),
    .A(_00835_),
    .Y(_00838_));
 sg13g2_mux2_1 _06637_ (.A0(_00838_),
    .A1(net576),
    .S(net1203),
    .X(_00165_));
 sg13g2_nand2_1 _06638_ (.Y(_00839_),
    .A(net286),
    .B(net1205));
 sg13g2_a22oi_1 _06639_ (.Y(_00840_),
    .B1(net1267),
    .B2(\mac_inst.get_msu[13] ),
    .A2(net1315),
    .A1(\mac_inst.get_multiply[13] ));
 sg13g2_a22oi_1 _06640_ (.Y(_00841_),
    .B1(net1310),
    .B2(\cordic_atan2_result[13] ),
    .A2(net1274),
    .A1(\mac_inst.get_mac[13] ));
 sg13g2_nand2_1 _06641_ (.Y(_00842_),
    .A(_00840_),
    .B(_00841_));
 sg13g2_a21oi_2 _06642_ (.B1(_00842_),
    .Y(_00843_),
    .A2(net1228),
    .A1(\cordic_inst.cordic_state[69] ));
 sg13g2_o21ai_1 _06643_ (.B1(_00839_),
    .Y(_00166_),
    .A1(net1206),
    .A2(_00843_));
 sg13g2_nand2_1 _06644_ (.Y(_00844_),
    .A(\cordic_inst.cordic_state[70] ),
    .B(net1227));
 sg13g2_a22oi_1 _06645_ (.Y(_00845_),
    .B1(net1311),
    .B2(\cordic_atan2_result[14] ),
    .A2(net1275),
    .A1(\mac_inst.get_mac[14] ));
 sg13g2_a22oi_1 _06646_ (.Y(_00846_),
    .B1(net1267),
    .B2(net534),
    .A2(net1315),
    .A1(net404));
 sg13g2_nand3_1 _06647_ (.B(_00845_),
    .C(_00846_),
    .A(_00844_),
    .Y(_00847_));
 sg13g2_mux2_1 _06648_ (.A0(_00847_),
    .A1(net566),
    .S(net1204),
    .X(_00167_));
 sg13g2_nand2_1 _06649_ (.Y(_00848_),
    .A(\cordic_inst.cordic_state[71] ),
    .B(net1228));
 sg13g2_a22oi_1 _06650_ (.Y(_00849_),
    .B1(net1311),
    .B2(\cordic_atan2_result[15] ),
    .A2(net1275),
    .A1(\mac_inst.get_mac[15] ));
 sg13g2_a22oi_1 _06651_ (.Y(_00850_),
    .B1(net1269),
    .B2(\mac_inst.get_msu[15] ),
    .A2(net1316),
    .A1(\mac_inst.get_multiply[15] ));
 sg13g2_nand3_1 _06652_ (.B(_00849_),
    .C(_00850_),
    .A(_00848_),
    .Y(_00851_));
 sg13g2_mux2_1 _06653_ (.A0(_00851_),
    .A1(net571),
    .S(net1206),
    .X(_00168_));
 sg13g2_nand2_1 _06654_ (.Y(_00852_),
    .A(\cordic_inst.cordic_state[72] ),
    .B(net1228));
 sg13g2_a22oi_1 _06655_ (.Y(_00853_),
    .B1(net1269),
    .B2(\mac_inst.get_msu[16] ),
    .A2(net1316),
    .A1(\mac_inst.get_multiply[16] ));
 sg13g2_a22oi_1 _06656_ (.Y(_00854_),
    .B1(net1311),
    .B2(\cordic_atan2_result[16] ),
    .A2(net1275),
    .A1(\mac_inst.get_mac[16] ));
 sg13g2_nand3_1 _06657_ (.B(_00853_),
    .C(_00854_),
    .A(_00852_),
    .Y(_00855_));
 sg13g2_mux2_1 _06658_ (.A0(_00855_),
    .A1(net605),
    .S(net1206),
    .X(_00169_));
 sg13g2_nand2_1 _06659_ (.Y(_00856_),
    .A(net387),
    .B(net1208));
 sg13g2_a22oi_1 _06660_ (.Y(_00857_),
    .B1(net1269),
    .B2(\mac_inst.get_msu[17] ),
    .A2(net1316),
    .A1(net362));
 sg13g2_a22oi_1 _06661_ (.Y(_00858_),
    .B1(net1309),
    .B2(\cordic_atan2_result[17] ),
    .A2(net1273),
    .A1(\mac_inst.get_mac[17] ));
 sg13g2_nand2_1 _06662_ (.Y(_00859_),
    .A(_00857_),
    .B(_00858_));
 sg13g2_a21oi_2 _06663_ (.B1(_00859_),
    .Y(_00860_),
    .A2(net1228),
    .A1(\cordic_inst.cordic_state[73] ));
 sg13g2_o21ai_1 _06664_ (.B1(_00856_),
    .Y(_00170_),
    .A1(net1208),
    .A2(_00860_));
 sg13g2_nand2_1 _06665_ (.Y(_00861_),
    .A(net298),
    .B(net1206));
 sg13g2_a22oi_1 _06666_ (.Y(_00862_),
    .B1(net1270),
    .B2(\mac_inst.get_msu[18] ),
    .A2(net1317),
    .A1(\mac_inst.get_multiply[18] ));
 sg13g2_a22oi_1 _06667_ (.Y(_00863_),
    .B1(net1309),
    .B2(\cordic_atan2_result[18] ),
    .A2(net1273),
    .A1(\mac_inst.get_mac[18] ));
 sg13g2_nand2_2 _06668_ (.Y(_00864_),
    .A(_00862_),
    .B(_00863_));
 sg13g2_a21oi_1 _06669_ (.A1(\cordic_inst.cordic_state[74] ),
    .A2(net1228),
    .Y(_00865_),
    .B1(_00864_));
 sg13g2_o21ai_1 _06670_ (.B1(_00861_),
    .Y(_00171_),
    .A1(net1205),
    .A2(_00865_));
 sg13g2_nand2_1 _06671_ (.Y(_00866_),
    .A(net338),
    .B(net1204));
 sg13g2_a22oi_1 _06672_ (.Y(_00867_),
    .B1(net1273),
    .B2(\mac_inst.get_mac[19] ),
    .A2(net1317),
    .A1(\mac_inst.get_multiply[19] ));
 sg13g2_a22oi_1 _06673_ (.Y(_00868_),
    .B1(net1309),
    .B2(\cordic_atan2_result[19] ),
    .A2(net1269),
    .A1(\mac_inst.get_msu[19] ));
 sg13g2_nand2_2 _06674_ (.Y(_00869_),
    .A(_00867_),
    .B(_00868_));
 sg13g2_a21oi_2 _06675_ (.B1(_00869_),
    .Y(_00870_),
    .A2(net1227),
    .A1(\cordic_inst.cordic_state[75] ));
 sg13g2_o21ai_1 _06676_ (.B1(_00866_),
    .Y(_00172_),
    .A1(net1204),
    .A2(_00870_));
 sg13g2_nand2_1 _06677_ (.Y(_00871_),
    .A(net314),
    .B(net1209));
 sg13g2_a22oi_1 _06678_ (.Y(_00872_),
    .B1(net1270),
    .B2(\mac_inst.get_msu[20] ),
    .A2(net1317),
    .A1(\mac_inst.get_multiply[20] ));
 sg13g2_a22oi_1 _06679_ (.Y(_00873_),
    .B1(net1309),
    .B2(\cordic_atan2_result[20] ),
    .A2(net1273),
    .A1(\mac_inst.get_mac[20] ));
 sg13g2_nand2_2 _06680_ (.Y(_00874_),
    .A(_00872_),
    .B(_00873_));
 sg13g2_a21oi_2 _06681_ (.B1(_00874_),
    .Y(_00875_),
    .A2(net1228),
    .A1(net1406));
 sg13g2_o21ai_1 _06682_ (.B1(_00871_),
    .Y(_00173_),
    .A1(net1209),
    .A2(_00875_));
 sg13g2_nand2_1 _06683_ (.Y(_00876_),
    .A(net310),
    .B(net1207));
 sg13g2_a22oi_1 _06684_ (.Y(_00877_),
    .B1(net1270),
    .B2(\mac_inst.get_msu[21] ),
    .A2(net1317),
    .A1(\mac_inst.get_multiply[21] ));
 sg13g2_a22oi_1 _06685_ (.Y(_00878_),
    .B1(net1309),
    .B2(\cordic_atan2_result[21] ),
    .A2(net1273),
    .A1(\mac_inst.get_mac[21] ));
 sg13g2_nand2_2 _06686_ (.Y(_00879_),
    .A(_00877_),
    .B(_00878_));
 sg13g2_a21oi_1 _06687_ (.A1(\cordic_inst.cordic_state[77] ),
    .A2(net1228),
    .Y(_00880_),
    .B1(_00879_));
 sg13g2_o21ai_1 _06688_ (.B1(_00876_),
    .Y(_00174_),
    .A1(net1207),
    .A2(_00880_));
 sg13g2_nand2_1 _06689_ (.Y(_00881_),
    .A(net336),
    .B(net1207));
 sg13g2_a22oi_1 _06690_ (.Y(_00882_),
    .B1(net1309),
    .B2(\cordic_atan2_result[22] ),
    .A2(net1273),
    .A1(\mac_inst.get_mac[22] ));
 sg13g2_a22oi_1 _06691_ (.Y(_00883_),
    .B1(net1269),
    .B2(\mac_inst.get_msu[22] ),
    .A2(net1316),
    .A1(\mac_inst.get_multiply[22] ));
 sg13g2_nand2_2 _06692_ (.Y(_00884_),
    .A(_00882_),
    .B(_00883_));
 sg13g2_a21oi_1 _06693_ (.A1(\cordic_inst.cordic_state[78] ),
    .A2(net1229),
    .Y(_00885_),
    .B1(_00884_));
 sg13g2_o21ai_1 _06694_ (.B1(_00881_),
    .Y(_00175_),
    .A1(net1209),
    .A2(_00885_));
 sg13g2_nand2_1 _06695_ (.Y(_00886_),
    .A(net352),
    .B(net1207));
 sg13g2_a22oi_1 _06696_ (.Y(_00887_),
    .B1(net1270),
    .B2(\mac_inst.get_msu[23] ),
    .A2(net1316),
    .A1(\mac_inst.get_multiply[23] ));
 sg13g2_a22oi_1 _06697_ (.Y(_00888_),
    .B1(net1309),
    .B2(\cordic_atan2_result[23] ),
    .A2(net1273),
    .A1(\mac_inst.get_mac[23] ));
 sg13g2_nand2_1 _06698_ (.Y(_00889_),
    .A(_00887_),
    .B(_00888_));
 sg13g2_a21oi_1 _06699_ (.A1(net1405),
    .A2(net1229),
    .Y(_00890_),
    .B1(_00889_));
 sg13g2_o21ai_1 _06700_ (.B1(_00886_),
    .Y(_00176_),
    .A1(net1207),
    .A2(_00890_));
 sg13g2_a21oi_1 _06701_ (.A1(net1561),
    .A2(\state[1] ),
    .Y(_00891_),
    .B1(_00444_));
 sg13g2_a221oi_1 _06702_ (.B2(_05600_),
    .C1(_00767_),
    .B1(_00768_),
    .A1(net1307),
    .Y(_00892_),
    .A2(_00427_));
 sg13g2_nand3b_1 _06703_ (.B(_00891_),
    .C(_00892_),
    .Y(_00893_),
    .A_N(_00457_));
 sg13g2_or2_1 _06704_ (.X(_00894_),
    .B(_00893_),
    .A(_00416_));
 sg13g2_and2_1 _06705_ (.A(net1326),
    .B(_00417_),
    .X(_00895_));
 sg13g2_a21o_1 _06706_ (.A2(_00895_),
    .A1(_00543_),
    .B1(net813),
    .X(_00896_));
 sg13g2_nor2_1 _06707_ (.A(_05618_),
    .B(_05623_),
    .Y(_00897_));
 sg13g2_a21oi_1 _06708_ (.A1(_05619_),
    .A2(_00896_),
    .Y(_00898_),
    .B1(_00897_));
 sg13g2_mux2_1 _06709_ (.A0(_00898_),
    .A1(net1465),
    .S(_00894_),
    .X(_00177_));
 sg13g2_a21oi_1 _06710_ (.A1(\state[2] ),
    .A2(_05618_),
    .Y(_00899_),
    .B1(_05623_));
 sg13g2_a221oi_1 _06711_ (.B2(_00895_),
    .C1(_00899_),
    .B1(_00543_),
    .A1(_05626_),
    .Y(_00900_),
    .A2(_00422_));
 sg13g2_mux2_1 _06712_ (.A0(_00900_),
    .A1(net774),
    .S(_00894_),
    .X(_00178_));
 sg13g2_xor2_1 _06713_ (.B(_00680_),
    .A(net668),
    .X(_00901_));
 sg13g2_nor2_1 _06714_ (.A(_00899_),
    .B(_00901_),
    .Y(_00902_));
 sg13g2_mux2_1 _06715_ (.A0(_00902_),
    .A1(net668),
    .S(_00894_),
    .X(_00179_));
 sg13g2_xnor2_1 _06716_ (.Y(_00903_),
    .A(_05595_),
    .B(_00684_));
 sg13g2_nor3_1 _06717_ (.A(_00894_),
    .B(_00899_),
    .C(_00903_),
    .Y(_00904_));
 sg13g2_a21o_1 _06718_ (.A2(_00894_),
    .A1(net772),
    .B1(_00904_),
    .X(_00180_));
 sg13g2_nand2b_1 _06719_ (.Y(_00905_),
    .B(net685),
    .A_N(net1480));
 sg13g2_nand3_1 _06720_ (.B(_00461_),
    .C(_00905_),
    .A(net1754),
    .Y(_00181_));
 sg13g2_nor2_1 _06721_ (.A(net1437),
    .B(net1442),
    .Y(_00906_));
 sg13g2_or2_1 _06722_ (.X(_00907_),
    .B(net1445),
    .A(net1440));
 sg13g2_nand4_1 _06723_ (.B(net1348),
    .C(_00487_),
    .A(net1427),
    .Y(_00908_),
    .D(net1346));
 sg13g2_a21oi_1 _06724_ (.A1(net737),
    .A2(_00908_),
    .Y(_00909_),
    .B1(net1323));
 sg13g2_nor2_1 _06725_ (.A(net1746),
    .B(_00909_),
    .Y(_00182_));
 sg13g2_a21oi_1 _06726_ (.A1(_05592_),
    .A2(_00908_),
    .Y(_00183_),
    .B1(_00466_));
 sg13g2_o21ai_1 _06727_ (.B1(net1285),
    .Y(_00910_),
    .A1(net1480),
    .A2(\cordic_inst.CASE_cordic_state_BITS_7_TO_3_0_3217_1_1901_2__ETC__q3[0] ));
 sg13g2_nand2_2 _06728_ (.Y(_00911_),
    .A(net672),
    .B(\cordic_inst.CASE_cordic_state_BITS_7_TO_3_0_3217_1_1901_2__ETC__q3[0] ));
 sg13g2_and2_1 _06729_ (.A(net1559),
    .B(net1481),
    .X(_00912_));
 sg13g2_a22oi_1 _06730_ (.Y(_00913_),
    .B1(_00912_),
    .B2(_00461_),
    .A2(_00911_),
    .A1(_00486_));
 sg13g2_a221oi_1 _06731_ (.B2(net1285),
    .C1(net1736),
    .B1(_00913_),
    .A1(_05587_),
    .Y(_00189_),
    .A2(_00910_));
 sg13g2_nand2b_1 _06732_ (.Y(_00914_),
    .B(\cordic_atan2_result[23] ),
    .A_N(\cordic_inst.IF_IF_cordic_state_BITS_2_TO_1_EQ_1_THEN_NOT_c_ETC___d36[1] ));
 sg13g2_nor4_1 _06733_ (.A(net1414),
    .B(\cordic_inst.cordic_state[49] ),
    .C(net1415),
    .D(\cordic_inst.cordic_state[47] ),
    .Y(_00915_));
 sg13g2_nor3_1 _06734_ (.A(net1411),
    .B(net1412),
    .C(net1413),
    .Y(_00916_));
 sg13g2_nor3_1 _06735_ (.A(\cordic_inst.cordic_state[34] ),
    .B(\cordic_inst.cordic_state[33] ),
    .C(\cordic_inst.cordic_state[32] ),
    .Y(_00917_));
 sg13g2_nor4_1 _06736_ (.A(net1425),
    .B(net1426),
    .C(\cordic_inst.cordic_state[36] ),
    .D(\cordic_inst.cordic_state[35] ),
    .Y(_00918_));
 sg13g2_nor4_1 _06737_ (.A(net1421),
    .B(net1422),
    .C(net1423),
    .D(net1424),
    .Y(_00919_));
 sg13g2_nor4_1 _06738_ (.A(net1417),
    .B(net1418),
    .C(net1419),
    .D(net1420),
    .Y(_00920_));
 sg13g2_nand4_1 _06739_ (.B(_00916_),
    .C(_00917_),
    .A(_00915_),
    .Y(_00921_),
    .D(_00918_));
 sg13g2_nand3_1 _06740_ (.B(_00919_),
    .C(_00920_),
    .A(_05582_),
    .Y(_00922_));
 sg13g2_nor2b_1 _06741_ (.A(net1409),
    .B_N(\cordic_inst.IF_IF_cordic_state_BITS_2_TO_1_EQ_1_THEN_NOT_c_ETC___d36[1] ),
    .Y(_00923_));
 sg13g2_o21ai_1 _06742_ (.B1(_00923_),
    .Y(_00924_),
    .A1(_00921_),
    .A2(_00922_));
 sg13g2_and2_1 _06743_ (.A(_00914_),
    .B(_00924_),
    .X(_00925_));
 sg13g2_nand2_1 _06744_ (.Y(_00926_),
    .A(_00914_),
    .B(_00924_));
 sg13g2_nand3_1 _06745_ (.B(_00914_),
    .C(_00924_),
    .A(\cordic_inst.CASE_cordic_state_BITS_7_TO_3_0_3217_1_1901_2__ETC__q3[0] ),
    .Y(_00927_));
 sg13g2_xor2_1 _06746_ (.B(_00927_),
    .A(\cordic_inst.CASE_cordic_state_BITS_7_TO_3_0_3217_1_1901_2__ETC__q3[1] ),
    .X(_00928_));
 sg13g2_nand2b_1 _06747_ (.Y(_00929_),
    .B(\cordic_atan2_result[1] ),
    .A_N(_00928_));
 sg13g2_nor2b_1 _06748_ (.A(\cordic_atan2_result[1] ),
    .B_N(_00928_),
    .Y(_00930_));
 sg13g2_xor2_1 _06749_ (.B(_00928_),
    .A(\cordic_atan2_result[1] ),
    .X(_00931_));
 sg13g2_xnor2_1 _06750_ (.Y(_00932_),
    .A(_00911_),
    .B(_00931_));
 sg13g2_and2_1 _06751_ (.A(_00461_),
    .B(net1285),
    .X(_00933_));
 sg13g2_nand2_1 _06752_ (.Y(_00934_),
    .A(_00461_),
    .B(net1285));
 sg13g2_a22oi_1 _06753_ (.Y(_00935_),
    .B1(_00482_),
    .B2(_00932_),
    .A2(net1482),
    .A1(_05574_));
 sg13g2_a22oi_1 _06754_ (.Y(_00936_),
    .B1(_00933_),
    .B2(_00935_),
    .A2(net1297),
    .A1(net776));
 sg13g2_nand2_1 _06755_ (.Y(_00190_),
    .A(net1761),
    .B(_00936_));
 sg13g2_o21ai_1 _06756_ (.B1(_00929_),
    .Y(_00937_),
    .A1(_00911_),
    .A2(_00930_));
 sg13g2_o21ai_1 _06757_ (.B1(net1243),
    .Y(_00938_),
    .A1(\cordic_inst.CASE_cordic_state_BITS_7_TO_3_0_3217_1_1901_2__ETC__q3[0] ),
    .A2(\cordic_inst.CASE_cordic_state_BITS_7_TO_3_0_3217_1_1901_2__ETC__q3[1] ));
 sg13g2_xor2_1 _06758_ (.B(_00938_),
    .A(\cordic_inst.CASE_cordic_state_BITS_7_TO_3_0_3217_1_1901_2__ETC__q3[2] ),
    .X(_00939_));
 sg13g2_nor2b_1 _06759_ (.A(_00939_),
    .B_N(\cordic_atan2_result[2] ),
    .Y(_00940_));
 sg13g2_xnor2_1 _06760_ (.Y(_00941_),
    .A(\cordic_atan2_result[2] ),
    .B(_00939_));
 sg13g2_o21ai_1 _06761_ (.B1(net1283),
    .Y(_00942_),
    .A1(_00937_),
    .A2(_00941_));
 sg13g2_a21oi_1 _06762_ (.A1(_00937_),
    .A2(_00941_),
    .Y(_00943_),
    .B1(_00942_));
 sg13g2_a21o_1 _06763_ (.A2(net1481),
    .A1(net1544),
    .B1(_00943_),
    .X(_00944_));
 sg13g2_a22oi_1 _06764_ (.Y(_00945_),
    .B1(net1235),
    .B2(_00944_),
    .A2(net1299),
    .A1(net695));
 sg13g2_nor2_1 _06765_ (.A(net1737),
    .B(net696),
    .Y(_00191_));
 sg13g2_a21oi_1 _06766_ (.A1(_00937_),
    .A2(_00941_),
    .Y(_00946_),
    .B1(_00940_));
 sg13g2_nor3_1 _06767_ (.A(\cordic_inst.CASE_cordic_state_BITS_7_TO_3_0_3217_1_1901_2__ETC__q3[0] ),
    .B(\cordic_inst.CASE_cordic_state_BITS_7_TO_3_0_3217_1_1901_2__ETC__q3[1] ),
    .C(\cordic_inst.CASE_cordic_state_BITS_7_TO_3_0_3217_1_1901_2__ETC__q3[2] ),
    .Y(_00947_));
 sg13g2_nor2_1 _06768_ (.A(net1237),
    .B(_00947_),
    .Y(_00948_));
 sg13g2_xor2_1 _06769_ (.B(_00948_),
    .A(\cordic_inst.CASE_cordic_state_BITS_7_TO_3_0_3217_1_1901_2__ETC__q3[3] ),
    .X(_00949_));
 sg13g2_nand2_1 _06770_ (.Y(_00950_),
    .A(\cordic_atan2_result[3] ),
    .B(_00949_));
 sg13g2_xnor2_1 _06771_ (.Y(_00951_),
    .A(\cordic_atan2_result[3] ),
    .B(_00949_));
 sg13g2_xnor2_1 _06772_ (.Y(_00952_),
    .A(_00946_),
    .B(_00951_));
 sg13g2_a221oi_1 _06773_ (.B2(_00952_),
    .C1(net1233),
    .B1(net1283),
    .A1(_05572_),
    .Y(_00953_),
    .A2(net1481));
 sg13g2_a21oi_1 _06774_ (.A1(net709),
    .A2(net1299),
    .Y(_00954_),
    .B1(_00953_));
 sg13g2_nand2_1 _06775_ (.Y(_00192_),
    .A(net1755),
    .B(net710));
 sg13g2_o21ai_1 _06776_ (.B1(_00950_),
    .Y(_00955_),
    .A1(_00946_),
    .A2(_00951_));
 sg13g2_nor2b_1 _06777_ (.A(\cordic_inst.CASE_cordic_state_BITS_7_TO_3_0_3217_1_1901_2__ETC__q3[3] ),
    .B_N(_00947_),
    .Y(_00956_));
 sg13g2_nor2_1 _06778_ (.A(net1237),
    .B(_00956_),
    .Y(_00957_));
 sg13g2_xnor2_1 _06779_ (.Y(_00958_),
    .A(\cordic_inst.CASE_cordic_state_BITS_7_TO_3_0_3217_1_1901_2__ETC__q3[4] ),
    .B(_00957_));
 sg13g2_nor2b_1 _06780_ (.A(_00958_),
    .B_N(\cordic_atan2_result[4] ),
    .Y(_00959_));
 sg13g2_xnor2_1 _06781_ (.Y(_00960_),
    .A(\cordic_atan2_result[4] ),
    .B(_00958_));
 sg13g2_o21ai_1 _06782_ (.B1(net1283),
    .Y(_00961_),
    .A1(_00955_),
    .A2(_00960_));
 sg13g2_a21oi_1 _06783_ (.A1(_00955_),
    .A2(_00960_),
    .Y(_00962_),
    .B1(_00961_));
 sg13g2_a21o_1 _06784_ (.A2(net1481),
    .A1(net1531),
    .B1(_00962_),
    .X(_00963_));
 sg13g2_a22oi_1 _06785_ (.Y(_00964_),
    .B1(net1235),
    .B2(_00963_),
    .A2(net1295),
    .A1(net657));
 sg13g2_nor2_1 _06786_ (.A(net1737),
    .B(_00964_),
    .Y(_00193_));
 sg13g2_a21oi_1 _06787_ (.A1(_00955_),
    .A2(_00960_),
    .Y(_00965_),
    .B1(_00959_));
 sg13g2_nor2b_1 _06788_ (.A(\cordic_inst.CASE_cordic_state_BITS_7_TO_3_0_3217_1_1901_2__ETC__q3[4] ),
    .B_N(_00956_),
    .Y(_00966_));
 sg13g2_nor2_1 _06789_ (.A(net1237),
    .B(_00966_),
    .Y(_00967_));
 sg13g2_xor2_1 _06790_ (.B(_00967_),
    .A(\cordic_inst.CASE_cordic_state_BITS_7_TO_3_0_3217_1_1901_2__ETC__q3[5] ),
    .X(_00968_));
 sg13g2_nand2_1 _06791_ (.Y(_00969_),
    .A(\cordic_atan2_result[5] ),
    .B(_00968_));
 sg13g2_xnor2_1 _06792_ (.Y(_00970_),
    .A(\cordic_atan2_result[5] ),
    .B(_00968_));
 sg13g2_xnor2_1 _06793_ (.Y(_00971_),
    .A(_00965_),
    .B(_00970_));
 sg13g2_a221oi_1 _06794_ (.B2(_00971_),
    .C1(net1233),
    .B1(net1284),
    .A1(_05571_),
    .Y(_00972_),
    .A2(net1481));
 sg13g2_a21oi_1 _06795_ (.A1(net682),
    .A2(net1296),
    .Y(_00973_),
    .B1(_00972_));
 sg13g2_nand2_1 _06796_ (.Y(_00194_),
    .A(net1755),
    .B(net683));
 sg13g2_o21ai_1 _06797_ (.B1(_00969_),
    .Y(_00974_),
    .A1(_00965_),
    .A2(_00970_));
 sg13g2_nor2b_1 _06798_ (.A(\cordic_inst.CASE_cordic_state_BITS_7_TO_3_0_3217_1_1901_2__ETC__q3[5] ),
    .B_N(_00966_),
    .Y(_00975_));
 sg13g2_nor2_1 _06799_ (.A(net1237),
    .B(_00975_),
    .Y(_00976_));
 sg13g2_xnor2_1 _06800_ (.Y(_00977_),
    .A(\cordic_inst.CASE_cordic_state_BITS_7_TO_3_0_3217_1_1901_2__ETC__q3[6] ),
    .B(_00976_));
 sg13g2_nor2b_1 _06801_ (.A(_00977_),
    .B_N(\cordic_atan2_result[6] ),
    .Y(_00978_));
 sg13g2_xnor2_1 _06802_ (.Y(_00979_),
    .A(\cordic_atan2_result[6] ),
    .B(_00977_));
 sg13g2_o21ai_1 _06803_ (.B1(net1283),
    .Y(_00980_),
    .A1(_00974_),
    .A2(_00979_));
 sg13g2_a21oi_1 _06804_ (.A1(_00974_),
    .A2(_00979_),
    .Y(_00981_),
    .B1(_00980_));
 sg13g2_a21o_1 _06805_ (.A2(net1480),
    .A1(net1525),
    .B1(_00981_),
    .X(_00982_));
 sg13g2_a22oi_1 _06806_ (.Y(_00983_),
    .B1(net1235),
    .B2(_00982_),
    .A2(net1296),
    .A1(net670));
 sg13g2_nor2_1 _06807_ (.A(net1736),
    .B(net671),
    .Y(_00195_));
 sg13g2_a21oi_1 _06808_ (.A1(_00974_),
    .A2(_00979_),
    .Y(_00984_),
    .B1(_00978_));
 sg13g2_nor2b_1 _06809_ (.A(\cordic_inst.CASE_cordic_state_BITS_7_TO_3_0_3217_1_1901_2__ETC__q3[6] ),
    .B_N(_00975_),
    .Y(_00985_));
 sg13g2_nor2_1 _06810_ (.A(net1237),
    .B(_00985_),
    .Y(_00986_));
 sg13g2_xor2_1 _06811_ (.B(_00986_),
    .A(\cordic_inst.CASE_cordic_state_BITS_7_TO_3_0_3217_1_1901_2__ETC__q3[7] ),
    .X(_00987_));
 sg13g2_nand2_1 _06812_ (.Y(_00988_),
    .A(\cordic_atan2_result[7] ),
    .B(_00987_));
 sg13g2_xnor2_1 _06813_ (.Y(_00989_),
    .A(\cordic_atan2_result[7] ),
    .B(_00987_));
 sg13g2_xnor2_1 _06814_ (.Y(_00990_),
    .A(_00984_),
    .B(_00989_));
 sg13g2_a221oi_1 _06815_ (.B2(_00990_),
    .C1(net1233),
    .B1(net1283),
    .A1(_05570_),
    .Y(_00991_),
    .A2(net1480));
 sg13g2_a21oi_1 _06816_ (.A1(net690),
    .A2(net1293),
    .Y(_00992_),
    .B1(_00991_));
 sg13g2_nand2_1 _06817_ (.Y(_00196_),
    .A(net1753),
    .B(_00992_));
 sg13g2_nand2_1 _06818_ (.Y(_00993_),
    .A(net1733),
    .B(net1480));
 sg13g2_o21ai_1 _06819_ (.B1(_00988_),
    .Y(_00994_),
    .A1(_00984_),
    .A2(_00989_));
 sg13g2_nand2b_1 _06820_ (.Y(_00995_),
    .B(_00985_),
    .A_N(\cordic_inst.CASE_cordic_state_BITS_7_TO_3_0_3217_1_1901_2__ETC__q3[7] ));
 sg13g2_nand2_1 _06821_ (.Y(_00996_),
    .A(net1243),
    .B(_00995_));
 sg13g2_xor2_1 _06822_ (.B(_00996_),
    .A(\cordic_inst.CASE_cordic_state_BITS_7_TO_3_0_3217_1_1901_2__ETC__q3[8] ),
    .X(_00997_));
 sg13g2_nor2b_1 _06823_ (.A(_00997_),
    .B_N(\cordic_atan2_result[8] ),
    .Y(_00998_));
 sg13g2_xnor2_1 _06824_ (.Y(_00999_),
    .A(\cordic_atan2_result[8] ),
    .B(_00997_));
 sg13g2_and2_1 _06825_ (.A(_00994_),
    .B(_00999_),
    .X(_01000_));
 sg13g2_o21ai_1 _06826_ (.B1(net1283),
    .Y(_01001_),
    .A1(_00994_),
    .A2(_00999_));
 sg13g2_o21ai_1 _06827_ (.B1(_00993_),
    .Y(_01002_),
    .A1(_01000_),
    .A2(_01001_));
 sg13g2_a22oi_1 _06828_ (.Y(_01003_),
    .B1(net1235),
    .B2(_01002_),
    .A2(net1293),
    .A1(net707));
 sg13g2_nor2_1 _06829_ (.A(net1736),
    .B(net708),
    .Y(_00197_));
 sg13g2_a21oi_1 _06830_ (.A1(_00994_),
    .A2(_00999_),
    .Y(_01004_),
    .B1(_00998_));
 sg13g2_o21ai_1 _06831_ (.B1(net1243),
    .Y(_01005_),
    .A1(\cordic_inst.CASE_cordic_state_BITS_7_TO_3_0_3217_1_1901_2__ETC__q3[8] ),
    .A2(_00995_));
 sg13g2_xor2_1 _06832_ (.B(_01005_),
    .A(\cordic_inst.CASE_cordic_state_BITS_7_TO_3_0_3217_1_1901_2__ETC__q3[9] ),
    .X(_01006_));
 sg13g2_inv_1 _06833_ (.Y(_01007_),
    .A(_01006_));
 sg13g2_nor2_1 _06834_ (.A(\cordic_atan2_result[9] ),
    .B(_01007_),
    .Y(_01008_));
 sg13g2_xnor2_1 _06835_ (.Y(_01009_),
    .A(\cordic_atan2_result[9] ),
    .B(_01006_));
 sg13g2_xor2_1 _06836_ (.B(_01009_),
    .A(_01004_),
    .X(_01010_));
 sg13g2_a221oi_1 _06837_ (.B2(_01010_),
    .C1(net1233),
    .B1(net1283),
    .A1(_05569_),
    .Y(_01011_),
    .A2(net1480));
 sg13g2_a21oi_1 _06838_ (.A1(net728),
    .A2(net1293),
    .Y(_01012_),
    .B1(_01011_));
 sg13g2_nand2_1 _06839_ (.Y(_00198_),
    .A(net1753),
    .B(_01012_));
 sg13g2_nand2_1 _06840_ (.Y(_01013_),
    .A(net584),
    .B(net1293));
 sg13g2_nand2_1 _06841_ (.Y(_01014_),
    .A(net1720),
    .B(net1480));
 sg13g2_nor3_1 _06842_ (.A(\cordic_inst.CASE_cordic_state_BITS_7_TO_3_0_3217_1_1901_2__ETC__q3[8] ),
    .B(\cordic_inst.CASE_cordic_state_BITS_7_TO_3_0_3217_1_1901_2__ETC__q3[9] ),
    .C(_00995_),
    .Y(_01015_));
 sg13g2_nor2_1 _06843_ (.A(net1237),
    .B(_01015_),
    .Y(_01016_));
 sg13g2_xnor2_1 _06844_ (.Y(_01017_),
    .A(\cordic_inst.CASE_cordic_state_BITS_7_TO_3_0_3217_1_1901_2__ETC__q3[10] ),
    .B(_01016_));
 sg13g2_xnor2_1 _06845_ (.Y(_01018_),
    .A(_05586_),
    .B(_01017_));
 sg13g2_a221oi_1 _06846_ (.B2(\cordic_atan2_result[9] ),
    .C1(_00998_),
    .B1(_01007_),
    .A1(_00994_),
    .Y(_01019_),
    .A2(_00999_));
 sg13g2_o21ai_1 _06847_ (.B1(_01018_),
    .Y(_01020_),
    .A1(_01008_),
    .A2(_01019_));
 sg13g2_or3_1 _06848_ (.A(_01008_),
    .B(_01018_),
    .C(_01019_),
    .X(_01021_));
 sg13g2_nand3_1 _06849_ (.B(_01020_),
    .C(_01021_),
    .A(net1283),
    .Y(_01022_));
 sg13g2_a21o_1 _06850_ (.A2(_01022_),
    .A1(_01014_),
    .B1(net1233),
    .X(_01023_));
 sg13g2_a21oi_1 _06851_ (.A1(_01013_),
    .A2(_01023_),
    .Y(_00199_),
    .B1(net1736));
 sg13g2_o21ai_1 _06852_ (.B1(_01021_),
    .Y(_01024_),
    .A1(_05586_),
    .A2(_01017_));
 sg13g2_nand2b_1 _06853_ (.Y(_01025_),
    .B(_01015_),
    .A_N(\cordic_inst.CASE_cordic_state_BITS_7_TO_3_0_3217_1_1901_2__ETC__q3[10] ));
 sg13g2_nand2_1 _06854_ (.Y(_01026_),
    .A(net1243),
    .B(_01025_));
 sg13g2_xor2_1 _06855_ (.B(_01026_),
    .A(\cordic_inst.CASE_cordic_state_BITS_7_TO_3_0_3217_1_1901_2__ETC__q3[11] ),
    .X(_01027_));
 sg13g2_nor2b_1 _06856_ (.A(_01027_),
    .B_N(\cordic_atan2_result[11] ),
    .Y(_01028_));
 sg13g2_nor2b_1 _06857_ (.A(\cordic_atan2_result[11] ),
    .B_N(_01027_),
    .Y(_01029_));
 sg13g2_inv_1 _06858_ (.Y(_01030_),
    .A(_01029_));
 sg13g2_nor2_1 _06859_ (.A(_01028_),
    .B(_01029_),
    .Y(_01031_));
 sg13g2_xnor2_1 _06860_ (.Y(_01032_),
    .A(_01024_),
    .B(_01031_));
 sg13g2_a221oi_1 _06861_ (.B2(_01032_),
    .C1(net1233),
    .B1(net1284),
    .A1(_05568_),
    .Y(_01033_),
    .A2(net1481));
 sg13g2_a21oi_1 _06862_ (.A1(net686),
    .A2(net1295),
    .Y(_01034_),
    .B1(_01033_));
 sg13g2_nand2_1 _06863_ (.Y(_00200_),
    .A(net1755),
    .B(net687));
 sg13g2_nand2_1 _06864_ (.Y(_01035_),
    .A(net1709),
    .B(net1483));
 sg13g2_nor2_2 _06865_ (.A(\cordic_inst.CASE_cordic_state_BITS_7_TO_3_0_3217_1_1901_2__ETC__q3[11] ),
    .B(_01025_),
    .Y(_01036_));
 sg13g2_nor2_2 _06866_ (.A(net1239),
    .B(_01036_),
    .Y(_01037_));
 sg13g2_xnor2_1 _06867_ (.Y(_01038_),
    .A(\cordic_atan2_result[12] ),
    .B(_01037_));
 sg13g2_a21oi_1 _06868_ (.A1(_01024_),
    .A2(_01030_),
    .Y(_01039_),
    .B1(_01028_));
 sg13g2_nor2_1 _06869_ (.A(_01038_),
    .B(_01039_),
    .Y(_01040_));
 sg13g2_a21o_1 _06870_ (.A2(_01039_),
    .A1(_01038_),
    .B1(_00483_),
    .X(_01041_));
 sg13g2_o21ai_1 _06871_ (.B1(_01035_),
    .Y(_01042_),
    .A1(_01040_),
    .A2(_01041_));
 sg13g2_a22oi_1 _06872_ (.Y(_01043_),
    .B1(net1235),
    .B2(_01042_),
    .A2(net1299),
    .A1(net697));
 sg13g2_nor2_1 _06873_ (.A(net1743),
    .B(net698),
    .Y(_00201_));
 sg13g2_a21oi_1 _06874_ (.A1(\cordic_atan2_result[12] ),
    .A2(_01037_),
    .Y(_01044_),
    .B1(_01040_));
 sg13g2_nor2_2 _06875_ (.A(\cordic_inst.CASE_cordic_state_BITS_7_TO_3_0_262144_1_13107_ETC__q2[19] ),
    .B(_01037_),
    .Y(_01045_));
 sg13g2_and2_1 _06876_ (.A(\cordic_inst.CASE_cordic_state_BITS_7_TO_3_0_262144_1_13107_ETC__q2[19] ),
    .B(net1246),
    .X(_01046_));
 sg13g2_nand2_1 _06877_ (.Y(_01047_),
    .A(\cordic_inst.CASE_cordic_state_BITS_7_TO_3_0_262144_1_13107_ETC__q2[19] ),
    .B(net1246));
 sg13g2_nor2_1 _06878_ (.A(_01036_),
    .B(_01047_),
    .Y(_01048_));
 sg13g2_nor2_1 _06879_ (.A(_01045_),
    .B(_01048_),
    .Y(_01049_));
 sg13g2_or2_1 _06880_ (.X(_01050_),
    .B(_01049_),
    .A(\cordic_atan2_result[13] ));
 sg13g2_inv_1 _06881_ (.Y(_01051_),
    .A(_01050_));
 sg13g2_nand2_1 _06882_ (.Y(_01052_),
    .A(\cordic_atan2_result[13] ),
    .B(_01049_));
 sg13g2_nand2_1 _06883_ (.Y(_01053_),
    .A(_01050_),
    .B(_01052_));
 sg13g2_xnor2_1 _06884_ (.Y(_01054_),
    .A(_01044_),
    .B(_01053_));
 sg13g2_a221oi_1 _06885_ (.B2(_01054_),
    .C1(net1233),
    .B1(net1284),
    .A1(_05566_),
    .Y(_01055_),
    .A2(net1483));
 sg13g2_a21oi_1 _06886_ (.A1(net674),
    .A2(net1299),
    .Y(_01056_),
    .B1(_01055_));
 sg13g2_nand2_1 _06887_ (.Y(_00202_),
    .A(net1761),
    .B(net675));
 sg13g2_nand2_1 _06888_ (.Y(_01057_),
    .A(net1698),
    .B(net1483));
 sg13g2_o21ai_1 _06889_ (.B1(_01047_),
    .Y(_01058_),
    .A1(net1239),
    .A2(_01036_));
 sg13g2_and2_1 _06890_ (.A(\cordic_atan2_result[14] ),
    .B(net1202),
    .X(_01059_));
 sg13g2_xor2_1 _06891_ (.B(net1202),
    .A(\cordic_atan2_result[14] ),
    .X(_01060_));
 sg13g2_a21oi_1 _06892_ (.A1(_01044_),
    .A2(_01052_),
    .Y(_01061_),
    .B1(_01051_));
 sg13g2_and2_1 _06893_ (.A(_01060_),
    .B(_01061_),
    .X(_01062_));
 sg13g2_o21ai_1 _06894_ (.B1(net1284),
    .Y(_01063_),
    .A1(_01060_),
    .A2(_01061_));
 sg13g2_o21ai_1 _06895_ (.B1(_01057_),
    .Y(_01064_),
    .A1(_01062_),
    .A2(_01063_));
 sg13g2_a22oi_1 _06896_ (.Y(_01065_),
    .B1(net1235),
    .B2(_01064_),
    .A2(net1299),
    .A1(net653));
 sg13g2_nor2_1 _06897_ (.A(net1744),
    .B(net654),
    .Y(_00203_));
 sg13g2_a21o_1 _06898_ (.A2(_01061_),
    .A1(_01060_),
    .B1(_01059_),
    .X(_01066_));
 sg13g2_nor2_2 _06899_ (.A(_01045_),
    .B(_01046_),
    .Y(_01067_));
 sg13g2_and2_1 _06900_ (.A(\cordic_atan2_result[15] ),
    .B(_01067_),
    .X(_01068_));
 sg13g2_nor2_1 _06901_ (.A(\cordic_atan2_result[15] ),
    .B(_01067_),
    .Y(_01069_));
 sg13g2_inv_1 _06902_ (.Y(_01070_),
    .A(_01069_));
 sg13g2_nor2_1 _06903_ (.A(_01068_),
    .B(_01069_),
    .Y(_01071_));
 sg13g2_xnor2_1 _06904_ (.Y(_01072_),
    .A(_01066_),
    .B(_01071_));
 sg13g2_a221oi_1 _06905_ (.B2(_01072_),
    .C1(net1233),
    .B1(net1284),
    .A1(_05565_),
    .Y(_01073_),
    .A2(net1482));
 sg13g2_a21oi_1 _06906_ (.A1(net703),
    .A2(net1297),
    .Y(_01074_),
    .B1(_01073_));
 sg13g2_nand2_1 _06907_ (.Y(_00204_),
    .A(net1761),
    .B(_01074_));
 sg13g2_nand2_1 _06908_ (.Y(_01075_),
    .A(net1684),
    .B(net1482));
 sg13g2_nand2_1 _06909_ (.Y(_01076_),
    .A(\cordic_atan2_result[16] ),
    .B(net1202));
 sg13g2_xor2_1 _06910_ (.B(net1202),
    .A(\cordic_atan2_result[16] ),
    .X(_01077_));
 sg13g2_inv_1 _06911_ (.Y(_01078_),
    .A(_01077_));
 sg13g2_a21oi_1 _06912_ (.A1(_01066_),
    .A2(_01070_),
    .Y(_01079_),
    .B1(_01068_));
 sg13g2_nor2_1 _06913_ (.A(_01078_),
    .B(_01079_),
    .Y(_01080_));
 sg13g2_a21o_1 _06914_ (.A2(_01079_),
    .A1(_01078_),
    .B1(_00483_),
    .X(_01081_));
 sg13g2_o21ai_1 _06915_ (.B1(_01075_),
    .Y(_01082_),
    .A1(_01080_),
    .A2(_01081_));
 sg13g2_a22oi_1 _06916_ (.Y(_01083_),
    .B1(net1235),
    .B2(_01082_),
    .A2(net1297),
    .A1(net681));
 sg13g2_nor2_1 _06917_ (.A(net1744),
    .B(_01083_),
    .Y(_00205_));
 sg13g2_o21ai_1 _06918_ (.B1(_01076_),
    .Y(_01084_),
    .A1(_01078_),
    .A2(_01079_));
 sg13g2_and2_1 _06919_ (.A(\cordic_atan2_result[17] ),
    .B(_01067_),
    .X(_01085_));
 sg13g2_nor2_1 _06920_ (.A(\cordic_atan2_result[17] ),
    .B(_01067_),
    .Y(_01086_));
 sg13g2_inv_1 _06921_ (.Y(_01087_),
    .A(_01086_));
 sg13g2_nor2_1 _06922_ (.A(_01085_),
    .B(_01086_),
    .Y(_01088_));
 sg13g2_xnor2_1 _06923_ (.Y(_01089_),
    .A(_01084_),
    .B(_01088_));
 sg13g2_a221oi_1 _06924_ (.B2(_01089_),
    .C1(net1234),
    .B1(net1284),
    .A1(_05563_),
    .Y(_01090_),
    .A2(net1482));
 sg13g2_a21oi_1 _06925_ (.A1(net676),
    .A2(net1297),
    .Y(_01091_),
    .B1(_01090_));
 sg13g2_nand2_1 _06926_ (.Y(_00206_),
    .A(net1761),
    .B(_01091_));
 sg13g2_nand2_1 _06927_ (.Y(_01092_),
    .A(net1674),
    .B(net1482));
 sg13g2_nand2_1 _06928_ (.Y(_01093_),
    .A(\cordic_atan2_result[18] ),
    .B(net1202));
 sg13g2_xor2_1 _06929_ (.B(net1202),
    .A(\cordic_atan2_result[18] ),
    .X(_01094_));
 sg13g2_inv_1 _06930_ (.Y(_01095_),
    .A(_01094_));
 sg13g2_a21oi_1 _06931_ (.A1(_01084_),
    .A2(_01087_),
    .Y(_01096_),
    .B1(_01085_));
 sg13g2_a21oi_1 _06932_ (.A1(_01095_),
    .A2(_01096_),
    .Y(_01097_),
    .B1(_00483_));
 sg13g2_o21ai_1 _06933_ (.B1(_01097_),
    .Y(_01098_),
    .A1(_01095_),
    .A2(_01096_));
 sg13g2_a21oi_1 _06934_ (.A1(_01092_),
    .A2(_01098_),
    .Y(_01099_),
    .B1(net1234));
 sg13g2_a21oi_1 _06935_ (.A1(net646),
    .A2(net1297),
    .Y(_01100_),
    .B1(_01099_));
 sg13g2_nor2_1 _06936_ (.A(net1743),
    .B(_01100_),
    .Y(_00207_));
 sg13g2_o21ai_1 _06937_ (.B1(_01093_),
    .Y(_01101_),
    .A1(_01095_),
    .A2(_01096_));
 sg13g2_nor3_1 _06938_ (.A(_05585_),
    .B(_01045_),
    .C(_01046_),
    .Y(_01102_));
 sg13g2_o21ai_1 _06939_ (.B1(_05585_),
    .Y(_01103_),
    .A1(_01045_),
    .A2(_01046_));
 sg13g2_nor2b_1 _06940_ (.A(_01102_),
    .B_N(_01103_),
    .Y(_01104_));
 sg13g2_xnor2_1 _06941_ (.Y(_01105_),
    .A(_01101_),
    .B(_01104_));
 sg13g2_a221oi_1 _06942_ (.B2(_01105_),
    .C1(net1234),
    .B1(net1284),
    .A1(_05562_),
    .Y(_01106_),
    .A2(net1482));
 sg13g2_a21oi_1 _06943_ (.A1(net711),
    .A2(net1297),
    .Y(_01107_),
    .B1(_01106_));
 sg13g2_nand2_1 _06944_ (.Y(_00208_),
    .A(net1758),
    .B(_01107_));
 sg13g2_nand2_1 _06945_ (.Y(_01108_),
    .A(net1666),
    .B(net1483));
 sg13g2_nand2_1 _06946_ (.Y(_01109_),
    .A(\cordic_atan2_result[20] ),
    .B(_01058_));
 sg13g2_xor2_1 _06947_ (.B(_01058_),
    .A(\cordic_atan2_result[20] ),
    .X(_01110_));
 sg13g2_inv_1 _06948_ (.Y(_01111_),
    .A(_01110_));
 sg13g2_a21oi_1 _06949_ (.A1(_01101_),
    .A2(_01103_),
    .Y(_01112_),
    .B1(_01102_));
 sg13g2_a21oi_1 _06950_ (.A1(_01111_),
    .A2(_01112_),
    .Y(_01113_),
    .B1(_00483_));
 sg13g2_o21ai_1 _06951_ (.B1(_01113_),
    .Y(_01114_),
    .A1(_01111_),
    .A2(_01112_));
 sg13g2_nand2_1 _06952_ (.Y(_01115_),
    .A(_01108_),
    .B(_01114_));
 sg13g2_a22oi_1 _06953_ (.Y(_01116_),
    .B1(_00933_),
    .B2(_01115_),
    .A2(net1298),
    .A1(net731));
 sg13g2_nor2_1 _06954_ (.A(net1744),
    .B(_01116_),
    .Y(_00209_));
 sg13g2_o21ai_1 _06955_ (.B1(_01109_),
    .Y(_01117_),
    .A1(_01111_),
    .A2(_01112_));
 sg13g2_and2_1 _06956_ (.A(\cordic_atan2_result[21] ),
    .B(_01067_),
    .X(_01118_));
 sg13g2_or2_1 _06957_ (.X(_01119_),
    .B(_01067_),
    .A(\cordic_atan2_result[21] ));
 sg13g2_nor2b_1 _06958_ (.A(_01118_),
    .B_N(_01119_),
    .Y(_01120_));
 sg13g2_xnor2_1 _06959_ (.Y(_01121_),
    .A(_01117_),
    .B(_01120_));
 sg13g2_a221oi_1 _06960_ (.B2(_01121_),
    .C1(net1234),
    .B1(_00482_),
    .A1(_05561_),
    .Y(_01122_),
    .A2(net1482));
 sg13g2_a21oi_1 _06961_ (.A1(net766),
    .A2(net1298),
    .Y(_01123_),
    .B1(_01122_));
 sg13g2_nand2_1 _06962_ (.Y(_00210_),
    .A(net1762),
    .B(_01123_));
 sg13g2_nand2_1 _06963_ (.Y(_01124_),
    .A(net1658),
    .B(net1484));
 sg13g2_xnor2_1 _06964_ (.Y(_01125_),
    .A(\cordic_atan2_result[22] ),
    .B(net1202));
 sg13g2_a21oi_1 _06965_ (.A1(_01117_),
    .A2(_01119_),
    .Y(_01126_),
    .B1(_01118_));
 sg13g2_nor2_1 _06966_ (.A(_01125_),
    .B(_01126_),
    .Y(_01127_));
 sg13g2_a21o_1 _06967_ (.A2(_01126_),
    .A1(_01125_),
    .B1(_00483_),
    .X(_01128_));
 sg13g2_o21ai_1 _06968_ (.B1(_01124_),
    .Y(_01129_),
    .A1(_01127_),
    .A2(_01128_));
 sg13g2_a22oi_1 _06969_ (.Y(_01130_),
    .B1(net1235),
    .B2(_01129_),
    .A2(net1297),
    .A1(net679));
 sg13g2_nor2_1 _06970_ (.A(net1744),
    .B(_01130_),
    .Y(_00211_));
 sg13g2_a21oi_1 _06971_ (.A1(net679),
    .A2(net1202),
    .Y(_01131_),
    .B1(_01127_));
 sg13g2_xnor2_1 _06972_ (.Y(_01132_),
    .A(\cordic_atan2_result[23] ),
    .B(_01067_));
 sg13g2_xnor2_1 _06973_ (.Y(_01133_),
    .A(_01131_),
    .B(_01132_));
 sg13g2_a221oi_1 _06974_ (.B2(_01133_),
    .C1(net1234),
    .B1(_00482_),
    .A1(_05560_),
    .Y(_01134_),
    .A2(net1482));
 sg13g2_a21oi_1 _06975_ (.A1(net738),
    .A2(net1297),
    .Y(_01135_),
    .B1(net1744));
 sg13g2_nand2b_1 _06976_ (.Y(_00212_),
    .B(_01135_),
    .A_N(_01134_));
 sg13g2_mux4_1 _06977_ (.S0(net1460),
    .A0(\cordic_inst.cordic_state[64] ),
    .A1(\cordic_inst.cordic_state[65] ),
    .A2(\cordic_inst.cordic_state[66] ),
    .A3(\cordic_inst.cordic_state[67] ),
    .S1(net1451),
    .X(_01136_));
 sg13g2_mux4_1 _06978_ (.S0(net1459),
    .A0(\cordic_inst.cordic_state[68] ),
    .A1(\cordic_inst.cordic_state[69] ),
    .A2(\cordic_inst.cordic_state[70] ),
    .A3(\cordic_inst.cordic_state[71] ),
    .S1(net1451),
    .X(_01137_));
 sg13g2_mux2_1 _06979_ (.A0(_01136_),
    .A1(_01137_),
    .S(net1444),
    .X(_01138_));
 sg13g2_nand2_1 _06980_ (.Y(_01139_),
    .A(net1439),
    .B(_01138_));
 sg13g2_mux4_1 _06981_ (.S0(net1461),
    .A0(\cordic_inst.cordic_state[56] ),
    .A1(\cordic_inst.cordic_state[57] ),
    .A2(\cordic_inst.cordic_state[58] ),
    .A3(\cordic_inst.cordic_state[59] ),
    .S1(net1453),
    .X(_01140_));
 sg13g2_nor2b_2 _06982_ (.A(net1440),
    .B_N(net1444),
    .Y(_01141_));
 sg13g2_nand2b_2 _06983_ (.Y(_01142_),
    .B(net1444),
    .A_N(\cordic_inst.cordic_state[6] ));
 sg13g2_mux4_1 _06984_ (.S0(net1461),
    .A0(\cordic_inst.cordic_state[60] ),
    .A1(\cordic_inst.cordic_state[61] ),
    .A2(\cordic_inst.cordic_state[62] ),
    .A3(\cordic_inst.cordic_state[63] ),
    .S1(net1452),
    .X(_01143_));
 sg13g2_a22oi_1 _06985_ (.Y(_01144_),
    .B1(_01141_),
    .B2(_01143_),
    .A2(_01140_),
    .A1(net1346));
 sg13g2_a21oi_2 _06986_ (.B1(net1431),
    .Y(_01145_),
    .A2(_01144_),
    .A1(_01139_));
 sg13g2_nor2_2 _06987_ (.A(_05576_),
    .B(net1394),
    .Y(_01146_));
 sg13g2_nand2_1 _06988_ (.Y(_01147_),
    .A(_00499_),
    .B(_01146_));
 sg13g2_mux4_1 _06989_ (.S0(net1460),
    .A0(\cordic_inst.cordic_state[72] ),
    .A1(\cordic_inst.cordic_state[73] ),
    .A2(\cordic_inst.cordic_state[74] ),
    .A3(\cordic_inst.cordic_state[75] ),
    .S1(net1451),
    .X(_01148_));
 sg13g2_mux2_1 _06990_ (.A0(\cordic_inst.cordic_state[78] ),
    .A1(net1404),
    .S(net1457),
    .X(_01149_));
 sg13g2_mux4_1 _06991_ (.S0(net1459),
    .A0(net1406),
    .A1(\cordic_inst.cordic_state[77] ),
    .A2(\cordic_inst.cordic_state[78] ),
    .A3(net1404),
    .S1(net1451),
    .X(_01150_));
 sg13g2_mux2_1 _06992_ (.A0(_01148_),
    .A1(_01150_),
    .S(net1444),
    .X(_01151_));
 sg13g2_inv_1 _06993_ (.Y(_01152_),
    .A(_01151_));
 sg13g2_nand2_1 _06994_ (.Y(_01153_),
    .A(net1392),
    .B(_01151_));
 sg13g2_o21ai_1 _06995_ (.B1(_01147_),
    .Y(_01154_),
    .A1(net1395),
    .A2(_01153_));
 sg13g2_nor2_2 _06996_ (.A(_01145_),
    .B(_01154_),
    .Y(_01155_));
 sg13g2_nor2_1 _06997_ (.A(\cordic_inst.cordic_state[32] ),
    .B(_01155_),
    .Y(_01156_));
 sg13g2_or2_1 _06998_ (.X(_01157_),
    .B(_01155_),
    .A(\cordic_inst.cordic_state[32] ));
 sg13g2_xnor2_1 _06999_ (.Y(_01158_),
    .A(\cordic_inst.cordic_state[32] ),
    .B(_01155_));
 sg13g2_a22oi_1 _07000_ (.Y(_01159_),
    .B1(net1280),
    .B2(_01158_),
    .A2(net1476),
    .A1(net1559));
 sg13g2_nand2_1 _07001_ (.Y(_01160_),
    .A(net1371),
    .B(_01159_));
 sg13g2_o21ai_1 _07002_ (.B1(_01160_),
    .Y(_01161_),
    .A1(net1654),
    .A2(net1371));
 sg13g2_o21ai_1 _07003_ (.B1(net1766),
    .Y(_01162_),
    .A1(net786),
    .A2(net1289));
 sg13g2_a21oi_1 _07004_ (.A1(net1289),
    .A2(_01161_),
    .Y(_00213_),
    .B1(_01162_));
 sg13g2_mux2_1 _07005_ (.A0(\cordic_inst.cordic_state[73] ),
    .A1(\cordic_inst.cordic_state[74] ),
    .S(net1460),
    .X(_01163_));
 sg13g2_nand2_1 _07006_ (.Y(_01164_),
    .A(net1406),
    .B(net1460));
 sg13g2_o21ai_1 _07007_ (.B1(_01164_),
    .Y(_01165_),
    .A1(_05578_),
    .A2(net1460));
 sg13g2_mux4_1 _07008_ (.S0(net1459),
    .A0(\cordic_inst.cordic_state[73] ),
    .A1(\cordic_inst.cordic_state[74] ),
    .A2(\cordic_inst.cordic_state[75] ),
    .A3(net1406),
    .S1(net1451),
    .X(_01166_));
 sg13g2_nor2_1 _07009_ (.A(net1444),
    .B(_01166_),
    .Y(_01167_));
 sg13g2_mux2_1 _07010_ (.A0(\cordic_inst.cordic_state[77] ),
    .A1(\cordic_inst.cordic_state[78] ),
    .S(net1458),
    .X(_01168_));
 sg13g2_nor2b_2 _07011_ (.A(net1457),
    .B_N(net1446),
    .Y(_01169_));
 sg13g2_a22oi_1 _07012_ (.Y(_01170_),
    .B1(_01169_),
    .B2(net1404),
    .A2(_01168_),
    .A1(net1385));
 sg13g2_a221oi_1 _07013_ (.B2(net1404),
    .C1(net1388),
    .B1(_01169_),
    .A1(net1385),
    .Y(_01171_),
    .A2(_01168_));
 sg13g2_or2_1 _07014_ (.X(_01172_),
    .B(_01171_),
    .A(_01167_));
 sg13g2_nand2b_1 _07015_ (.Y(_01173_),
    .B(net1391),
    .A_N(_01172_));
 sg13g2_or4_1 _07016_ (.A(net1396),
    .B(net1441),
    .C(_01167_),
    .D(_01171_),
    .X(_01174_));
 sg13g2_mux2_1 _07017_ (.A0(\cordic_inst.cordic_state[69] ),
    .A1(\cordic_inst.cordic_state[70] ),
    .S(net1458),
    .X(_01175_));
 sg13g2_mux2_1 _07018_ (.A0(\cordic_inst.cordic_state[71] ),
    .A1(\cordic_inst.cordic_state[72] ),
    .S(net1459),
    .X(_01176_));
 sg13g2_mux2_1 _07019_ (.A0(_01175_),
    .A1(_01176_),
    .S(net1450),
    .X(_01177_));
 sg13g2_mux2_1 _07020_ (.A0(\cordic_inst.cordic_state[65] ),
    .A1(\cordic_inst.cordic_state[66] ),
    .S(net1458),
    .X(_01178_));
 sg13g2_mux2_1 _07021_ (.A0(\cordic_inst.cordic_state[67] ),
    .A1(\cordic_inst.cordic_state[68] ),
    .S(net1458),
    .X(_01179_));
 sg13g2_mux2_1 _07022_ (.A0(_01178_),
    .A1(_01179_),
    .S(net1446),
    .X(_01180_));
 sg13g2_mux4_1 _07023_ (.S0(net1450),
    .A0(_01175_),
    .A1(_01176_),
    .A2(_01178_),
    .A3(_01179_),
    .S1(net1389),
    .X(_01181_));
 sg13g2_nor2_1 _07024_ (.A(net1392),
    .B(_01181_),
    .Y(_01182_));
 sg13g2_mux2_1 _07025_ (.A0(\cordic_inst.cordic_state[59] ),
    .A1(\cordic_inst.cordic_state[60] ),
    .S(net1461),
    .X(_01183_));
 sg13g2_mux2_1 _07026_ (.A0(\cordic_inst.cordic_state[57] ),
    .A1(\cordic_inst.cordic_state[58] ),
    .S(net1461),
    .X(_01184_));
 sg13g2_mux2_1 _07027_ (.A0(\cordic_inst.cordic_state[63] ),
    .A1(\cordic_inst.cordic_state[64] ),
    .S(net1459),
    .X(_01185_));
 sg13g2_mux2_1 _07028_ (.A0(\cordic_inst.cordic_state[61] ),
    .A1(\cordic_inst.cordic_state[62] ),
    .S(net1461),
    .X(_01186_));
 sg13g2_mux2_1 _07029_ (.A0(_01185_),
    .A1(_01186_),
    .S(net1387),
    .X(_01187_));
 sg13g2_mux4_1 _07030_ (.S0(net1387),
    .A0(_01183_),
    .A1(_01184_),
    .A2(_01185_),
    .A3(_01186_),
    .S1(net1444),
    .X(_01188_));
 sg13g2_o21ai_1 _07031_ (.B1(net1395),
    .Y(_01189_),
    .A1(net1439),
    .A2(_01188_));
 sg13g2_o21ai_1 _07032_ (.B1(_01174_),
    .Y(_01190_),
    .A1(_01182_),
    .A2(_01189_));
 sg13g2_nor2b_1 _07033_ (.A(_01190_),
    .B_N(_01147_),
    .Y(_01191_));
 sg13g2_o21ai_1 _07034_ (.B1(net1244),
    .Y(_01192_),
    .A1(_01145_),
    .A2(_01154_));
 sg13g2_xnor2_1 _07035_ (.Y(_01193_),
    .A(_01191_),
    .B(_01192_));
 sg13g2_nand2_1 _07036_ (.Y(_01194_),
    .A(\cordic_inst.cordic_state[33] ),
    .B(_01193_));
 sg13g2_inv_1 _07037_ (.Y(_01195_),
    .A(_01194_));
 sg13g2_nor2_1 _07038_ (.A(\cordic_inst.cordic_state[33] ),
    .B(_01193_),
    .Y(_01196_));
 sg13g2_nor2_1 _07039_ (.A(_01195_),
    .B(_01196_),
    .Y(_01197_));
 sg13g2_a21oi_1 _07040_ (.A1(_01157_),
    .A2(_01197_),
    .Y(_01198_),
    .B1(net1324));
 sg13g2_o21ai_1 _07041_ (.B1(_01198_),
    .Y(_01199_),
    .A1(_01157_),
    .A2(_01197_));
 sg13g2_a22oi_1 _07042_ (.Y(_01200_),
    .B1(net1321),
    .B2(net1554),
    .A2(net1366),
    .A1(net1635));
 sg13g2_a21oi_1 _07043_ (.A1(_01199_),
    .A2(_01200_),
    .Y(_01201_),
    .B1(net1302));
 sg13g2_a21oi_1 _07044_ (.A1(net767),
    .A2(net1302),
    .Y(_01202_),
    .B1(_01201_));
 sg13g2_nand2_1 _07045_ (.Y(_00214_),
    .A(net1778),
    .B(_01202_));
 sg13g2_mux4_1 _07046_ (.S0(net1459),
    .A0(\cordic_inst.cordic_state[70] ),
    .A1(\cordic_inst.cordic_state[71] ),
    .A2(\cordic_inst.cordic_state[72] ),
    .A3(\cordic_inst.cordic_state[73] ),
    .S1(net1451),
    .X(_01203_));
 sg13g2_mux4_1 _07047_ (.S0(net1458),
    .A0(\cordic_inst.cordic_state[66] ),
    .A1(\cordic_inst.cordic_state[67] ),
    .A2(\cordic_inst.cordic_state[68] ),
    .A3(\cordic_inst.cordic_state[69] ),
    .S1(net1451),
    .X(_01204_));
 sg13g2_mux2_1 _07048_ (.A0(_01203_),
    .A1(_01204_),
    .S(net1389),
    .X(_01205_));
 sg13g2_mux4_1 _07049_ (.S0(net1461),
    .A0(\cordic_inst.cordic_state[58] ),
    .A1(\cordic_inst.cordic_state[59] ),
    .A2(\cordic_inst.cordic_state[60] ),
    .A3(\cordic_inst.cordic_state[61] ),
    .S1(net1453),
    .X(_01206_));
 sg13g2_and2_1 _07050_ (.A(net1346),
    .B(_01206_),
    .X(_01207_));
 sg13g2_mux4_1 _07051_ (.S0(net1459),
    .A0(\cordic_inst.cordic_state[62] ),
    .A1(\cordic_inst.cordic_state[63] ),
    .A2(\cordic_inst.cordic_state[64] ),
    .A3(\cordic_inst.cordic_state[65] ),
    .S1(net1452),
    .X(_01208_));
 sg13g2_a221oi_1 _07052_ (.B2(_01141_),
    .C1(_01207_),
    .B1(_01208_),
    .A1(net1439),
    .Y(_01209_),
    .A2(_01205_));
 sg13g2_nand2_1 _07053_ (.Y(_01210_),
    .A(net1385),
    .B(_01149_));
 sg13g2_mux4_1 _07054_ (.S0(net1459),
    .A0(\cordic_inst.cordic_state[74] ),
    .A1(\cordic_inst.cordic_state[75] ),
    .A2(net1406),
    .A3(\cordic_inst.cordic_state[77] ),
    .S1(net1451),
    .X(_01211_));
 sg13g2_nand2_1 _07055_ (.Y(_01212_),
    .A(net1389),
    .B(_01211_));
 sg13g2_o21ai_1 _07056_ (.B1(_01212_),
    .Y(_01213_),
    .A1(net1389),
    .A2(_01210_));
 sg13g2_and2_1 _07057_ (.A(net1392),
    .B(_01213_),
    .X(_01214_));
 sg13g2_o21ai_1 _07058_ (.B1(net1392),
    .Y(_01215_),
    .A1(net1389),
    .A2(_00506_));
 sg13g2_nand2_1 _07059_ (.Y(_01216_),
    .A(_01146_),
    .B(_01215_));
 sg13g2_o21ai_1 _07060_ (.B1(_01216_),
    .Y(_01217_),
    .A1(net1431),
    .A2(_01209_));
 sg13g2_a21o_1 _07061_ (.A2(_01214_),
    .A1(net1431),
    .B1(_01217_),
    .X(_01218_));
 sg13g2_nor3_1 _07062_ (.A(_01145_),
    .B(_01154_),
    .C(_01190_),
    .Y(_01219_));
 sg13g2_nor2_1 _07063_ (.A(net1238),
    .B(_01219_),
    .Y(_01220_));
 sg13g2_xnor2_1 _07064_ (.Y(_01221_),
    .A(_01218_),
    .B(_01220_));
 sg13g2_and2_1 _07065_ (.A(\cordic_inst.cordic_state[34] ),
    .B(_01221_),
    .X(_01222_));
 sg13g2_xor2_1 _07066_ (.B(_01221_),
    .A(\cordic_inst.cordic_state[34] ),
    .X(_01223_));
 sg13g2_o21ai_1 _07067_ (.B1(_01194_),
    .Y(_01224_),
    .A1(_01156_),
    .A2(_01196_));
 sg13g2_and2_1 _07068_ (.A(_01223_),
    .B(_01224_),
    .X(_01225_));
 sg13g2_o21ai_1 _07069_ (.B1(net1280),
    .Y(_01226_),
    .A1(_01223_),
    .A2(_01224_));
 sg13g2_a21oi_1 _07070_ (.A1(net1548),
    .A2(net1476),
    .Y(_01227_),
    .B1(net1368));
 sg13g2_o21ai_1 _07071_ (.B1(_01227_),
    .Y(_01228_),
    .A1(_01225_),
    .A2(_01226_));
 sg13g2_o21ai_1 _07072_ (.B1(_01228_),
    .Y(_01229_),
    .A1(net1629),
    .A2(net1371));
 sg13g2_nand2_1 _07073_ (.Y(_01230_),
    .A(net699),
    .B(net1302));
 sg13g2_a21oi_1 _07074_ (.A1(_01229_),
    .A2(_01230_),
    .Y(_00215_),
    .B1(net1748));
 sg13g2_a21oi_1 _07075_ (.A1(_01223_),
    .A2(_01224_),
    .Y(_01231_),
    .B1(_01222_));
 sg13g2_mux2_1 _07076_ (.A0(_01163_),
    .A1(_01176_),
    .S(net1385),
    .X(_01232_));
 sg13g2_mux2_1 _07077_ (.A0(_01175_),
    .A1(_01179_),
    .S(net1385),
    .X(_01233_));
 sg13g2_mux2_1 _07078_ (.A0(_01232_),
    .A1(_01233_),
    .S(_05590_),
    .X(_01234_));
 sg13g2_nor2_1 _07079_ (.A(net1393),
    .B(_01234_),
    .Y(_01235_));
 sg13g2_nand2_1 _07080_ (.Y(_01236_),
    .A(net1452),
    .B(_01186_));
 sg13g2_a21oi_1 _07081_ (.A1(net1387),
    .A2(_01183_),
    .Y(_01237_),
    .B1(net1345));
 sg13g2_mux2_1 _07082_ (.A0(_01178_),
    .A1(_01185_),
    .S(net1387),
    .X(_01238_));
 sg13g2_nor2_1 _07083_ (.A(net1342),
    .B(_01238_),
    .Y(_01239_));
 sg13g2_a21o_1 _07084_ (.A2(_01237_),
    .A1(_01236_),
    .B1(net1431),
    .X(_01240_));
 sg13g2_nor3_1 _07085_ (.A(_01235_),
    .B(_01239_),
    .C(_01240_),
    .Y(_01241_));
 sg13g2_mux2_1 _07086_ (.A0(_01165_),
    .A1(_01168_),
    .S(net1450),
    .X(_01242_));
 sg13g2_nor2_1 _07087_ (.A(net1388),
    .B(_00507_),
    .Y(_01243_));
 sg13g2_a22oi_1 _07088_ (.Y(_01244_),
    .B1(_01243_),
    .B2(net1403),
    .A2(_01242_),
    .A1(net1388));
 sg13g2_nor2_1 _07089_ (.A(net1441),
    .B(_01244_),
    .Y(_01245_));
 sg13g2_a221oi_1 _07090_ (.B2(net1430),
    .C1(_01241_),
    .B1(_01245_),
    .A1(_01146_),
    .Y(_01246_),
    .A2(_01215_));
 sg13g2_nor2b_1 _07091_ (.A(_01218_),
    .B_N(_01219_),
    .Y(_01247_));
 sg13g2_nor2_1 _07092_ (.A(net1238),
    .B(_01247_),
    .Y(_01248_));
 sg13g2_xnor2_1 _07093_ (.Y(_01249_),
    .A(_01246_),
    .B(_01248_));
 sg13g2_nand2b_1 _07094_ (.Y(_01250_),
    .B(\cordic_inst.cordic_state[35] ),
    .A_N(_01249_));
 sg13g2_xnor2_1 _07095_ (.Y(_01251_),
    .A(_05584_),
    .B(_01249_));
 sg13g2_xnor2_1 _07096_ (.Y(_01252_),
    .A(_01231_),
    .B(_01251_));
 sg13g2_a22oi_1 _07097_ (.Y(_01253_),
    .B1(_00476_),
    .B2(net1541),
    .A2(net1368),
    .A1(net1627));
 sg13g2_o21ai_1 _07098_ (.B1(_01253_),
    .Y(_01254_),
    .A1(net1324),
    .A2(_01252_));
 sg13g2_a21oi_1 _07099_ (.A1(net1289),
    .A2(_01254_),
    .Y(_01255_),
    .B1(net1747));
 sg13g2_o21ai_1 _07100_ (.B1(_01255_),
    .Y(_00216_),
    .A1(_05584_),
    .A2(net1289));
 sg13g2_o21ai_1 _07101_ (.B1(_01250_),
    .Y(_01256_),
    .A1(_01231_),
    .A2(_01251_));
 sg13g2_mux2_1 _07102_ (.A0(_01137_),
    .A1(_01148_),
    .S(net1444),
    .X(_01257_));
 sg13g2_nor2_1 _07103_ (.A(_01136_),
    .B(net1342),
    .Y(_01258_));
 sg13g2_o21ai_1 _07104_ (.B1(net1396),
    .Y(_01259_),
    .A1(net1345),
    .A2(_01143_));
 sg13g2_nor2_1 _07105_ (.A(_01258_),
    .B(_01259_),
    .Y(_01260_));
 sg13g2_o21ai_1 _07106_ (.B1(_01260_),
    .Y(_01261_),
    .A1(net1393),
    .A2(_01257_));
 sg13g2_nand2b_2 _07107_ (.Y(_01262_),
    .B(net1346),
    .A_N(_00487_));
 sg13g2_nand2_1 _07108_ (.Y(_01263_),
    .A(net1346),
    .B(_01150_));
 sg13g2_o21ai_1 _07109_ (.B1(_01261_),
    .Y(_01264_),
    .A1(net1396),
    .A2(_01263_));
 sg13g2_a21oi_1 _07110_ (.A1(_01146_),
    .A2(_01262_),
    .Y(_01265_),
    .B1(_01264_));
 sg13g2_inv_1 _07111_ (.Y(_01266_),
    .A(_01265_));
 sg13g2_nand2_1 _07112_ (.Y(_01267_),
    .A(_01246_),
    .B(_01247_));
 sg13g2_nand2_1 _07113_ (.Y(_01268_),
    .A(net1244),
    .B(_01267_));
 sg13g2_xnor2_1 _07114_ (.Y(_01269_),
    .A(_01266_),
    .B(_01268_));
 sg13g2_nor2b_1 _07115_ (.A(_01269_),
    .B_N(\cordic_inst.cordic_state[36] ),
    .Y(_01270_));
 sg13g2_xnor2_1 _07116_ (.Y(_01271_),
    .A(\cordic_inst.cordic_state[36] ),
    .B(_01269_));
 sg13g2_and2_1 _07117_ (.A(_01256_),
    .B(_01271_),
    .X(_01272_));
 sg13g2_o21ai_1 _07118_ (.B1(net1280),
    .Y(_01273_),
    .A1(_01256_),
    .A2(_01271_));
 sg13g2_a21oi_1 _07119_ (.A1(net1531),
    .A2(net1476),
    .Y(_01274_),
    .B1(net1368));
 sg13g2_o21ai_1 _07120_ (.B1(_01274_),
    .Y(_01275_),
    .A1(_01272_),
    .A2(_01273_));
 sg13g2_a21oi_1 _07121_ (.A1(_05557_),
    .A2(net1368),
    .Y(_01276_),
    .B1(net1303));
 sg13g2_a22oi_1 _07122_ (.Y(_01277_),
    .B1(_01275_),
    .B2(_01276_),
    .A2(net1303),
    .A1(net742));
 sg13g2_nor2_1 _07123_ (.A(net1748),
    .B(_01277_),
    .Y(_00217_));
 sg13g2_a21oi_1 _07124_ (.A1(_01256_),
    .A2(_01271_),
    .Y(_01278_),
    .B1(_01270_));
 sg13g2_mux2_1 _07125_ (.A0(_01166_),
    .A1(_01177_),
    .S(_05590_),
    .X(_01279_));
 sg13g2_nor2_1 _07126_ (.A(net1393),
    .B(_01279_),
    .Y(_01280_));
 sg13g2_nor2_1 _07127_ (.A(net1342),
    .B(_01180_),
    .Y(_01281_));
 sg13g2_o21ai_1 _07128_ (.B1(net1396),
    .Y(_01282_),
    .A1(net1343),
    .A2(_01187_));
 sg13g2_nor3_1 _07129_ (.A(_01280_),
    .B(_01281_),
    .C(_01282_),
    .Y(_01283_));
 sg13g2_nor2_1 _07130_ (.A(net1343),
    .B(_01170_),
    .Y(_01284_));
 sg13g2_inv_1 _07131_ (.Y(_01285_),
    .A(_01284_));
 sg13g2_a221oi_1 _07132_ (.B2(net1431),
    .C1(_01283_),
    .B1(_01284_),
    .A1(_01146_),
    .Y(_01286_),
    .A2(_01262_));
 sg13g2_o21ai_1 _07133_ (.B1(net1244),
    .Y(_01287_),
    .A1(_01266_),
    .A2(_01267_));
 sg13g2_xnor2_1 _07134_ (.Y(_01288_),
    .A(_01286_),
    .B(_01287_));
 sg13g2_nand2_1 _07135_ (.Y(_01289_),
    .A(net1426),
    .B(_01288_));
 sg13g2_nor2_1 _07136_ (.A(net1426),
    .B(_01288_),
    .Y(_01290_));
 sg13g2_xnor2_1 _07137_ (.Y(_01291_),
    .A(net1426),
    .B(_01288_));
 sg13g2_xnor2_1 _07138_ (.Y(_01292_),
    .A(_01278_),
    .B(_01291_));
 sg13g2_a221oi_1 _07139_ (.B2(net1526),
    .C1(net1303),
    .B1(_00476_),
    .A1(net1615),
    .Y(_01293_),
    .A2(net1368));
 sg13g2_o21ai_1 _07140_ (.B1(_01293_),
    .Y(_01294_),
    .A1(net1324),
    .A2(_01292_));
 sg13g2_o21ai_1 _07141_ (.B1(_01294_),
    .Y(_01295_),
    .A1(net757),
    .A2(net1289));
 sg13g2_nand2_1 _07142_ (.Y(_00218_),
    .A(net1766),
    .B(_01295_));
 sg13g2_nand4_1 _07143_ (.B(_01247_),
    .C(_01265_),
    .A(_01246_),
    .Y(_01296_),
    .D(_01286_));
 sg13g2_nand2_1 _07144_ (.Y(_01297_),
    .A(net1242),
    .B(_01296_));
 sg13g2_mux2_1 _07145_ (.A0(_01203_),
    .A1(_01211_),
    .S(net1444),
    .X(_01298_));
 sg13g2_and2_1 _07146_ (.A(net1346),
    .B(_01208_),
    .X(_01299_));
 sg13g2_a221oi_1 _07147_ (.B2(net1439),
    .C1(_01299_),
    .B1(_01298_),
    .A1(_01141_),
    .Y(_01300_),
    .A2(_01204_));
 sg13g2_nor2_1 _07148_ (.A(net1343),
    .B(_01210_),
    .Y(_01301_));
 sg13g2_nand2_1 _07149_ (.Y(_01302_),
    .A(_00506_),
    .B(net1346));
 sg13g2_a22oi_1 _07150_ (.Y(_01303_),
    .B1(_01302_),
    .B2(_01146_),
    .A2(_01301_),
    .A1(net1429));
 sg13g2_o21ai_1 _07151_ (.B1(_01303_),
    .Y(_01304_),
    .A1(net1431),
    .A2(_01300_));
 sg13g2_xor2_1 _07152_ (.B(_01304_),
    .A(_01297_),
    .X(_01305_));
 sg13g2_and2_1 _07153_ (.A(net1425),
    .B(_01305_),
    .X(_01306_));
 sg13g2_xor2_1 _07154_ (.B(_01305_),
    .A(net1425),
    .X(_01307_));
 sg13g2_o21ai_1 _07155_ (.B1(_01289_),
    .Y(_01308_),
    .A1(_01278_),
    .A2(_01290_));
 sg13g2_nor2_1 _07156_ (.A(_01307_),
    .B(_01308_),
    .Y(_01309_));
 sg13g2_a21o_1 _07157_ (.A2(_01308_),
    .A1(_01307_),
    .B1(_00485_),
    .X(_01310_));
 sg13g2_a21oi_1 _07158_ (.A1(net1525),
    .A2(net1474),
    .Y(_01311_),
    .B1(net1362));
 sg13g2_o21ai_1 _07159_ (.B1(_01311_),
    .Y(_01312_),
    .A1(_01309_),
    .A2(_01310_));
 sg13g2_o21ai_1 _07160_ (.B1(_01312_),
    .Y(_01313_),
    .A1(net1611),
    .A2(net1371));
 sg13g2_o21ai_1 _07161_ (.B1(net1766),
    .Y(_01314_),
    .A1(net701),
    .A2(net1288));
 sg13g2_a21oi_1 _07162_ (.A1(net1289),
    .A2(_01313_),
    .Y(_00219_),
    .B1(_01314_));
 sg13g2_a21oi_1 _07163_ (.A1(_01307_),
    .A2(_01308_),
    .Y(_01315_),
    .B1(_01306_));
 sg13g2_mux2_1 _07164_ (.A0(_01232_),
    .A1(_01242_),
    .S(net1443),
    .X(_01316_));
 sg13g2_nor2_1 _07165_ (.A(net1393),
    .B(_01316_),
    .Y(_01317_));
 sg13g2_nor2_1 _07166_ (.A(net1342),
    .B(_01233_),
    .Y(_01318_));
 sg13g2_o21ai_1 _07167_ (.B1(net1396),
    .Y(_01319_),
    .A1(net1343),
    .A2(_01238_));
 sg13g2_nor3_1 _07168_ (.A(_01317_),
    .B(_01318_),
    .C(_01319_),
    .Y(_01320_));
 sg13g2_nor2_1 _07169_ (.A(_01146_),
    .B(_01320_),
    .Y(_01321_));
 sg13g2_nor2_1 _07170_ (.A(_01296_),
    .B(_01304_),
    .Y(_01322_));
 sg13g2_nor2_1 _07171_ (.A(net1240),
    .B(_01322_),
    .Y(_01323_));
 sg13g2_xor2_1 _07172_ (.B(_01323_),
    .A(_01321_),
    .X(_01324_));
 sg13g2_nand2_1 _07173_ (.Y(_01325_),
    .A(net1424),
    .B(_01324_));
 sg13g2_xnor2_1 _07174_ (.Y(_01326_),
    .A(net1424),
    .B(_01324_));
 sg13g2_xnor2_1 _07175_ (.Y(_01327_),
    .A(_01315_),
    .B(_01326_));
 sg13g2_nand2_1 _07176_ (.Y(_01328_),
    .A(net1348),
    .B(_01327_));
 sg13g2_a221oi_1 _07177_ (.B2(_01328_),
    .C1(net1366),
    .B1(net1359),
    .A1(net1518),
    .Y(_01329_),
    .A2(net1477));
 sg13g2_o21ai_1 _07178_ (.B1(net1290),
    .Y(_01330_),
    .A1(net1606),
    .A2(net1371));
 sg13g2_a21oi_1 _07179_ (.A1(net1424),
    .A2(net1302),
    .Y(_01331_),
    .B1(net1748));
 sg13g2_o21ai_1 _07180_ (.B1(_01331_),
    .Y(_00220_),
    .A1(_01329_),
    .A2(_01330_));
 sg13g2_o21ai_1 _07181_ (.B1(_01325_),
    .Y(_01332_),
    .A1(_01315_),
    .A2(_01326_));
 sg13g2_and2_1 _07182_ (.A(_01321_),
    .B(_01322_),
    .X(_01333_));
 sg13g2_nor2_1 _07183_ (.A(net1236),
    .B(_01333_),
    .Y(_01334_));
 sg13g2_o21ai_1 _07184_ (.B1(net1396),
    .Y(_01335_),
    .A1(net1439),
    .A2(_01138_));
 sg13g2_a21oi_1 _07185_ (.A1(net1439),
    .A2(_01152_),
    .Y(_01336_),
    .B1(_01335_));
 sg13g2_nor2_2 _07186_ (.A(_01146_),
    .B(_01336_),
    .Y(_01337_));
 sg13g2_xnor2_1 _07187_ (.Y(_01338_),
    .A(_01334_),
    .B(_01337_));
 sg13g2_nor2b_1 _07188_ (.A(_01338_),
    .B_N(net1423),
    .Y(_01339_));
 sg13g2_xnor2_1 _07189_ (.Y(_01340_),
    .A(net1423),
    .B(_01338_));
 sg13g2_and2_1 _07190_ (.A(_01332_),
    .B(_01340_),
    .X(_01341_));
 sg13g2_o21ai_1 _07191_ (.B1(net1282),
    .Y(_01342_),
    .A1(_01332_),
    .A2(_01340_));
 sg13g2_a21oi_1 _07192_ (.A1(net1733),
    .A2(net1474),
    .Y(_01343_),
    .B1(net1361));
 sg13g2_o21ai_1 _07193_ (.B1(_01343_),
    .Y(_01344_),
    .A1(_01341_),
    .A2(_01342_));
 sg13g2_o21ai_1 _07194_ (.B1(_01344_),
    .Y(_01345_),
    .A1(net1602),
    .A2(net1370));
 sg13g2_o21ai_1 _07195_ (.B1(net1765),
    .Y(_01346_),
    .A1(net1423),
    .A2(net1287));
 sg13g2_a21oi_1 _07196_ (.A1(net1287),
    .A2(_01345_),
    .Y(_00221_),
    .B1(_01346_));
 sg13g2_a21oi_1 _07197_ (.A1(_01332_),
    .A2(_01340_),
    .Y(_01347_),
    .B1(_01339_));
 sg13g2_a21oi_2 _07198_ (.B1(net1428),
    .Y(_01348_),
    .A2(net1442),
    .A1(net1437));
 sg13g2_a21oi_1 _07199_ (.A1(net1397),
    .A2(net1385),
    .Y(_01349_),
    .B1(_01348_));
 sg13g2_nand2_1 _07200_ (.Y(_01350_),
    .A(net1403),
    .B(_01349_));
 sg13g2_a21oi_1 _07201_ (.A1(net1435),
    .A2(_01172_),
    .Y(_01351_),
    .B1(net1428));
 sg13g2_o21ai_1 _07202_ (.B1(_01351_),
    .Y(_01352_),
    .A1(net1435),
    .A2(_01181_));
 sg13g2_nand2_1 _07203_ (.Y(_01353_),
    .A(_01350_),
    .B(_01352_));
 sg13g2_inv_1 _07204_ (.Y(_01354_),
    .A(_01353_));
 sg13g2_a21oi_1 _07205_ (.A1(_01333_),
    .A2(_01337_),
    .Y(_01355_),
    .B1(net1236));
 sg13g2_xnor2_1 _07206_ (.Y(_01356_),
    .A(_01354_),
    .B(_01355_));
 sg13g2_nand2b_1 _07207_ (.Y(_01357_),
    .B(net1422),
    .A_N(_01356_));
 sg13g2_xor2_1 _07208_ (.B(_01356_),
    .A(net1422),
    .X(_01358_));
 sg13g2_xnor2_1 _07209_ (.Y(_01359_),
    .A(_01347_),
    .B(_01358_));
 sg13g2_nand2_1 _07210_ (.Y(_01360_),
    .A(net688),
    .B(net1296));
 sg13g2_a22oi_1 _07211_ (.Y(_01361_),
    .B1(net1322),
    .B2(net1727),
    .A2(net1361),
    .A1(net1597));
 sg13g2_o21ai_1 _07212_ (.B1(_01361_),
    .Y(_01362_),
    .A1(net1323),
    .A2(_01359_));
 sg13g2_nand2_1 _07213_ (.Y(_01363_),
    .A(net1287),
    .B(_01362_));
 sg13g2_nand3_1 _07214_ (.B(_01360_),
    .C(_01363_),
    .A(net1765),
    .Y(_00222_));
 sg13g2_o21ai_1 _07215_ (.B1(_01357_),
    .Y(_01364_),
    .A1(_01347_),
    .A2(_01358_));
 sg13g2_nor2_1 _07216_ (.A(net1439),
    .B(_01205_),
    .Y(_01365_));
 sg13g2_nor2_1 _07217_ (.A(net1429),
    .B(_01365_),
    .Y(_01366_));
 sg13g2_o21ai_1 _07218_ (.B1(_01366_),
    .Y(_01367_),
    .A1(net1392),
    .A2(_01213_));
 sg13g2_nand2_1 _07219_ (.Y(_01368_),
    .A(_01350_),
    .B(_01367_));
 sg13g2_and2_1 _07220_ (.A(_01337_),
    .B(_01354_),
    .X(_01369_));
 sg13g2_a21oi_1 _07221_ (.A1(_01333_),
    .A2(_01369_),
    .Y(_01370_),
    .B1(net1236));
 sg13g2_xor2_1 _07222_ (.B(_01370_),
    .A(_01368_),
    .X(_01371_));
 sg13g2_nor2b_1 _07223_ (.A(_01371_),
    .B_N(net1421),
    .Y(_01372_));
 sg13g2_xnor2_1 _07224_ (.Y(_01373_),
    .A(net1421),
    .B(_01371_));
 sg13g2_o21ai_1 _07225_ (.B1(net1282),
    .Y(_01374_),
    .A1(_01364_),
    .A2(_01373_));
 sg13g2_a21o_1 _07226_ (.A2(_01373_),
    .A1(_01364_),
    .B1(_01374_),
    .X(_01375_));
 sg13g2_a21oi_1 _07227_ (.A1(net1720),
    .A2(net1474),
    .Y(_01376_),
    .B1(net1361));
 sg13g2_o21ai_1 _07228_ (.B1(net1287),
    .Y(_01377_),
    .A1(net1590),
    .A2(net1370));
 sg13g2_a21oi_1 _07229_ (.A1(_01375_),
    .A2(_01376_),
    .Y(_01378_),
    .B1(_01377_));
 sg13g2_a21oi_1 _07230_ (.A1(net1421),
    .A2(net1296),
    .Y(_01379_),
    .B1(_01378_));
 sg13g2_nor2_1 _07231_ (.A(net1746),
    .B(net799),
    .Y(_00223_));
 sg13g2_a21oi_1 _07232_ (.A1(_01364_),
    .A2(_01373_),
    .Y(_01380_),
    .B1(_01372_));
 sg13g2_nor2_1 _07233_ (.A(net1428),
    .B(_00507_),
    .Y(_01381_));
 sg13g2_nor2_1 _07234_ (.A(_01348_),
    .B(_01381_),
    .Y(_01382_));
 sg13g2_nand2_1 _07235_ (.Y(_01383_),
    .A(net1403),
    .B(_01382_));
 sg13g2_a21oi_1 _07236_ (.A1(net1436),
    .A2(_01244_),
    .Y(_01384_),
    .B1(net1428));
 sg13g2_o21ai_1 _07237_ (.B1(_01384_),
    .Y(_01385_),
    .A1(net1435),
    .A2(_01234_));
 sg13g2_nand2_1 _07238_ (.Y(_01386_),
    .A(_01383_),
    .B(_01385_));
 sg13g2_nand3_1 _07239_ (.B(_01367_),
    .C(_01369_),
    .A(_01333_),
    .Y(_01387_));
 sg13g2_nand2_1 _07240_ (.Y(_01388_),
    .A(net1241),
    .B(_01387_));
 sg13g2_xor2_1 _07241_ (.B(_01388_),
    .A(_01386_),
    .X(_01389_));
 sg13g2_nor2_1 _07242_ (.A(net1420),
    .B(_01389_),
    .Y(_01390_));
 sg13g2_xor2_1 _07243_ (.B(_01389_),
    .A(net1420),
    .X(_01391_));
 sg13g2_o21ai_1 _07244_ (.B1(net1348),
    .Y(_01392_),
    .A1(_01380_),
    .A2(_01391_));
 sg13g2_a21oi_1 _07245_ (.A1(_01380_),
    .A2(_01391_),
    .Y(_01393_),
    .B1(_01392_));
 sg13g2_a22oi_1 _07246_ (.Y(_01394_),
    .B1(net1322),
    .B2(net1714),
    .A2(net1361),
    .A1(net1583));
 sg13g2_o21ai_1 _07247_ (.B1(_01394_),
    .Y(_01395_),
    .A1(net1323),
    .A2(_01393_));
 sg13g2_o21ai_1 _07248_ (.B1(_01395_),
    .Y(_01396_),
    .A1(net732),
    .A2(net1287));
 sg13g2_nand2_1 _07249_ (.Y(_00224_),
    .A(net1765),
    .B(_01396_));
 sg13g2_a21oi_1 _07250_ (.A1(net1438),
    .A2(_00495_),
    .Y(_01397_),
    .B1(net1427));
 sg13g2_nor2_1 _07251_ (.A(_05576_),
    .B(_01397_),
    .Y(_01398_));
 sg13g2_mux2_1 _07252_ (.A0(_01150_),
    .A1(_01257_),
    .S(net1393),
    .X(_01399_));
 sg13g2_a21o_1 _07253_ (.A2(_01399_),
    .A1(_01348_),
    .B1(_01398_),
    .X(_01400_));
 sg13g2_inv_1 _07254_ (.Y(_01401_),
    .A(_01400_));
 sg13g2_o21ai_1 _07255_ (.B1(net1241),
    .Y(_01402_),
    .A1(_01386_),
    .A2(_01387_));
 sg13g2_xnor2_1 _07256_ (.Y(_01403_),
    .A(_01401_),
    .B(_01402_));
 sg13g2_and2_1 _07257_ (.A(net1419),
    .B(_01403_),
    .X(_01404_));
 sg13g2_xor2_1 _07258_ (.B(_01403_),
    .A(net1419),
    .X(_01405_));
 sg13g2_a221oi_1 _07259_ (.B2(net1420),
    .C1(_01372_),
    .B1(_01389_),
    .A1(_01364_),
    .Y(_01406_),
    .A2(_01373_));
 sg13g2_nor2_1 _07260_ (.A(_01390_),
    .B(_01406_),
    .Y(_01407_));
 sg13g2_and2_1 _07261_ (.A(_01405_),
    .B(_01407_),
    .X(_01408_));
 sg13g2_or2_1 _07262_ (.X(_01409_),
    .B(_01407_),
    .A(_01405_));
 sg13g2_nand3b_1 _07263_ (.B(_01409_),
    .C(net1282),
    .Y(_01410_),
    .A_N(_01408_));
 sg13g2_a21oi_1 _07264_ (.A1(net1709),
    .A2(net1479),
    .Y(_01411_),
    .B1(net1361));
 sg13g2_o21ai_1 _07265_ (.B1(net1287),
    .Y(_01412_),
    .A1(net1578),
    .A2(net1370));
 sg13g2_a21oi_1 _07266_ (.A1(_01410_),
    .A2(_01411_),
    .Y(_01413_),
    .B1(_01412_));
 sg13g2_a21oi_1 _07267_ (.A1(net1419),
    .A2(net1296),
    .Y(_01414_),
    .B1(_01413_));
 sg13g2_nor2_1 _07268_ (.A(net1746),
    .B(net803),
    .Y(_00225_));
 sg13g2_nor2_1 _07269_ (.A(_01404_),
    .B(_01408_),
    .Y(_01415_));
 sg13g2_o21ai_1 _07270_ (.B1(_01348_),
    .Y(_01416_),
    .A1(net1435),
    .A2(_01279_));
 sg13g2_a21o_1 _07271_ (.A2(_01170_),
    .A1(net1435),
    .B1(_01416_),
    .X(_01417_));
 sg13g2_nand2b_1 _07272_ (.Y(_01418_),
    .B(_01417_),
    .A_N(_01398_));
 sg13g2_o21ai_1 _07273_ (.B1(_01402_),
    .Y(_01419_),
    .A1(net1236),
    .A2(_01401_));
 sg13g2_xnor2_1 _07274_ (.Y(_01420_),
    .A(_01418_),
    .B(_01419_));
 sg13g2_nor2_1 _07275_ (.A(net1418),
    .B(_01420_),
    .Y(_01421_));
 sg13g2_xor2_1 _07276_ (.B(_01420_),
    .A(net1418),
    .X(_01422_));
 sg13g2_o21ai_1 _07277_ (.B1(net1348),
    .Y(_01423_),
    .A1(_01415_),
    .A2(_01422_));
 sg13g2_a21oi_1 _07278_ (.A1(_01415_),
    .A2(_01422_),
    .Y(_01424_),
    .B1(_01423_));
 sg13g2_a22oi_1 _07279_ (.Y(_01425_),
    .B1(net1322),
    .B2(net1703),
    .A2(net1361),
    .A1(net1573));
 sg13g2_o21ai_1 _07280_ (.B1(_01425_),
    .Y(_01426_),
    .A1(net1323),
    .A2(_01424_));
 sg13g2_o21ai_1 _07281_ (.B1(_01426_),
    .Y(_01427_),
    .A1(net743),
    .A2(net1287));
 sg13g2_nand2_1 _07282_ (.Y(_00226_),
    .A(net1765),
    .B(_01427_));
 sg13g2_o21ai_1 _07283_ (.B1(_01348_),
    .Y(_01428_),
    .A1(net1391),
    .A2(_00506_));
 sg13g2_nand2_1 _07284_ (.Y(_01429_),
    .A(net1403),
    .B(_01428_));
 sg13g2_a21oi_1 _07285_ (.A1(net1385),
    .A2(_01149_),
    .Y(_01430_),
    .B1(net1390));
 sg13g2_o21ai_1 _07286_ (.B1(_01348_),
    .Y(_01431_),
    .A1(net1435),
    .A2(_01298_));
 sg13g2_o21ai_1 _07287_ (.B1(_01429_),
    .Y(_01432_),
    .A1(_01430_),
    .A2(_01431_));
 sg13g2_nor2_1 _07288_ (.A(net1236),
    .B(_01417_),
    .Y(_01433_));
 sg13g2_nor2_1 _07289_ (.A(_01419_),
    .B(_01433_),
    .Y(_01434_));
 sg13g2_xor2_1 _07290_ (.B(_01434_),
    .A(_01432_),
    .X(_01435_));
 sg13g2_and2_1 _07291_ (.A(net1417),
    .B(_01435_),
    .X(_01436_));
 sg13g2_xor2_1 _07292_ (.B(_01435_),
    .A(net1417),
    .X(_01437_));
 sg13g2_a221oi_1 _07293_ (.B2(net1418),
    .C1(_01404_),
    .B1(_01420_),
    .A1(_01405_),
    .Y(_01438_),
    .A2(_01407_));
 sg13g2_nor2_1 _07294_ (.A(_01421_),
    .B(_01438_),
    .Y(_01439_));
 sg13g2_and2_1 _07295_ (.A(_01437_),
    .B(_01439_),
    .X(_01440_));
 sg13g2_o21ai_1 _07296_ (.B1(net1282),
    .Y(_01441_),
    .A1(_01437_),
    .A2(_01439_));
 sg13g2_a21oi_1 _07297_ (.A1(net1698),
    .A2(net1474),
    .Y(_01442_),
    .B1(net1361));
 sg13g2_o21ai_1 _07298_ (.B1(_01442_),
    .Y(_01443_),
    .A1(_01440_),
    .A2(_01441_));
 sg13g2_a21oi_1 _07299_ (.A1(_05555_),
    .A2(net1361),
    .Y(_01444_),
    .B1(net1305));
 sg13g2_a22oi_1 _07300_ (.Y(_01445_),
    .B1(_01443_),
    .B2(_01444_),
    .A2(net1305),
    .A1(net1417));
 sg13g2_nor2_1 _07301_ (.A(net1746),
    .B(_01445_),
    .Y(_00227_));
 sg13g2_a21o_1 _07302_ (.A2(_01439_),
    .A1(_01437_),
    .B1(_01436_),
    .X(_01446_));
 sg13g2_nor3_1 _07303_ (.A(net1391),
    .B(net1443),
    .C(_00507_),
    .Y(_01447_));
 sg13g2_a22oi_1 _07304_ (.Y(_01448_),
    .B1(_01447_),
    .B2(net1403),
    .A2(_01316_),
    .A1(net1391));
 sg13g2_o21ai_1 _07305_ (.B1(_01429_),
    .Y(_01449_),
    .A1(net1427),
    .A2(_01448_));
 sg13g2_nand2_1 _07306_ (.Y(_01450_),
    .A(net1241),
    .B(_01432_));
 sg13g2_and2_1 _07307_ (.A(_01434_),
    .B(_01450_),
    .X(_01451_));
 sg13g2_xnor2_1 _07308_ (.Y(_01452_),
    .A(_01449_),
    .B(_01451_));
 sg13g2_nor2b_1 _07309_ (.A(_01452_),
    .B_N(net1416),
    .Y(_01453_));
 sg13g2_xnor2_1 _07310_ (.Y(_01454_),
    .A(net1416),
    .B(_01452_));
 sg13g2_xnor2_1 _07311_ (.Y(_01455_),
    .A(_01446_),
    .B(_01454_));
 sg13g2_a22oi_1 _07312_ (.Y(_01456_),
    .B1(net1322),
    .B2(net1693),
    .A2(net1362),
    .A1(net1565));
 sg13g2_o21ai_1 _07313_ (.B1(_01456_),
    .Y(_01457_),
    .A1(net1324),
    .A2(_01455_));
 sg13g2_mux2_1 _07314_ (.A0(net1416),
    .A1(_01457_),
    .S(net1287),
    .X(_01458_));
 sg13g2_nand2b_1 _07315_ (.Y(_00228_),
    .B(net1765),
    .A_N(_01458_));
 sg13g2_a21o_1 _07316_ (.A2(_01454_),
    .A1(_01446_),
    .B1(_01453_),
    .X(_01459_));
 sg13g2_o21ai_1 _07317_ (.B1(net1403),
    .Y(_01460_),
    .A1(net1430),
    .A2(_00499_));
 sg13g2_o21ai_1 _07318_ (.B1(_01460_),
    .Y(_01461_),
    .A1(net1430),
    .A2(_01153_));
 sg13g2_nand2_1 _07319_ (.Y(_01462_),
    .A(net1241),
    .B(_01449_));
 sg13g2_nand2_1 _07320_ (.Y(_01463_),
    .A(_01451_),
    .B(_01462_));
 sg13g2_xnor2_1 _07321_ (.Y(_01464_),
    .A(_01461_),
    .B(_01463_));
 sg13g2_and2_1 _07322_ (.A(net1415),
    .B(_01464_),
    .X(_01465_));
 sg13g2_xor2_1 _07323_ (.B(_01464_),
    .A(net1415),
    .X(_01466_));
 sg13g2_and2_1 _07324_ (.A(_01459_),
    .B(_01466_),
    .X(_01467_));
 sg13g2_o21ai_1 _07325_ (.B1(net1282),
    .Y(_01468_),
    .A1(_01459_),
    .A2(_01466_));
 sg13g2_a21oi_2 _07326_ (.B1(net1367),
    .Y(_01469_),
    .A2(net1477),
    .A1(net1685));
 sg13g2_o21ai_1 _07327_ (.B1(_01469_),
    .Y(_01470_),
    .A1(_01467_),
    .A2(_01468_));
 sg13g2_a21oi_1 _07328_ (.A1(_05554_),
    .A2(net1362),
    .Y(_01471_),
    .B1(net1296));
 sg13g2_a22oi_1 _07329_ (.Y(_01472_),
    .B1(_01470_),
    .B2(_01471_),
    .A2(net1305),
    .A1(net677));
 sg13g2_nor2_1 _07330_ (.A(net1746),
    .B(_01472_),
    .Y(_00229_));
 sg13g2_or2_1 _07331_ (.X(_01473_),
    .B(_01467_),
    .A(_01465_));
 sg13g2_o21ai_1 _07332_ (.B1(_01460_),
    .Y(_01474_),
    .A1(net1430),
    .A2(_01173_));
 sg13g2_a21o_1 _07333_ (.A2(_01461_),
    .A1(net1242),
    .B1(_01463_),
    .X(_01475_));
 sg13g2_xnor2_1 _07334_ (.Y(_01476_),
    .A(_01474_),
    .B(_01475_));
 sg13g2_or2_1 _07335_ (.X(_01477_),
    .B(_01476_),
    .A(\cordic_inst.cordic_state[49] ));
 sg13g2_inv_1 _07336_ (.Y(_01478_),
    .A(_01477_));
 sg13g2_xnor2_1 _07337_ (.Y(_01479_),
    .A(_05583_),
    .B(_01476_));
 sg13g2_xnor2_1 _07338_ (.Y(_01480_),
    .A(_01473_),
    .B(_01479_));
 sg13g2_a22oi_1 _07339_ (.Y(_01481_),
    .B1(net1321),
    .B2(net1679),
    .A2(net1367),
    .A1(net1507));
 sg13g2_o21ai_1 _07340_ (.B1(_01481_),
    .Y(_01482_),
    .A1(net1324),
    .A2(_01480_));
 sg13g2_a21oi_1 _07341_ (.A1(net1288),
    .A2(_01482_),
    .Y(_01483_),
    .B1(net1746));
 sg13g2_o21ai_1 _07342_ (.B1(_01483_),
    .Y(_00230_),
    .A1(_05583_),
    .A2(net1288));
 sg13g2_nor2_1 _07343_ (.A(net1430),
    .B(_01215_),
    .Y(_01484_));
 sg13g2_inv_1 _07344_ (.Y(_01485_),
    .A(_01484_));
 sg13g2_a22oi_1 _07345_ (.Y(_01486_),
    .B1(_01485_),
    .B2(net1403),
    .A2(_01214_),
    .A1(net1394));
 sg13g2_a21oi_1 _07346_ (.A1(net1242),
    .A2(_01474_),
    .Y(_01487_),
    .B1(_01475_));
 sg13g2_xnor2_1 _07347_ (.Y(_01488_),
    .A(_01486_),
    .B(_01487_));
 sg13g2_nand2_1 _07348_ (.Y(_01489_),
    .A(net1414),
    .B(_01488_));
 sg13g2_xor2_1 _07349_ (.B(_01488_),
    .A(net1414),
    .X(_01490_));
 sg13g2_inv_1 _07350_ (.Y(_01491_),
    .A(_01490_));
 sg13g2_a221oi_1 _07351_ (.B2(\cordic_inst.cordic_state[49] ),
    .C1(_01465_),
    .B1(_01476_),
    .A1(_01459_),
    .Y(_01492_),
    .A2(_01466_));
 sg13g2_or3_1 _07352_ (.A(_01478_),
    .B(_01491_),
    .C(_01492_),
    .X(_01493_));
 sg13g2_o21ai_1 _07353_ (.B1(_01491_),
    .Y(_01494_),
    .A1(_01478_),
    .A2(_01492_));
 sg13g2_nand3_1 _07354_ (.B(_01493_),
    .C(_01494_),
    .A(net1282),
    .Y(_01495_));
 sg13g2_a21oi_1 _07355_ (.A1(net1674),
    .A2(net1479),
    .Y(_01496_),
    .B1(net1362));
 sg13g2_nand2_1 _07356_ (.Y(_01497_),
    .A(_01495_),
    .B(_01496_));
 sg13g2_o21ai_1 _07357_ (.B1(_01497_),
    .Y(_01498_),
    .A1(net1506),
    .A2(net1370));
 sg13g2_o21ai_1 _07358_ (.B1(net1765),
    .Y(_01499_),
    .A1(net705),
    .A2(net1288));
 sg13g2_a21oi_1 _07359_ (.A1(net1288),
    .A2(_01498_),
    .Y(_00231_),
    .B1(_01499_));
 sg13g2_nand2_1 _07360_ (.Y(_01500_),
    .A(net1394),
    .B(_01245_));
 sg13g2_o21ai_1 _07361_ (.B1(_01500_),
    .Y(_01501_),
    .A1(_05576_),
    .A2(_01484_));
 sg13g2_a21o_1 _07362_ (.A2(_01487_),
    .A1(_01486_),
    .B1(net1240),
    .X(_01502_));
 sg13g2_xnor2_1 _07363_ (.Y(_01503_),
    .A(_01501_),
    .B(_01502_));
 sg13g2_nand2b_1 _07364_ (.Y(_01504_),
    .B(\cordic_inst.cordic_state[51] ),
    .A_N(_01503_));
 sg13g2_xnor2_1 _07365_ (.Y(_01505_),
    .A(_05582_),
    .B(_01503_));
 sg13g2_nand2_1 _07366_ (.Y(_01506_),
    .A(_01489_),
    .B(_01493_));
 sg13g2_o21ai_1 _07367_ (.B1(net1348),
    .Y(_01507_),
    .A1(_01505_),
    .A2(_01506_));
 sg13g2_a21oi_1 _07368_ (.A1(_01505_),
    .A2(_01506_),
    .Y(_01508_),
    .B1(_01507_));
 sg13g2_nand2b_1 _07369_ (.Y(_01509_),
    .B(net1359),
    .A_N(_01508_));
 sg13g2_a21oi_1 _07370_ (.A1(net1670),
    .A2(net1476),
    .Y(_01510_),
    .B1(net1362));
 sg13g2_o21ai_1 _07371_ (.B1(net1288),
    .Y(_01511_),
    .A1(net1502),
    .A2(net1370));
 sg13g2_a21oi_1 _07372_ (.A1(_01509_),
    .A2(_01510_),
    .Y(_01512_),
    .B1(_01511_));
 sg13g2_a21oi_1 _07373_ (.A1(net758),
    .A2(net1296),
    .Y(_01513_),
    .B1(_01512_));
 sg13g2_nand2_1 _07374_ (.Y(_00232_),
    .A(net1765),
    .B(net759));
 sg13g2_o21ai_1 _07375_ (.B1(net1405),
    .Y(_01514_),
    .A1(net1433),
    .A2(_01262_));
 sg13g2_o21ai_1 _07376_ (.B1(_01514_),
    .Y(_01515_),
    .A1(net1433),
    .A2(_01263_));
 sg13g2_o21ai_1 _07377_ (.B1(_01502_),
    .Y(_01516_),
    .A1(net1237),
    .A2(_01500_));
 sg13g2_or2_1 _07378_ (.X(_01517_),
    .B(_01516_),
    .A(_01515_));
 sg13g2_xnor2_1 _07379_ (.Y(_01518_),
    .A(_01515_),
    .B(_01516_));
 sg13g2_nand2_1 _07380_ (.Y(_01519_),
    .A(net1413),
    .B(_01518_));
 sg13g2_xor2_1 _07381_ (.B(_01518_),
    .A(net1413),
    .X(_01520_));
 sg13g2_and2_1 _07382_ (.A(_01489_),
    .B(_01504_),
    .X(_01521_));
 sg13g2_a22oi_1 _07383_ (.Y(_01522_),
    .B1(_01521_),
    .B2(_01493_),
    .A2(_01503_),
    .A1(_05582_));
 sg13g2_nand2_1 _07384_ (.Y(_01523_),
    .A(_01520_),
    .B(_01522_));
 sg13g2_o21ai_1 _07385_ (.B1(net1281),
    .Y(_01524_),
    .A1(_01520_),
    .A2(_01522_));
 sg13g2_nand2b_1 _07386_ (.Y(_01525_),
    .B(_01523_),
    .A_N(_01524_));
 sg13g2_a21oi_1 _07387_ (.A1(net1666),
    .A2(net1477),
    .Y(_01526_),
    .B1(net1366));
 sg13g2_o21ai_1 _07388_ (.B1(net1290),
    .Y(_01527_),
    .A1(net1497),
    .A2(net1371));
 sg13g2_a21oi_1 _07389_ (.A1(_01525_),
    .A2(_01526_),
    .Y(_01528_),
    .B1(_01527_));
 sg13g2_a21oi_1 _07390_ (.A1(net627),
    .A2(net1302),
    .Y(_01529_),
    .B1(_01528_));
 sg13g2_nor2_1 _07391_ (.A(net1749),
    .B(_01529_),
    .Y(_00233_));
 sg13g2_and2_1 _07392_ (.A(_01519_),
    .B(_01523_),
    .X(_01530_));
 sg13g2_nor2_1 _07393_ (.A(net1433),
    .B(_01285_),
    .Y(_01531_));
 sg13g2_o21ai_1 _07394_ (.B1(_01514_),
    .Y(_01532_),
    .A1(net1433),
    .A2(_01285_));
 sg13g2_nand2_1 _07395_ (.Y(_01533_),
    .A(net1245),
    .B(_01517_));
 sg13g2_xor2_1 _07396_ (.B(_01533_),
    .A(_01532_),
    .X(_01534_));
 sg13g2_nor2_1 _07397_ (.A(net1412),
    .B(_01534_),
    .Y(_01535_));
 sg13g2_nand2_1 _07398_ (.Y(_01536_),
    .A(\cordic_inst.cordic_state[53] ),
    .B(_01534_));
 sg13g2_nor2b_1 _07399_ (.A(_01535_),
    .B_N(_01536_),
    .Y(_01537_));
 sg13g2_and2_1 _07400_ (.A(_01519_),
    .B(_01536_),
    .X(_01538_));
 sg13g2_and2_1 _07401_ (.A(_01530_),
    .B(_01537_),
    .X(_01539_));
 sg13g2_o21ai_1 _07402_ (.B1(net1348),
    .Y(_01540_),
    .A1(_01530_),
    .A2(_01537_));
 sg13g2_o21ai_1 _07403_ (.B1(_00462_),
    .Y(_01541_),
    .A1(_01539_),
    .A2(_01540_));
 sg13g2_a21oi_1 _07404_ (.A1(net1662),
    .A2(net1476),
    .Y(_01542_),
    .B1(net1366));
 sg13g2_nand2_1 _07405_ (.Y(_01543_),
    .A(_01541_),
    .B(_01542_));
 sg13g2_a21oi_1 _07406_ (.A1(_05553_),
    .A2(net1367),
    .Y(_01544_),
    .B1(net1301));
 sg13g2_a22oi_1 _07407_ (.Y(_01545_),
    .B1(_01543_),
    .B2(_01544_),
    .A2(net1300),
    .A1(net1412));
 sg13g2_nand2_1 _07408_ (.Y(_00234_),
    .A(net1780),
    .B(_01545_));
 sg13g2_a21oi_1 _07409_ (.A1(net1346),
    .A2(_01381_),
    .Y(_01546_),
    .B1(_05576_));
 sg13g2_a21o_1 _07410_ (.A2(_01301_),
    .A1(net1394),
    .B1(_01546_),
    .X(_01547_));
 sg13g2_inv_1 _07411_ (.Y(_01548_),
    .A(_01547_));
 sg13g2_o21ai_1 _07412_ (.B1(net1245),
    .Y(_01549_),
    .A1(_01517_),
    .A2(_01531_));
 sg13g2_xnor2_1 _07413_ (.Y(_01550_),
    .A(_01548_),
    .B(_01549_));
 sg13g2_xor2_1 _07414_ (.B(_01550_),
    .A(net1411),
    .X(_01551_));
 sg13g2_a21oi_1 _07415_ (.A1(_01523_),
    .A2(_01538_),
    .Y(_01552_),
    .B1(_01535_));
 sg13g2_and2_1 _07416_ (.A(_01551_),
    .B(_01552_),
    .X(_01553_));
 sg13g2_o21ai_1 _07417_ (.B1(net1281),
    .Y(_01554_),
    .A1(_01551_),
    .A2(_01552_));
 sg13g2_a21oi_1 _07418_ (.A1(net1658),
    .A2(net1477),
    .Y(_01555_),
    .B1(net1366));
 sg13g2_o21ai_1 _07419_ (.B1(_01555_),
    .Y(_01556_),
    .A1(_01553_),
    .A2(_01554_));
 sg13g2_a21oi_1 _07420_ (.A1(_05552_),
    .A2(net1366),
    .Y(_01557_),
    .B1(net1301));
 sg13g2_a22oi_1 _07421_ (.Y(_01558_),
    .B1(_01556_),
    .B2(_01557_),
    .A2(net1300),
    .A1(net1411));
 sg13g2_nor2_1 _07422_ (.A(net1748),
    .B(_01558_),
    .Y(_00235_));
 sg13g2_a21oi_1 _07423_ (.A1(net1411),
    .A2(_01550_),
    .Y(_01559_),
    .B1(_01553_));
 sg13g2_a21oi_1 _07424_ (.A1(_01548_),
    .A2(_01549_),
    .Y(_01560_),
    .B1(net1238));
 sg13g2_xor2_1 _07425_ (.B(net1410),
    .A(net1405),
    .X(_01561_));
 sg13g2_xor2_1 _07426_ (.B(_01561_),
    .A(_01560_),
    .X(_01562_));
 sg13g2_inv_1 _07427_ (.Y(_01563_),
    .A(_01562_));
 sg13g2_nand2b_1 _07428_ (.Y(_01564_),
    .B(_01562_),
    .A_N(_01559_));
 sg13g2_a21oi_1 _07429_ (.A1(_01559_),
    .A2(_01563_),
    .Y(_01565_),
    .B1(_00479_));
 sg13g2_a21oi_1 _07430_ (.A1(_01564_),
    .A2(_01565_),
    .Y(_01566_),
    .B1(_00464_));
 sg13g2_a221oi_1 _07431_ (.B2(net1656),
    .C1(_01566_),
    .B1(net1321),
    .A1(net1486),
    .Y(_01567_),
    .A2(net1369));
 sg13g2_a21oi_1 _07432_ (.A1(net1410),
    .A2(net1300),
    .Y(_01568_),
    .B1(net1749));
 sg13g2_o21ai_1 _07433_ (.B1(_01568_),
    .Y(_00236_),
    .A1(net1300),
    .A2(_01567_));
 sg13g2_mux4_1 _07434_ (.S0(net1454),
    .A0(net1423),
    .A1(net1422),
    .A2(net1421),
    .A3(net1420),
    .S1(net1448),
    .X(_01569_));
 sg13g2_mux4_1 _07435_ (.S0(net1454),
    .A0(net1419),
    .A1(net1418),
    .A2(net1417),
    .A3(net1416),
    .S1(net1447),
    .X(_01570_));
 sg13g2_mux2_1 _07436_ (.A0(_01569_),
    .A1(_01570_),
    .S(net1445),
    .X(_01571_));
 sg13g2_nand2b_1 _07437_ (.Y(_01572_),
    .B(\cordic_inst.cordic_state[32] ),
    .A_N(net1461));
 sg13g2_a21oi_1 _07438_ (.A1(\cordic_inst.cordic_state[33] ),
    .A2(net1462),
    .Y(_01573_),
    .B1(net1453));
 sg13g2_mux2_1 _07439_ (.A0(\cordic_inst.cordic_state[34] ),
    .A1(\cordic_inst.cordic_state[35] ),
    .S(net1462),
    .X(_01574_));
 sg13g2_a21oi_1 _07440_ (.A1(_01572_),
    .A2(_01573_),
    .Y(_01575_),
    .B1(net1345));
 sg13g2_o21ai_1 _07441_ (.B1(_01575_),
    .Y(_01576_),
    .A1(net1386),
    .A2(_01574_));
 sg13g2_mux2_1 _07442_ (.A0(\cordic_inst.cordic_state[36] ),
    .A1(net1426),
    .S(net1462),
    .X(_01577_));
 sg13g2_mux2_1 _07443_ (.A0(net1425),
    .A1(net1424),
    .S(net1462),
    .X(_01578_));
 sg13g2_mux2_1 _07444_ (.A0(_01577_),
    .A1(_01578_),
    .S(net1453),
    .X(_01579_));
 sg13g2_a22oi_1 _07445_ (.Y(_01580_),
    .B1(_01579_),
    .B2(_01141_),
    .A2(_01571_),
    .A1(net1439));
 sg13g2_a21o_1 _07446_ (.A2(_01580_),
    .A1(_01576_),
    .B1(net1432),
    .X(_01581_));
 sg13g2_and2_1 _07447_ (.A(net1410),
    .B(net1432),
    .X(_01582_));
 sg13g2_nand2_1 _07448_ (.Y(_01583_),
    .A(_00499_),
    .B(net1341));
 sg13g2_mux2_1 _07449_ (.A0(net1411),
    .A1(net1407),
    .S(net1456),
    .X(_01584_));
 sg13g2_mux4_1 _07450_ (.S0(net1454),
    .A0(net1413),
    .A1(net1412),
    .A2(net1411),
    .A3(net1408),
    .S1(net1448),
    .X(_01585_));
 sg13g2_mux4_1 _07451_ (.S0(net1457),
    .A0(net1415),
    .A1(\cordic_inst.cordic_state[49] ),
    .A2(net1414),
    .A3(\cordic_inst.cordic_state[51] ),
    .S1(net1449),
    .X(_01586_));
 sg13g2_mux2_1 _07452_ (.A0(_01585_),
    .A1(_01586_),
    .S(net1389),
    .X(_01587_));
 sg13g2_and2_1 _07453_ (.A(net1393),
    .B(_01587_),
    .X(_01588_));
 sg13g2_inv_1 _07454_ (.Y(_01589_),
    .A(_01588_));
 sg13g2_a22oi_1 _07455_ (.Y(_01590_),
    .B1(_01588_),
    .B2(net1432),
    .A2(net1341),
    .A1(_00499_));
 sg13g2_and2_1 _07456_ (.A(_01581_),
    .B(_01590_),
    .X(_01591_));
 sg13g2_nand2b_2 _07457_ (.Y(_01592_),
    .B(net764),
    .A_N(_01591_));
 sg13g2_nand2b_1 _07458_ (.Y(_01593_),
    .B(_01591_),
    .A_N(\cordic_inst.cordic_state[56] ));
 sg13g2_nand3_1 _07459_ (.B(_01592_),
    .C(_01593_),
    .A(net1349),
    .Y(_01594_));
 sg13g2_a22oi_1 _07460_ (.Y(_01595_),
    .B1(net1359),
    .B2(_01594_),
    .A2(net1476),
    .A1(_05559_));
 sg13g2_nand2_1 _07461_ (.Y(_01596_),
    .A(net1372),
    .B(_01595_));
 sg13g2_a21oi_1 _07462_ (.A1(net1559),
    .A2(net1367),
    .Y(_01597_),
    .B1(net1301));
 sg13g2_o21ai_1 _07463_ (.B1(net1780),
    .Y(_01598_),
    .A1(net764),
    .A2(net1290));
 sg13g2_a21oi_1 _07464_ (.A1(_01596_),
    .A2(_01597_),
    .Y(_00237_),
    .B1(_01598_));
 sg13g2_mux4_1 _07465_ (.S0(net1455),
    .A0(\cordic_inst.cordic_state[49] ),
    .A1(net1414),
    .A2(\cordic_inst.cordic_state[51] ),
    .A3(net1413),
    .S1(net1447),
    .X(_01599_));
 sg13g2_nor2_1 _07466_ (.A(net1442),
    .B(_01599_),
    .Y(_01600_));
 sg13g2_mux2_1 _07467_ (.A0(net1412),
    .A1(net1411),
    .S(net1456),
    .X(_01601_));
 sg13g2_a22oi_1 _07468_ (.Y(_01602_),
    .B1(_01601_),
    .B2(net1385),
    .A2(_01169_),
    .A1(net1407));
 sg13g2_a221oi_1 _07469_ (.B2(net1386),
    .C1(net1388),
    .B1(_01601_),
    .A1(net1407),
    .Y(_01603_),
    .A2(_01169_));
 sg13g2_or3_1 _07470_ (.A(net1436),
    .B(_01600_),
    .C(_01603_),
    .X(_01604_));
 sg13g2_mux4_1 _07471_ (.S0(net1454),
    .A0(net1418),
    .A1(net1417),
    .A2(net1416),
    .A3(net1415),
    .S1(net1447),
    .X(_01605_));
 sg13g2_mux4_1 _07472_ (.S0(net1454),
    .A0(net1422),
    .A1(net1421),
    .A2(net1420),
    .A3(net1419),
    .S1(net1447),
    .X(_01606_));
 sg13g2_mux2_1 _07473_ (.A0(_01605_),
    .A1(_01606_),
    .S(net1388),
    .X(_01607_));
 sg13g2_nand2b_1 _07474_ (.Y(_01608_),
    .B(\cordic_inst.cordic_state[33] ),
    .A_N(net1461));
 sg13g2_a21oi_1 _07475_ (.A1(\cordic_inst.cordic_state[34] ),
    .A2(net1462),
    .Y(_01609_),
    .B1(net1453));
 sg13g2_mux2_1 _07476_ (.A0(\cordic_inst.cordic_state[35] ),
    .A1(\cordic_inst.cordic_state[36] ),
    .S(net1462),
    .X(_01610_));
 sg13g2_or2_1 _07477_ (.X(_01611_),
    .B(_01610_),
    .A(net1386));
 sg13g2_a21oi_1 _07478_ (.A1(_01608_),
    .A2(_01609_),
    .Y(_01612_),
    .B1(net1345));
 sg13g2_mux2_1 _07479_ (.A0(net1426),
    .A1(net1425),
    .S(net1462),
    .X(_01613_));
 sg13g2_mux4_1 _07480_ (.S0(net1457),
    .A0(net1426),
    .A1(net1425),
    .A2(net1424),
    .A3(net1423),
    .S1(net1449),
    .X(_01614_));
 sg13g2_and2_1 _07481_ (.A(_01141_),
    .B(_01614_),
    .X(_01615_));
 sg13g2_a221oi_1 _07482_ (.B2(_01612_),
    .C1(_01615_),
    .B1(_01611_),
    .A1(net1440),
    .Y(_01616_),
    .A2(_01607_));
 sg13g2_mux2_1 _07483_ (.A0(_01604_),
    .A1(_01616_),
    .S(net1395),
    .X(_01617_));
 sg13g2_nand2_1 _07484_ (.Y(_01618_),
    .A(_01583_),
    .B(_01617_));
 sg13g2_a21oi_1 _07485_ (.A1(_01581_),
    .A2(_01590_),
    .Y(_01619_),
    .B1(net1238));
 sg13g2_xnor2_1 _07486_ (.Y(_01620_),
    .A(_01618_),
    .B(_01619_));
 sg13g2_or2_1 _07487_ (.X(_01621_),
    .B(_01620_),
    .A(_05581_));
 sg13g2_xnor2_1 _07488_ (.Y(_01622_),
    .A(_05581_),
    .B(_01620_));
 sg13g2_xnor2_1 _07489_ (.Y(_01623_),
    .A(_01592_),
    .B(_01622_));
 sg13g2_nand2b_1 _07490_ (.Y(_01624_),
    .B(net1475),
    .A_N(net1635));
 sg13g2_a21oi_1 _07491_ (.A1(net1280),
    .A2(_01623_),
    .Y(_01625_),
    .B1(net1369));
 sg13g2_a22oi_1 _07492_ (.Y(_01626_),
    .B1(_01624_),
    .B2(_01625_),
    .A2(net1364),
    .A1(net1550));
 sg13g2_a21oi_1 _07493_ (.A1(net722),
    .A2(net1300),
    .Y(_01627_),
    .B1(net1748));
 sg13g2_o21ai_1 _07494_ (.B1(_01627_),
    .Y(_00238_),
    .A1(net1301),
    .A2(_01626_));
 sg13g2_o21ai_1 _07495_ (.B1(_01621_),
    .Y(_01628_),
    .A1(_01592_),
    .A2(_01622_));
 sg13g2_mux4_1 _07496_ (.S0(net1455),
    .A0(net1417),
    .A1(net1416),
    .A2(net1415),
    .A3(\cordic_inst.cordic_state[49] ),
    .S1(net1448),
    .X(_01629_));
 sg13g2_mux4_1 _07497_ (.S0(net1454),
    .A0(net1421),
    .A1(net1420),
    .A2(net1419),
    .A3(net1418),
    .S1(net1447),
    .X(_01630_));
 sg13g2_mux2_1 _07498_ (.A0(_01629_),
    .A1(_01630_),
    .S(net1388),
    .X(_01631_));
 sg13g2_or2_1 _07499_ (.X(_01632_),
    .B(_01631_),
    .A(net1390));
 sg13g2_nand2_1 _07500_ (.Y(_01633_),
    .A(net1453),
    .B(_01577_));
 sg13g2_a21oi_1 _07501_ (.A1(net1386),
    .A2(_01574_),
    .Y(_01634_),
    .B1(net1345));
 sg13g2_mux4_1 _07502_ (.S0(net1457),
    .A0(net1425),
    .A1(net1424),
    .A2(net1423),
    .A3(net1422),
    .S1(net1449),
    .X(_01635_));
 sg13g2_o21ai_1 _07503_ (.B1(net1394),
    .Y(_01636_),
    .A1(net1342),
    .A2(_01635_));
 sg13g2_a21oi_1 _07504_ (.A1(_01633_),
    .A2(_01634_),
    .Y(_01637_),
    .B1(_01636_));
 sg13g2_nand2_2 _07505_ (.Y(_01638_),
    .A(net1386),
    .B(_01584_));
 sg13g2_mux4_1 _07506_ (.S0(net1455),
    .A0(net1414),
    .A1(\cordic_inst.cordic_state[51] ),
    .A2(net1413),
    .A3(net1412),
    .S1(net1447),
    .X(_01639_));
 sg13g2_nor2_1 _07507_ (.A(net1442),
    .B(_01639_),
    .Y(_01640_));
 sg13g2_a21oi_1 _07508_ (.A1(net1386),
    .A2(_01584_),
    .Y(_01641_),
    .B1(net1388));
 sg13g2_nor3_2 _07509_ (.A(net1436),
    .B(_01640_),
    .C(_01641_),
    .Y(_01642_));
 sg13g2_and2_1 _07510_ (.A(_01215_),
    .B(net1341),
    .X(_01643_));
 sg13g2_a221oi_1 _07511_ (.B2(net1429),
    .C1(_01643_),
    .B1(_01642_),
    .A1(_01632_),
    .Y(_01644_),
    .A2(_01637_));
 sg13g2_a21oi_1 _07512_ (.A1(_01591_),
    .A2(_01617_),
    .Y(_01645_),
    .B1(net1238));
 sg13g2_xnor2_1 _07513_ (.Y(_01646_),
    .A(_01644_),
    .B(_01645_));
 sg13g2_and2_1 _07514_ (.A(\cordic_inst.cordic_state[58] ),
    .B(_01646_),
    .X(_01647_));
 sg13g2_xor2_1 _07515_ (.B(_01646_),
    .A(\cordic_inst.cordic_state[58] ),
    .X(_01648_));
 sg13g2_and2_1 _07516_ (.A(_01628_),
    .B(_01648_),
    .X(_01649_));
 sg13g2_o21ai_1 _07517_ (.B1(net1349),
    .Y(_01650_),
    .A1(_01628_),
    .A2(_01648_));
 sg13g2_o21ai_1 _07518_ (.B1(net1359),
    .Y(_01651_),
    .A1(_01649_),
    .A2(_01650_));
 sg13g2_a21oi_1 _07519_ (.A1(_05558_),
    .A2(net1476),
    .Y(_01652_),
    .B1(net1366));
 sg13g2_a221oi_1 _07520_ (.B2(_01652_),
    .C1(net1303),
    .B1(_01651_),
    .A1(net1548),
    .Y(_01653_),
    .A2(net1366));
 sg13g2_o21ai_1 _07521_ (.B1(net1780),
    .Y(_01654_),
    .A1(net779),
    .A2(net1290));
 sg13g2_nor2_1 _07522_ (.A(_01653_),
    .B(_01654_),
    .Y(_00239_));
 sg13g2_a21oi_1 _07523_ (.A1(_01628_),
    .A2(_01648_),
    .Y(_01655_),
    .B1(_01647_));
 sg13g2_mux4_1 _07524_ (.S0(net1454),
    .A0(net1420),
    .A1(net1419),
    .A2(net1418),
    .A3(net1417),
    .S1(net1447),
    .X(_01656_));
 sg13g2_mux4_1 _07525_ (.S0(net1455),
    .A0(net1416),
    .A1(net1415),
    .A2(\cordic_inst.cordic_state[49] ),
    .A3(net1414),
    .S1(net1448),
    .X(_01657_));
 sg13g2_mux2_1 _07526_ (.A0(_01656_),
    .A1(_01657_),
    .S(net1442),
    .X(_01658_));
 sg13g2_nand2_1 _07527_ (.Y(_01659_),
    .A(net1449),
    .B(_01613_));
 sg13g2_a21oi_1 _07528_ (.A1(net1386),
    .A2(_01610_),
    .Y(_01660_),
    .B1(net1343));
 sg13g2_mux4_1 _07529_ (.S0(net1457),
    .A0(net1424),
    .A1(\cordic_inst.cordic_state[40] ),
    .A2(net1422),
    .A3(\cordic_inst.cordic_state[42] ),
    .S1(net1449),
    .X(_01661_));
 sg13g2_nor2_1 _07530_ (.A(net1342),
    .B(_01661_),
    .Y(_01662_));
 sg13g2_a21oi_1 _07531_ (.A1(_01659_),
    .A2(_01660_),
    .Y(_01663_),
    .B1(_01662_));
 sg13g2_o21ai_1 _07532_ (.B1(_01663_),
    .Y(_01664_),
    .A1(net1392),
    .A2(_01658_));
 sg13g2_nand3_1 _07533_ (.B(net1442),
    .C(_00506_),
    .A(net1407),
    .Y(_01665_));
 sg13g2_mux4_1 _07534_ (.S0(net1454),
    .A0(\cordic_inst.cordic_state[51] ),
    .A1(net1413),
    .A2(net1412),
    .A3(net1411),
    .S1(net1447),
    .X(_01666_));
 sg13g2_nand2_1 _07535_ (.Y(_01667_),
    .A(net1388),
    .B(_01666_));
 sg13g2_a21oi_2 _07536_ (.B1(net1436),
    .Y(_01668_),
    .A2(_01667_),
    .A1(_01665_));
 sg13g2_a22oi_1 _07537_ (.Y(_01669_),
    .B1(_01668_),
    .B2(net1429),
    .A2(net1341),
    .A1(_01215_));
 sg13g2_o21ai_1 _07538_ (.B1(_01669_),
    .Y(_01670_),
    .A1(net1429),
    .A2(_01664_));
 sg13g2_nand4_1 _07539_ (.B(_01590_),
    .C(_01617_),
    .A(_01581_),
    .Y(_01671_),
    .D(_01644_));
 sg13g2_nand2_1 _07540_ (.Y(_01672_),
    .A(net1244),
    .B(_01671_));
 sg13g2_xnor2_1 _07541_ (.Y(_01673_),
    .A(_01670_),
    .B(_01672_));
 sg13g2_nand2_1 _07542_ (.Y(_01674_),
    .A(\cordic_inst.cordic_state[59] ),
    .B(_01673_));
 sg13g2_xnor2_1 _07543_ (.Y(_01675_),
    .A(\cordic_inst.cordic_state[59] ),
    .B(_01673_));
 sg13g2_xnor2_1 _07544_ (.Y(_01676_),
    .A(_01655_),
    .B(_01675_));
 sg13g2_a22oi_1 _07545_ (.Y(_01677_),
    .B1(net1321),
    .B2(net1627),
    .A2(net1368),
    .A1(net1541));
 sg13g2_o21ai_1 _07546_ (.B1(_01677_),
    .Y(_01678_),
    .A1(_00464_),
    .A2(_01676_));
 sg13g2_a21oi_1 _07547_ (.A1(net1289),
    .A2(_01678_),
    .Y(_01679_),
    .B1(net1748));
 sg13g2_o21ai_1 _07548_ (.B1(_01679_),
    .Y(_00240_),
    .A1(_05580_),
    .A2(net1289));
 sg13g2_o21ai_1 _07549_ (.B1(_01674_),
    .Y(_01680_),
    .A1(_01655_),
    .A2(_01675_));
 sg13g2_mux2_1 _07550_ (.A0(_01570_),
    .A1(_01586_),
    .S(net1442),
    .X(_01681_));
 sg13g2_nor2_1 _07551_ (.A(net1392),
    .B(_01681_),
    .Y(_01682_));
 sg13g2_nor2_1 _07552_ (.A(net1344),
    .B(_01579_),
    .Y(_01683_));
 sg13g2_o21ai_1 _07553_ (.B1(net1394),
    .Y(_01684_),
    .A1(net1342),
    .A2(_01569_));
 sg13g2_nor3_1 _07554_ (.A(_01682_),
    .B(_01683_),
    .C(_01684_),
    .Y(_01685_));
 sg13g2_and2_1 _07555_ (.A(_00906_),
    .B(_01585_),
    .X(_01686_));
 sg13g2_inv_1 _07556_ (.Y(_01687_),
    .A(_01686_));
 sg13g2_a22oi_1 _07557_ (.Y(_01688_),
    .B1(_01686_),
    .B2(net1434),
    .A2(net1341),
    .A1(_01262_));
 sg13g2_inv_1 _07558_ (.Y(_01689_),
    .A(_01688_));
 sg13g2_nor2_1 _07559_ (.A(_01685_),
    .B(_01689_),
    .Y(_01690_));
 sg13g2_o21ai_1 _07560_ (.B1(net1244),
    .Y(_01691_),
    .A1(_01670_),
    .A2(_01671_));
 sg13g2_xor2_1 _07561_ (.B(_01691_),
    .A(_01690_),
    .X(_01692_));
 sg13g2_and2_1 _07562_ (.A(\cordic_inst.cordic_state[60] ),
    .B(_01692_),
    .X(_01693_));
 sg13g2_xor2_1 _07563_ (.B(_01692_),
    .A(\cordic_inst.cordic_state[60] ),
    .X(_01694_));
 sg13g2_a21oi_1 _07564_ (.A1(_01680_),
    .A2(_01694_),
    .Y(_01695_),
    .B1(_00479_));
 sg13g2_o21ai_1 _07565_ (.B1(_01695_),
    .Y(_01696_),
    .A1(_01680_),
    .A2(_01694_));
 sg13g2_a221oi_1 _07566_ (.B2(_01696_),
    .C1(net1368),
    .B1(_00462_),
    .A1(_05557_),
    .Y(_01697_),
    .A2(net1476));
 sg13g2_a221oi_1 _07567_ (.B2(_00479_),
    .C1(_01697_),
    .B1(_00463_),
    .A1(net1531),
    .Y(_01698_),
    .A2(net1368));
 sg13g2_o21ai_1 _07568_ (.B1(net1780),
    .Y(_01699_),
    .A1(net781),
    .A2(net1290));
 sg13g2_nor2_1 _07569_ (.A(_01698_),
    .B(_01699_),
    .Y(_00241_));
 sg13g2_a21oi_1 _07570_ (.A1(_01680_),
    .A2(_01694_),
    .Y(_01700_),
    .B1(_01693_));
 sg13g2_mux2_1 _07571_ (.A0(_01599_),
    .A1(_01605_),
    .S(net1389),
    .X(_01701_));
 sg13g2_nor2_1 _07572_ (.A(net1390),
    .B(_01701_),
    .Y(_01702_));
 sg13g2_nor2_1 _07573_ (.A(net1342),
    .B(_01606_),
    .Y(_01703_));
 sg13g2_o21ai_1 _07574_ (.B1(net1395),
    .Y(_01704_),
    .A1(net1344),
    .A2(_01614_));
 sg13g2_nor3_1 _07575_ (.A(_01702_),
    .B(_01703_),
    .C(_01704_),
    .Y(_01705_));
 sg13g2_nor2_1 _07576_ (.A(net1343),
    .B(_01602_),
    .Y(_01706_));
 sg13g2_a221oi_1 _07577_ (.B2(net1431),
    .C1(_01705_),
    .B1(_01706_),
    .A1(_01262_),
    .Y(_01707_),
    .A2(net1341));
 sg13g2_nor4_1 _07578_ (.A(_01670_),
    .B(_01671_),
    .C(_01685_),
    .D(_01689_),
    .Y(_01708_));
 sg13g2_nor2_1 _07579_ (.A(net1238),
    .B(_01708_),
    .Y(_01709_));
 sg13g2_xnor2_1 _07580_ (.Y(_01710_),
    .A(_01707_),
    .B(_01709_));
 sg13g2_nand2_1 _07581_ (.Y(_01711_),
    .A(\cordic_inst.cordic_state[61] ),
    .B(_01710_));
 sg13g2_xnor2_1 _07582_ (.Y(_01712_),
    .A(\cordic_inst.cordic_state[61] ),
    .B(_01710_));
 sg13g2_xnor2_1 _07583_ (.Y(_01713_),
    .A(_01700_),
    .B(_01712_));
 sg13g2_nand2b_1 _07584_ (.Y(_01714_),
    .B(net1475),
    .A_N(net1615));
 sg13g2_a21oi_1 _07585_ (.A1(net1280),
    .A2(_01713_),
    .Y(_01715_),
    .B1(net1365));
 sg13g2_a22oi_1 _07586_ (.Y(_01716_),
    .B1(_01714_),
    .B2(_01715_),
    .A2(net1365),
    .A1(net1526));
 sg13g2_a21oi_1 _07587_ (.A1(net749),
    .A2(net1303),
    .Y(_01717_),
    .B1(net1748));
 sg13g2_o21ai_1 _07588_ (.B1(_01717_),
    .Y(_00242_),
    .A1(net1303),
    .A2(_01716_));
 sg13g2_o21ai_1 _07589_ (.B1(_01711_),
    .Y(_01718_),
    .A1(_01700_),
    .A2(_01712_));
 sg13g2_mux2_1 _07590_ (.A0(_01629_),
    .A1(_01639_),
    .S(net1445),
    .X(_01719_));
 sg13g2_nor2_1 _07591_ (.A(net1390),
    .B(_01719_),
    .Y(_01720_));
 sg13g2_nor2_1 _07592_ (.A(_01142_),
    .B(_01630_),
    .Y(_01721_));
 sg13g2_o21ai_1 _07593_ (.B1(net1395),
    .Y(_01722_),
    .A1(net1344),
    .A2(_01635_));
 sg13g2_nor3_1 _07594_ (.A(_01720_),
    .B(_01721_),
    .C(_01722_),
    .Y(_01723_));
 sg13g2_nor2_1 _07595_ (.A(net1343),
    .B(_01638_),
    .Y(_01724_));
 sg13g2_a221oi_1 _07596_ (.B2(net1429),
    .C1(_01723_),
    .B1(_01724_),
    .A1(_01302_),
    .Y(_01725_),
    .A2(net1341));
 sg13g2_and2_1 _07597_ (.A(_01707_),
    .B(_01708_),
    .X(_01726_));
 sg13g2_nor2_1 _07598_ (.A(net1238),
    .B(_01726_),
    .Y(_01727_));
 sg13g2_xnor2_1 _07599_ (.Y(_01728_),
    .A(_01725_),
    .B(_01727_));
 sg13g2_and2_1 _07600_ (.A(\cordic_inst.cordic_state[62] ),
    .B(_01728_),
    .X(_01729_));
 sg13g2_xor2_1 _07601_ (.B(_01728_),
    .A(\cordic_inst.cordic_state[62] ),
    .X(_01730_));
 sg13g2_nand2_1 _07602_ (.Y(_01731_),
    .A(_01718_),
    .B(_01730_));
 sg13g2_nor2_1 _07603_ (.A(_01718_),
    .B(_01730_),
    .Y(_01732_));
 sg13g2_nand3b_1 _07604_ (.B(net1280),
    .C(_01731_),
    .Y(_01733_),
    .A_N(_01732_));
 sg13g2_a21oi_1 _07605_ (.A1(net1611),
    .A2(net1475),
    .Y(_01734_),
    .B1(net1365));
 sg13g2_nand2_1 _07606_ (.Y(_01735_),
    .A(_01733_),
    .B(_01734_));
 sg13g2_o21ai_1 _07607_ (.B1(_01735_),
    .Y(_01736_),
    .A1(net1525),
    .A2(net1372));
 sg13g2_nand2_1 _07608_ (.Y(_01737_),
    .A(net680),
    .B(net1299));
 sg13g2_a21oi_1 _07609_ (.A1(_01736_),
    .A2(_01737_),
    .Y(_00243_),
    .B1(net1747));
 sg13g2_mux2_1 _07610_ (.A0(_01657_),
    .A1(_01666_),
    .S(net1442),
    .X(_01738_));
 sg13g2_nand2b_1 _07611_ (.Y(_01739_),
    .B(net1436),
    .A_N(_01738_));
 sg13g2_nor2_1 _07612_ (.A(_01142_),
    .B(_01656_),
    .Y(_01740_));
 sg13g2_o21ai_1 _07613_ (.B1(net1395),
    .Y(_01741_),
    .A1(net1344),
    .A2(_01661_));
 sg13g2_nor2_1 _07614_ (.A(_01740_),
    .B(_01741_),
    .Y(_01742_));
 sg13g2_a21oi_2 _07615_ (.B1(net1341),
    .Y(_01743_),
    .A2(_01742_),
    .A1(_01739_));
 sg13g2_and2_1 _07616_ (.A(_01725_),
    .B(_01726_),
    .X(_01744_));
 sg13g2_nor2_1 _07617_ (.A(net1238),
    .B(_01744_),
    .Y(_01745_));
 sg13g2_xnor2_1 _07618_ (.Y(_01746_),
    .A(_01743_),
    .B(_01745_));
 sg13g2_nand2_1 _07619_ (.Y(_01747_),
    .A(\cordic_inst.cordic_state[63] ),
    .B(_01746_));
 sg13g2_xnor2_1 _07620_ (.Y(_01748_),
    .A(\cordic_inst.cordic_state[63] ),
    .B(_01746_));
 sg13g2_a21oi_1 _07621_ (.A1(_01718_),
    .A2(_01730_),
    .Y(_01749_),
    .B1(_01729_));
 sg13g2_xnor2_1 _07622_ (.Y(_01750_),
    .A(_01748_),
    .B(_01749_));
 sg13g2_a221oi_1 _07623_ (.B2(_01750_),
    .C1(net1364),
    .B1(net1281),
    .A1(_05556_),
    .Y(_01751_),
    .A2(net1475));
 sg13g2_a21oi_1 _07624_ (.A1(net1515),
    .A2(net1364),
    .Y(_01752_),
    .B1(_01751_));
 sg13g2_a21oi_1 _07625_ (.A1(net762),
    .A2(net1300),
    .Y(_01753_),
    .B1(net1748));
 sg13g2_o21ai_1 _07626_ (.B1(_01753_),
    .Y(_00244_),
    .A1(net1302),
    .A2(_01752_));
 sg13g2_o21ai_1 _07627_ (.B1(_01747_),
    .Y(_01754_),
    .A1(_01748_),
    .A2(_01749_));
 sg13g2_nor2_1 _07628_ (.A(net1440),
    .B(_01571_),
    .Y(_01755_));
 sg13g2_or2_1 _07629_ (.X(_01756_),
    .B(_01587_),
    .A(net1392));
 sg13g2_nor2_1 _07630_ (.A(net1431),
    .B(_01755_),
    .Y(_01757_));
 sg13g2_a21oi_1 _07631_ (.A1(_01756_),
    .A2(_01757_),
    .Y(_01758_),
    .B1(_01582_));
 sg13g2_nand2_1 _07632_ (.Y(_01759_),
    .A(_01743_),
    .B(_01744_));
 sg13g2_nand2_1 _07633_ (.Y(_01760_),
    .A(net1244),
    .B(_01759_));
 sg13g2_xor2_1 _07634_ (.B(_01760_),
    .A(_01758_),
    .X(_01761_));
 sg13g2_nand2_1 _07635_ (.Y(_01762_),
    .A(\cordic_inst.cordic_state[64] ),
    .B(_01761_));
 sg13g2_inv_1 _07636_ (.Y(_01763_),
    .A(_01762_));
 sg13g2_xor2_1 _07637_ (.B(_01761_),
    .A(\cordic_inst.cordic_state[64] ),
    .X(_01764_));
 sg13g2_and2_1 _07638_ (.A(_01754_),
    .B(_01764_),
    .X(_01765_));
 sg13g2_o21ai_1 _07639_ (.B1(net1349),
    .Y(_01766_),
    .A1(_01754_),
    .A2(_01764_));
 sg13g2_o21ai_1 _07640_ (.B1(net1359),
    .Y(_01767_),
    .A1(_01765_),
    .A2(_01766_));
 sg13g2_nand2b_1 _07641_ (.Y(_01768_),
    .B(net1474),
    .A_N(net1602));
 sg13g2_nand3_1 _07642_ (.B(_01767_),
    .C(_01768_),
    .A(net1372),
    .Y(_01769_));
 sg13g2_a21oi_1 _07643_ (.A1(net1733),
    .A2(net1363),
    .Y(_01770_),
    .B1(net1295));
 sg13g2_o21ai_1 _07644_ (.B1(net1755),
    .Y(_01771_),
    .A1(net769),
    .A2(net1286));
 sg13g2_a21oi_1 _07645_ (.A1(_01769_),
    .A2(_01770_),
    .Y(_00245_),
    .B1(_01771_));
 sg13g2_a21oi_2 _07646_ (.B1(_01763_),
    .Y(_01772_),
    .A2(_01764_),
    .A1(_01754_));
 sg13g2_nand2_1 _07647_ (.Y(_01773_),
    .A(net1407),
    .B(_01349_));
 sg13g2_o21ai_1 _07648_ (.B1(net1436),
    .Y(_01774_),
    .A1(_01600_),
    .A2(_01603_));
 sg13g2_o21ai_1 _07649_ (.B1(net1397),
    .Y(_01775_),
    .A1(net1437),
    .A2(_01607_));
 sg13g2_nand2b_1 _07650_ (.Y(_01776_),
    .B(_01774_),
    .A_N(_01775_));
 sg13g2_nand2_1 _07651_ (.Y(_01777_),
    .A(_01773_),
    .B(_01776_));
 sg13g2_a21o_2 _07652_ (.A2(_01757_),
    .A1(_01756_),
    .B1(_01759_),
    .X(_01778_));
 sg13g2_nand2_1 _07653_ (.Y(_01779_),
    .A(net1241),
    .B(_01778_));
 sg13g2_xor2_1 _07654_ (.B(_01779_),
    .A(_01777_),
    .X(_01780_));
 sg13g2_nand2b_1 _07655_ (.Y(_01781_),
    .B(\cordic_inst.cordic_state[65] ),
    .A_N(_01780_));
 sg13g2_xnor2_1 _07656_ (.Y(_01782_),
    .A(_05579_),
    .B(_01780_));
 sg13g2_xnor2_1 _07657_ (.Y(_01783_),
    .A(_01772_),
    .B(_01782_));
 sg13g2_a22oi_1 _07658_ (.Y(_01784_),
    .B1(net1322),
    .B2(net1597),
    .A2(net1360),
    .A1(net1727));
 sg13g2_o21ai_1 _07659_ (.B1(_01784_),
    .Y(_01785_),
    .A1(net1323),
    .A2(_01783_));
 sg13g2_a21oi_1 _07660_ (.A1(net1286),
    .A2(_01785_),
    .Y(_01786_),
    .B1(net1747));
 sg13g2_o21ai_1 _07661_ (.B1(_01786_),
    .Y(_00246_),
    .A1(_05579_),
    .A2(net1286));
 sg13g2_o21ai_1 _07662_ (.B1(_01781_),
    .Y(_01787_),
    .A1(_01772_),
    .A2(_01782_));
 sg13g2_o21ai_1 _07663_ (.B1(net1437),
    .Y(_01788_),
    .A1(_01640_),
    .A2(_01641_));
 sg13g2_nor2_1 _07664_ (.A(net1437),
    .B(_01631_),
    .Y(_01789_));
 sg13g2_nor2_1 _07665_ (.A(net1428),
    .B(_01789_),
    .Y(_01790_));
 sg13g2_a22oi_1 _07666_ (.Y(_01791_),
    .B1(_01788_),
    .B2(_01790_),
    .A2(_01349_),
    .A1(net1407));
 sg13g2_nor2b_1 _07667_ (.A(_01778_),
    .B_N(_01776_),
    .Y(_01792_));
 sg13g2_nor2_1 _07668_ (.A(net1236),
    .B(_01792_),
    .Y(_01793_));
 sg13g2_xnor2_1 _07669_ (.Y(_01794_),
    .A(_01791_),
    .B(_01793_));
 sg13g2_and2_1 _07670_ (.A(\cordic_inst.cordic_state[66] ),
    .B(_01794_),
    .X(_01795_));
 sg13g2_xor2_1 _07671_ (.B(_01794_),
    .A(\cordic_inst.cordic_state[66] ),
    .X(_01796_));
 sg13g2_o21ai_1 _07672_ (.B1(net1282),
    .Y(_01797_),
    .A1(_01787_),
    .A2(_01796_));
 sg13g2_a21o_1 _07673_ (.A2(_01796_),
    .A1(_01787_),
    .B1(_01797_),
    .X(_01798_));
 sg13g2_a21oi_1 _07674_ (.A1(net1590),
    .A2(net1474),
    .Y(_01799_),
    .B1(net1360));
 sg13g2_o21ai_1 _07675_ (.B1(net1285),
    .Y(_01800_),
    .A1(net1720),
    .A2(net1370));
 sg13g2_a21oi_1 _07676_ (.A1(_01798_),
    .A2(_01799_),
    .Y(_01801_),
    .B1(_01800_));
 sg13g2_a21oi_1 _07677_ (.A1(net739),
    .A2(net1294),
    .Y(_01802_),
    .B1(_01801_));
 sg13g2_nor2_1 _07678_ (.A(net1736),
    .B(net740),
    .Y(_00247_));
 sg13g2_a21oi_1 _07679_ (.A1(_01787_),
    .A2(_01796_),
    .Y(_01803_),
    .B1(_01795_));
 sg13g2_or2_1 _07680_ (.X(_01804_),
    .B(_01658_),
    .A(net1437));
 sg13g2_nand3_1 _07681_ (.B(_01665_),
    .C(_01667_),
    .A(net1437),
    .Y(_01805_));
 sg13g2_and3_1 _07682_ (.X(_01806_),
    .A(net1397),
    .B(_01804_),
    .C(_01805_));
 sg13g2_a21oi_1 _07683_ (.A1(net1407),
    .A2(_01382_),
    .Y(_01807_),
    .B1(_01806_));
 sg13g2_and2_1 _07684_ (.A(_01791_),
    .B(_01792_),
    .X(_01808_));
 sg13g2_nor2_1 _07685_ (.A(net1236),
    .B(_01808_),
    .Y(_01809_));
 sg13g2_xnor2_1 _07686_ (.Y(_01810_),
    .A(_01807_),
    .B(_01809_));
 sg13g2_nor2_1 _07687_ (.A(\cordic_inst.cordic_state[67] ),
    .B(_01810_),
    .Y(_01811_));
 sg13g2_xor2_1 _07688_ (.B(_01810_),
    .A(\cordic_inst.cordic_state[67] ),
    .X(_01812_));
 sg13g2_xnor2_1 _07689_ (.Y(_01813_),
    .A(_01803_),
    .B(_01812_));
 sg13g2_nor2_1 _07690_ (.A(_00485_),
    .B(_01813_),
    .Y(_01814_));
 sg13g2_a21oi_1 _07691_ (.A1(net1583),
    .A2(net1370),
    .Y(_01815_),
    .B1(_00461_));
 sg13g2_a21oi_1 _07692_ (.A1(net1714),
    .A2(net1360),
    .Y(_01816_),
    .B1(net1293));
 sg13g2_o21ai_1 _07693_ (.B1(_01816_),
    .Y(_01817_),
    .A1(_01814_),
    .A2(_01815_));
 sg13g2_o21ai_1 _07694_ (.B1(_01817_),
    .Y(_01818_),
    .A1(net820),
    .A2(net1285));
 sg13g2_nand2_1 _07695_ (.Y(_00248_),
    .A(net1754),
    .B(_01818_));
 sg13g2_nand2b_1 _07696_ (.Y(_01819_),
    .B(net1407),
    .A_N(_01397_));
 sg13g2_nor2_1 _07697_ (.A(net1390),
    .B(_01585_),
    .Y(_01820_));
 sg13g2_o21ai_1 _07698_ (.B1(_01348_),
    .Y(_01821_),
    .A1(net1436),
    .A2(_01681_));
 sg13g2_o21ai_1 _07699_ (.B1(_01819_),
    .Y(_01822_),
    .A1(_01820_),
    .A2(_01821_));
 sg13g2_a21oi_1 _07700_ (.A1(_01807_),
    .A2(_01808_),
    .Y(_01823_),
    .B1(net1236));
 sg13g2_xnor2_1 _07701_ (.Y(_01824_),
    .A(_01822_),
    .B(_01823_));
 sg13g2_nand2b_1 _07702_ (.Y(_01825_),
    .B(\cordic_inst.cordic_state[68] ),
    .A_N(_01824_));
 sg13g2_xor2_1 _07703_ (.B(_01824_),
    .A(\cordic_inst.cordic_state[68] ),
    .X(_01826_));
 sg13g2_a221oi_1 _07704_ (.B2(\cordic_inst.cordic_state[67] ),
    .C1(_01795_),
    .B1(_01810_),
    .A1(_01787_),
    .Y(_01827_),
    .A2(_01796_));
 sg13g2_or3_1 _07705_ (.A(_01811_),
    .B(_01826_),
    .C(_01827_),
    .X(_01828_));
 sg13g2_o21ai_1 _07706_ (.B1(_01826_),
    .Y(_01829_),
    .A1(_01811_),
    .A2(_01827_));
 sg13g2_nand3_1 _07707_ (.B(_01828_),
    .C(_01829_),
    .A(net1282),
    .Y(_01830_));
 sg13g2_a21oi_1 _07708_ (.A1(net1578),
    .A2(net1474),
    .Y(_01831_),
    .B1(net1360));
 sg13g2_nand2_1 _07709_ (.Y(_01832_),
    .A(_01830_),
    .B(_01831_));
 sg13g2_a21oi_1 _07710_ (.A1(_05567_),
    .A2(net1365),
    .Y(_01833_),
    .B1(net1299));
 sg13g2_a22oi_1 _07711_ (.Y(_01834_),
    .B1(_01832_),
    .B2(_01833_),
    .A2(net1295),
    .A1(net751));
 sg13g2_nor2_1 _07712_ (.A(net1736),
    .B(_01834_),
    .Y(_00249_));
 sg13g2_nand2_1 _07713_ (.Y(_01835_),
    .A(_01825_),
    .B(_01828_));
 sg13g2_nor3_1 _07714_ (.A(net1390),
    .B(net1443),
    .C(_01602_),
    .Y(_01836_));
 sg13g2_a21oi_1 _07715_ (.A1(net1390),
    .A2(_01701_),
    .Y(_01837_),
    .B1(_01836_));
 sg13g2_nor2_1 _07716_ (.A(net1427),
    .B(_01837_),
    .Y(_01838_));
 sg13g2_o21ai_1 _07717_ (.B1(_01819_),
    .Y(_01839_),
    .A1(net1427),
    .A2(_01837_));
 sg13g2_a21o_1 _07718_ (.A2(_01822_),
    .A1(net1241),
    .B1(_01823_),
    .X(_01840_));
 sg13g2_xnor2_1 _07719_ (.Y(_01841_),
    .A(_01839_),
    .B(_01840_));
 sg13g2_nor2b_1 _07720_ (.A(_01841_),
    .B_N(\cordic_inst.cordic_state[69] ),
    .Y(_01842_));
 sg13g2_inv_1 _07721_ (.Y(_01843_),
    .A(_01842_));
 sg13g2_nand2b_1 _07722_ (.Y(_01844_),
    .B(_01841_),
    .A_N(\cordic_inst.cordic_state[69] ));
 sg13g2_nand2_1 _07723_ (.Y(_01845_),
    .A(_01843_),
    .B(_01844_));
 sg13g2_xor2_1 _07724_ (.B(_01845_),
    .A(_01835_),
    .X(_01846_));
 sg13g2_a221oi_1 _07725_ (.B2(net1573),
    .C1(net1293),
    .B1(net1322),
    .A1(net1703),
    .Y(_01847_),
    .A2(net1360));
 sg13g2_o21ai_1 _07726_ (.B1(_01847_),
    .Y(_01848_),
    .A1(net1323),
    .A2(_01846_));
 sg13g2_o21ai_1 _07727_ (.B1(_01848_),
    .Y(_01849_),
    .A1(net791),
    .A2(net1285));
 sg13g2_nand2_1 _07728_ (.Y(_00250_),
    .A(net1754),
    .B(_01849_));
 sg13g2_nand2_1 _07729_ (.Y(_01850_),
    .A(net1408),
    .B(_01428_));
 sg13g2_nor2_1 _07730_ (.A(net1435),
    .B(_01719_),
    .Y(_01851_));
 sg13g2_nand2_1 _07731_ (.Y(_01852_),
    .A(net1435),
    .B(_01638_));
 sg13g2_nand2_1 _07732_ (.Y(_01853_),
    .A(_01348_),
    .B(_01852_));
 sg13g2_o21ai_1 _07733_ (.B1(_01850_),
    .Y(_01854_),
    .A1(_01851_),
    .A2(_01853_));
 sg13g2_a21o_1 _07734_ (.A2(_01838_),
    .A1(net1241),
    .B1(_01840_),
    .X(_01855_));
 sg13g2_xor2_1 _07735_ (.B(_01855_),
    .A(_01854_),
    .X(_01856_));
 sg13g2_and2_1 _07736_ (.A(\cordic_inst.cordic_state[70] ),
    .B(_01856_),
    .X(_01857_));
 sg13g2_inv_1 _07737_ (.Y(_01858_),
    .A(_01857_));
 sg13g2_xnor2_1 _07738_ (.Y(_01859_),
    .A(\cordic_inst.cordic_state[70] ),
    .B(_01856_));
 sg13g2_nand3_1 _07739_ (.B(_01828_),
    .C(_01843_),
    .A(_01825_),
    .Y(_01860_));
 sg13g2_nand2_1 _07740_ (.Y(_01861_),
    .A(_01844_),
    .B(_01860_));
 sg13g2_nand3b_1 _07741_ (.B(_01860_),
    .C(_01844_),
    .Y(_01862_),
    .A_N(_01859_));
 sg13g2_a21oi_1 _07742_ (.A1(_01859_),
    .A2(_01861_),
    .Y(_01863_),
    .B1(_00485_));
 sg13g2_a21oi_1 _07743_ (.A1(_05555_),
    .A2(_00459_),
    .Y(_01864_),
    .B1(_00461_));
 sg13g2_a21o_1 _07744_ (.A2(_01863_),
    .A1(_01862_),
    .B1(_01864_),
    .X(_01865_));
 sg13g2_o21ai_1 _07745_ (.B1(_01865_),
    .Y(_01866_),
    .A1(net1698),
    .A2(net1370));
 sg13g2_o21ai_1 _07746_ (.B1(net1756),
    .Y(_01867_),
    .A1(net752),
    .A2(net1286));
 sg13g2_a21oi_1 _07747_ (.A1(net1286),
    .A2(_01866_),
    .Y(_00251_),
    .B1(_01867_));
 sg13g2_a22oi_1 _07748_ (.Y(_01868_),
    .B1(_01738_),
    .B2(net1390),
    .A2(_01447_),
    .A1(net1408));
 sg13g2_o21ai_1 _07749_ (.B1(_01850_),
    .Y(_01869_),
    .A1(net1427),
    .A2(_01868_));
 sg13g2_a21o_1 _07750_ (.A2(_01854_),
    .A1(net1241),
    .B1(_01855_),
    .X(_01870_));
 sg13g2_xor2_1 _07751_ (.B(_01870_),
    .A(_01869_),
    .X(_01871_));
 sg13g2_nand2_1 _07752_ (.Y(_01872_),
    .A(\cordic_inst.cordic_state[71] ),
    .B(_01871_));
 sg13g2_inv_1 _07753_ (.Y(_01873_),
    .A(_01872_));
 sg13g2_xor2_1 _07754_ (.B(_01871_),
    .A(\cordic_inst.cordic_state[71] ),
    .X(_01874_));
 sg13g2_inv_1 _07755_ (.Y(_01875_),
    .A(_01874_));
 sg13g2_nand3_1 _07756_ (.B(_01862_),
    .C(_01875_),
    .A(_01858_),
    .Y(_01876_));
 sg13g2_a21oi_1 _07757_ (.A1(_01858_),
    .A2(_01862_),
    .Y(_01877_),
    .B1(_01875_));
 sg13g2_nand3b_1 _07758_ (.B(_00463_),
    .C(_01876_),
    .Y(_01878_),
    .A_N(_01877_));
 sg13g2_a22oi_1 _07759_ (.Y(_01879_),
    .B1(net1322),
    .B2(net1565),
    .A2(net1360),
    .A1(net1693));
 sg13g2_a21oi_1 _07760_ (.A1(_01878_),
    .A2(_01879_),
    .Y(_01880_),
    .B1(net1295));
 sg13g2_a21oi_1 _07761_ (.A1(net760),
    .A2(net1295),
    .Y(_01881_),
    .B1(_01880_));
 sg13g2_nand2_1 _07762_ (.Y(_00252_),
    .A(net1756),
    .B(_01881_));
 sg13g2_or2_1 _07763_ (.X(_01882_),
    .B(_01877_),
    .A(_01873_));
 sg13g2_o21ai_1 _07764_ (.B1(net1410),
    .Y(_01883_),
    .A1(net1432),
    .A2(_00499_));
 sg13g2_o21ai_1 _07765_ (.B1(_01883_),
    .Y(_01884_),
    .A1(net1433),
    .A2(_01589_));
 sg13g2_a21o_2 _07766_ (.A2(_01869_),
    .A1(net1242),
    .B1(_01870_),
    .X(_01885_));
 sg13g2_xor2_1 _07767_ (.B(_01885_),
    .A(_01884_),
    .X(_01886_));
 sg13g2_nand2_1 _07768_ (.Y(_01887_),
    .A(\cordic_inst.cordic_state[72] ),
    .B(_01886_));
 sg13g2_xor2_1 _07769_ (.B(_01886_),
    .A(\cordic_inst.cordic_state[72] ),
    .X(_01888_));
 sg13g2_and2_1 _07770_ (.A(_01882_),
    .B(_01888_),
    .X(_01889_));
 sg13g2_o21ai_1 _07771_ (.B1(_01888_),
    .Y(_01890_),
    .A1(_01873_),
    .A2(_01877_));
 sg13g2_o21ai_1 _07772_ (.B1(net1280),
    .Y(_01891_),
    .A1(_01882_),
    .A2(_01888_));
 sg13g2_a21oi_1 _07773_ (.A1(net1513),
    .A2(net1475),
    .Y(_01892_),
    .B1(net1363));
 sg13g2_o21ai_1 _07774_ (.B1(_01892_),
    .Y(_01893_),
    .A1(_01889_),
    .A2(_01891_));
 sg13g2_a21oi_1 _07775_ (.A1(_05564_),
    .A2(net1364),
    .Y(_01894_),
    .B1(net1298));
 sg13g2_a22oi_1 _07776_ (.Y(_01895_),
    .B1(_01893_),
    .B2(_01894_),
    .A2(net1298),
    .A1(net741));
 sg13g2_nor2_1 _07777_ (.A(net1743),
    .B(_01895_),
    .Y(_00253_));
 sg13g2_o21ai_1 _07778_ (.B1(_01883_),
    .Y(_01896_),
    .A1(net1433),
    .A2(_01604_));
 sg13g2_a21o_1 _07779_ (.A2(_01884_),
    .A1(net1244),
    .B1(_01885_),
    .X(_01897_));
 sg13g2_or2_1 _07780_ (.X(_01898_),
    .B(_01897_),
    .A(_01896_));
 sg13g2_nand2_1 _07781_ (.Y(_01899_),
    .A(_01896_),
    .B(_01897_));
 sg13g2_nand3_1 _07782_ (.B(_01898_),
    .C(_01899_),
    .A(net777),
    .Y(_01900_));
 sg13g2_inv_1 _07783_ (.Y(_01901_),
    .A(_01900_));
 sg13g2_nand2_1 _07784_ (.Y(_01902_),
    .A(_01887_),
    .B(_01890_));
 sg13g2_a21oi_1 _07785_ (.A1(_01898_),
    .A2(_01899_),
    .Y(_01903_),
    .B1(\cordic_inst.cordic_state[73] ));
 sg13g2_a21oi_1 _07786_ (.A1(_01887_),
    .A2(_01890_),
    .Y(_01904_),
    .B1(_01903_));
 sg13g2_nor2_1 _07787_ (.A(_01901_),
    .B(_01903_),
    .Y(_01905_));
 sg13g2_o21ai_1 _07788_ (.B1(_00463_),
    .Y(_01906_),
    .A1(_01902_),
    .A2(_01905_));
 sg13g2_a21oi_1 _07789_ (.A1(_01900_),
    .A2(_01904_),
    .Y(_01907_),
    .B1(_01906_));
 sg13g2_a221oi_1 _07790_ (.B2(net1507),
    .C1(_01907_),
    .B1(net1321),
    .A1(net1679),
    .Y(_01908_),
    .A2(net1364));
 sg13g2_a21oi_1 _07791_ (.A1(net777),
    .A2(net1298),
    .Y(_01909_),
    .B1(net1743));
 sg13g2_o21ai_1 _07792_ (.B1(_01909_),
    .Y(_00254_),
    .A1(net1298),
    .A2(_01908_));
 sg13g2_nor2b_2 _07793_ (.A(_01484_),
    .B_N(net1409),
    .Y(_01910_));
 sg13g2_a21oi_2 _07794_ (.B1(_01910_),
    .Y(_01911_),
    .A2(_01642_),
    .A1(net1394));
 sg13g2_nand2_1 _07795_ (.Y(_01912_),
    .A(net1244),
    .B(_01898_));
 sg13g2_xor2_1 _07796_ (.B(_01912_),
    .A(_01911_),
    .X(_01913_));
 sg13g2_nand2_1 _07797_ (.Y(_01914_),
    .A(\cordic_inst.cordic_state[74] ),
    .B(_01913_));
 sg13g2_xor2_1 _07798_ (.B(_01913_),
    .A(\cordic_inst.cordic_state[74] ),
    .X(_01915_));
 sg13g2_o21ai_1 _07799_ (.B1(_01915_),
    .Y(_01916_),
    .A1(_01901_),
    .A2(_01904_));
 sg13g2_or3_1 _07800_ (.A(_01901_),
    .B(_01904_),
    .C(_01915_),
    .X(_01917_));
 sg13g2_nand3_1 _07801_ (.B(_01916_),
    .C(_01917_),
    .A(net1280),
    .Y(_01918_));
 sg13g2_a21oi_1 _07802_ (.A1(net1506),
    .A2(net1475),
    .Y(_01919_),
    .B1(net1365));
 sg13g2_o21ai_1 _07803_ (.B1(net1291),
    .Y(_01920_),
    .A1(net1674),
    .A2(net1372));
 sg13g2_a21oi_1 _07804_ (.A1(_01918_),
    .A2(_01919_),
    .Y(_01921_),
    .B1(_01920_));
 sg13g2_a21oi_1 _07805_ (.A1(net729),
    .A2(net1299),
    .Y(_01922_),
    .B1(_01921_));
 sg13g2_nor2_1 _07806_ (.A(net1743),
    .B(net730),
    .Y(_00255_));
 sg13g2_nor2_1 _07807_ (.A(net784),
    .B(net1291),
    .Y(_01923_));
 sg13g2_a21oi_2 _07808_ (.B1(_01910_),
    .Y(_01924_),
    .A2(_01668_),
    .A1(net1394));
 sg13g2_o21ai_1 _07809_ (.B1(_01912_),
    .Y(_01925_),
    .A1(net1239),
    .A2(_01911_));
 sg13g2_xnor2_1 _07810_ (.Y(_01926_),
    .A(_01924_),
    .B(_01925_));
 sg13g2_inv_1 _07811_ (.Y(_01927_),
    .A(_01926_));
 sg13g2_nand2_1 _07812_ (.Y(_01928_),
    .A(_05578_),
    .B(_01927_));
 sg13g2_nand2_1 _07813_ (.Y(_01929_),
    .A(\cordic_inst.cordic_state[75] ),
    .B(_01926_));
 sg13g2_and2_1 _07814_ (.A(_01914_),
    .B(_01929_),
    .X(_01930_));
 sg13g2_nand2_1 _07815_ (.Y(_01931_),
    .A(_01916_),
    .B(_01930_));
 sg13g2_nand3_1 _07816_ (.B(_01928_),
    .C(_01930_),
    .A(_01916_),
    .Y(_01932_));
 sg13g2_a22oi_1 _07817_ (.Y(_01933_),
    .B1(_01928_),
    .B2(_01929_),
    .A2(_01916_),
    .A1(_01914_));
 sg13g2_nor2_1 _07818_ (.A(_00479_),
    .B(_01933_),
    .Y(_01934_));
 sg13g2_a21oi_1 _07819_ (.A1(_01932_),
    .A2(_01934_),
    .Y(_01935_),
    .B1(net1324));
 sg13g2_a221oi_1 _07820_ (.B2(net1502),
    .C1(_01935_),
    .B1(net1321),
    .A1(net1670),
    .Y(_01936_),
    .A2(net1365));
 sg13g2_o21ai_1 _07821_ (.B1(net1756),
    .Y(_00256_),
    .A1(_01923_),
    .A2(_01936_));
 sg13g2_o21ai_1 _07822_ (.B1(net1410),
    .Y(_01937_),
    .A1(net1433),
    .A2(_01262_));
 sg13g2_o21ai_1 _07823_ (.B1(_01937_),
    .Y(_01938_),
    .A1(net1433),
    .A2(_01687_));
 sg13g2_nor2_1 _07824_ (.A(net1239),
    .B(_01924_),
    .Y(_01939_));
 sg13g2_or2_1 _07825_ (.X(_01940_),
    .B(_01939_),
    .A(_01925_));
 sg13g2_xor2_1 _07826_ (.B(_01940_),
    .A(_01938_),
    .X(_01941_));
 sg13g2_nand2_1 _07827_ (.Y(_01942_),
    .A(net1406),
    .B(_01941_));
 sg13g2_xnor2_1 _07828_ (.Y(_01943_),
    .A(\cordic_inst.cordic_state[76] ),
    .B(_01941_));
 sg13g2_nand2_1 _07829_ (.Y(_01944_),
    .A(_01928_),
    .B(_01931_));
 sg13g2_a221oi_1 _07830_ (.B2(_01916_),
    .C1(_01943_),
    .B1(_01930_),
    .A1(_05578_),
    .Y(_01945_),
    .A2(_01927_));
 sg13g2_a21o_1 _07831_ (.A2(_01944_),
    .A1(_01943_),
    .B1(_00485_),
    .X(_01946_));
 sg13g2_a21oi_1 _07832_ (.A1(net1497),
    .A2(net1478),
    .Y(_01947_),
    .B1(net1364));
 sg13g2_o21ai_1 _07833_ (.B1(_01947_),
    .Y(_01948_),
    .A1(_01945_),
    .A2(_01946_));
 sg13g2_o21ai_1 _07834_ (.B1(_01948_),
    .Y(_01949_),
    .A1(net1666),
    .A2(net1372));
 sg13g2_nand2_1 _07835_ (.Y(_01950_),
    .A(net1406),
    .B(net1304));
 sg13g2_a21oi_1 _07836_ (.A1(_01949_),
    .A2(_01950_),
    .Y(_00257_),
    .B1(net1749));
 sg13g2_a22oi_1 _07837_ (.Y(_01951_),
    .B1(net1321),
    .B2(net1496),
    .A2(net1364),
    .A1(net1662));
 sg13g2_a21oi_1 _07838_ (.A1(net1406),
    .A2(_01941_),
    .Y(_01952_),
    .B1(_01945_));
 sg13g2_o21ai_1 _07839_ (.B1(net1245),
    .Y(_01953_),
    .A1(_01938_),
    .A2(_01940_));
 sg13g2_nand2_1 _07840_ (.Y(_01954_),
    .A(net1395),
    .B(_01706_));
 sg13g2_and2_1 _07841_ (.A(_01937_),
    .B(_01954_),
    .X(_01955_));
 sg13g2_xnor2_1 _07842_ (.Y(_01956_),
    .A(_01953_),
    .B(_01955_));
 sg13g2_and2_1 _07843_ (.A(_05577_),
    .B(_01956_),
    .X(_01957_));
 sg13g2_xnor2_1 _07844_ (.Y(_01958_),
    .A(_05577_),
    .B(_01956_));
 sg13g2_a21oi_1 _07845_ (.A1(_01952_),
    .A2(_01958_),
    .Y(_01959_),
    .B1(net1324));
 sg13g2_o21ai_1 _07846_ (.B1(_01959_),
    .Y(_01960_),
    .A1(_01952_),
    .A2(_01958_));
 sg13g2_o21ai_1 _07847_ (.B1(_01942_),
    .Y(_01961_),
    .A1(_05577_),
    .A2(_01956_));
 sg13g2_nor2_1 _07848_ (.A(_01945_),
    .B(_01961_),
    .Y(_01962_));
 sg13g2_a21oi_1 _07849_ (.A1(_01951_),
    .A2(_01960_),
    .Y(_01963_),
    .B1(net1298));
 sg13g2_a21oi_1 _07850_ (.A1(net744),
    .A2(net1304),
    .Y(_01964_),
    .B1(_01963_));
 sg13g2_nand2_1 _07851_ (.Y(_00258_),
    .A(net1763),
    .B(net745));
 sg13g2_nor3_1 _07852_ (.A(net1429),
    .B(net1343),
    .C(_01638_),
    .Y(_01965_));
 sg13g2_o21ai_1 _07853_ (.B1(net1409),
    .Y(_01966_),
    .A1(net1429),
    .A2(_01302_));
 sg13g2_nand2b_2 _07854_ (.Y(_01967_),
    .B(_01966_),
    .A_N(_01965_));
 sg13g2_o21ai_1 _07855_ (.B1(_01953_),
    .Y(_01968_),
    .A1(net1239),
    .A2(_01955_));
 sg13g2_xor2_1 _07856_ (.B(_01968_),
    .A(_01967_),
    .X(_01969_));
 sg13g2_xnor2_1 _07857_ (.Y(_01970_),
    .A(\cordic_inst.cordic_state[78] ),
    .B(_01969_));
 sg13g2_inv_1 _07858_ (.Y(_01971_),
    .A(_01970_));
 sg13g2_nor2_1 _07859_ (.A(_01957_),
    .B(_01962_),
    .Y(_01972_));
 sg13g2_nor3_1 _07860_ (.A(_01957_),
    .B(_01962_),
    .C(_01970_),
    .Y(_01973_));
 sg13g2_o21ai_1 _07861_ (.B1(net1281),
    .Y(_01974_),
    .A1(_01971_),
    .A2(_01972_));
 sg13g2_a21oi_1 _07862_ (.A1(net1492),
    .A2(net1475),
    .Y(_01975_),
    .B1(net1364));
 sg13g2_o21ai_1 _07863_ (.B1(_01975_),
    .Y(_01976_),
    .A1(_01973_),
    .A2(_01974_));
 sg13g2_o21ai_1 _07864_ (.B1(_01976_),
    .Y(_01977_),
    .A1(net1658),
    .A2(net1372));
 sg13g2_o21ai_1 _07865_ (.B1(net1763),
    .Y(_01978_),
    .A1(net782),
    .A2(net1291));
 sg13g2_a21oi_1 _07866_ (.A1(net1291),
    .A2(_01977_),
    .Y(_00259_),
    .B1(_01978_));
 sg13g2_a21oi_1 _07867_ (.A1(\cordic_inst.cordic_state[78] ),
    .A2(_01969_),
    .Y(_01979_),
    .B1(_01973_));
 sg13g2_a21oi_1 _07868_ (.A1(net1245),
    .A2(_01967_),
    .Y(_01980_),
    .B1(_01968_));
 sg13g2_xnor2_1 _07869_ (.Y(_01981_),
    .A(_01561_),
    .B(_01980_));
 sg13g2_o21ai_1 _07870_ (.B1(net1349),
    .Y(_01982_),
    .A1(_01979_),
    .A2(_01981_));
 sg13g2_a21oi_1 _07871_ (.A1(_01979_),
    .A2(_01981_),
    .Y(_01983_),
    .B1(_01982_));
 sg13g2_nor2_1 _07872_ (.A(_00464_),
    .B(_01983_),
    .Y(_01984_));
 sg13g2_a221oi_1 _07873_ (.B2(net1486),
    .C1(_01984_),
    .B1(net1321),
    .A1(net1656),
    .Y(_01985_),
    .A2(net1365));
 sg13g2_a21oi_1 _07874_ (.A1(net1405),
    .A2(net1300),
    .Y(_01986_),
    .B1(net1749));
 sg13g2_o21ai_1 _07875_ (.B1(_01986_),
    .Y(_00260_),
    .A1(net1300),
    .A2(_01985_));
 sg13g2_nor3_1 _07876_ (.A(\cordic_inst.result_ready ),
    .B(_05575_),
    .C(cordic_busy),
    .Y(_01987_));
 sg13g2_nand2b_1 _07877_ (.Y(_01988_),
    .B(net483),
    .A_N(net500));
 sg13g2_a21oi_1 _07878_ (.A1(_00463_),
    .A2(_01988_),
    .Y(_00261_),
    .B1(net1747));
 sg13g2_o21ai_1 _07879_ (.B1(\cordic_inst.operation_started ),
    .Y(_01989_),
    .A1(\cordic_inst.result_ready ),
    .A2(cordic_busy));
 sg13g2_nand2_1 _07880_ (.Y(_01990_),
    .A(net483),
    .B(cordic_busy));
 sg13g2_a21oi_1 _07881_ (.A1(_01989_),
    .A2(net484),
    .Y(_00262_),
    .B1(_00466_));
 sg13g2_nor2b_1 _07882_ (.A(net633),
    .B_N(\cordic_inst.result_ready ),
    .Y(_01991_));
 sg13g2_nor3_1 _07883_ (.A(cordic_en_get_normalize),
    .B(cordic_en_get_atan2),
    .C(cordic_en_get_sin_cos),
    .Y(_01992_));
 sg13g2_a21oi_1 _07884_ (.A1(net634),
    .A2(_01992_),
    .Y(_01993_),
    .B1(net500));
 sg13g2_nor2_1 _07885_ (.A(_00466_),
    .B(net635),
    .Y(_00263_));
 sg13g2_a22oi_1 _07886_ (.Y(_01994_),
    .B1(net1357),
    .B2(net418),
    .A2(net1380),
    .A1(net1559));
 sg13g2_inv_1 _07887_ (.Y(_00264_),
    .A(_01994_));
 sg13g2_a22oi_1 _07888_ (.Y(_01995_),
    .B1(net1356),
    .B2(net472),
    .A2(net1379),
    .A1(net1554));
 sg13g2_inv_1 _07889_ (.Y(_00265_),
    .A(net473));
 sg13g2_a22oi_1 _07890_ (.Y(_01996_),
    .B1(net1357),
    .B2(net397),
    .A2(net1376),
    .A1(net1548));
 sg13g2_inv_1 _07891_ (.Y(_00266_),
    .A(net398));
 sg13g2_a22oi_1 _07892_ (.Y(_01997_),
    .B1(net1353),
    .B2(net466),
    .A2(net1376),
    .A1(net1541));
 sg13g2_inv_1 _07893_ (.Y(_00267_),
    .A(_01997_));
 sg13g2_a22oi_1 _07894_ (.Y(_01998_),
    .B1(net1356),
    .B2(net434),
    .A2(net1379),
    .A1(net1531));
 sg13g2_inv_1 _07895_ (.Y(_00268_),
    .A(net435));
 sg13g2_a22oi_1 _07896_ (.Y(_01999_),
    .B1(net1352),
    .B2(net438),
    .A2(net1375),
    .A1(net1526));
 sg13g2_inv_1 _07897_ (.Y(_00269_),
    .A(net439));
 sg13g2_a22oi_1 _07898_ (.Y(_02000_),
    .B1(net1358),
    .B2(net492),
    .A2(net1375),
    .A1(net1525));
 sg13g2_inv_1 _07899_ (.Y(_00270_),
    .A(net493));
 sg13g2_a22oi_1 _07900_ (.Y(_02001_),
    .B1(net1353),
    .B2(net578),
    .A2(net1376),
    .A1(net1518));
 sg13g2_inv_1 _07901_ (.Y(_00271_),
    .A(net579));
 sg13g2_a22oi_1 _07902_ (.Y(_02002_),
    .B1(net1351),
    .B2(net453),
    .A2(net1374),
    .A1(net1733));
 sg13g2_inv_1 _07903_ (.Y(_00272_),
    .A(net454));
 sg13g2_a22oi_1 _07904_ (.Y(_02003_),
    .B1(net1353),
    .B2(net383),
    .A2(net1376),
    .A1(net1727));
 sg13g2_inv_1 _07905_ (.Y(_00273_),
    .A(_02003_));
 sg13g2_a22oi_1 _07906_ (.Y(_02004_),
    .B1(net1353),
    .B2(net459),
    .A2(net1376),
    .A1(net1720));
 sg13g2_inv_1 _07907_ (.Y(_00274_),
    .A(net460));
 sg13g2_a22oi_1 _07908_ (.Y(_02005_),
    .B1(net1350),
    .B2(net446),
    .A2(net1373),
    .A1(net1714));
 sg13g2_inv_1 _07909_ (.Y(_00275_),
    .A(net447));
 sg13g2_a22oi_1 _07910_ (.Y(_02006_),
    .B1(net1352),
    .B2(net416),
    .A2(net1375),
    .A1(net1709));
 sg13g2_inv_1 _07911_ (.Y(_00276_),
    .A(net417));
 sg13g2_a22oi_1 _07912_ (.Y(_02007_),
    .B1(net1356),
    .B2(net425),
    .A2(net1379),
    .A1(net1703));
 sg13g2_inv_1 _07913_ (.Y(_00277_),
    .A(net426));
 sg13g2_a22oi_1 _07914_ (.Y(_02008_),
    .B1(net1356),
    .B2(net358),
    .A2(net1379),
    .A1(net1698));
 sg13g2_inv_1 _07915_ (.Y(_00278_),
    .A(net359));
 sg13g2_a22oi_1 _07916_ (.Y(_02009_),
    .B1(net1356),
    .B2(net363),
    .A2(net1379),
    .A1(net1693));
 sg13g2_inv_1 _07917_ (.Y(_00279_),
    .A(_02009_));
 sg13g2_a22oi_1 _07918_ (.Y(_02010_),
    .B1(net1356),
    .B2(net429),
    .A2(net1379),
    .A1(net1685));
 sg13g2_inv_1 _07919_ (.Y(_00280_),
    .A(net430));
 sg13g2_a22oi_1 _07920_ (.Y(_02011_),
    .B1(net1355),
    .B2(net520),
    .A2(net1377),
    .A1(net1679));
 sg13g2_inv_1 _07921_ (.Y(_00281_),
    .A(net521));
 sg13g2_a22oi_1 _07922_ (.Y(_02012_),
    .B1(net1354),
    .B2(net399),
    .A2(net1378),
    .A1(net1674));
 sg13g2_inv_1 _07923_ (.Y(_00282_),
    .A(net400));
 sg13g2_a22oi_1 _07924_ (.Y(_02013_),
    .B1(net1352),
    .B2(net541),
    .A2(net1375),
    .A1(net1670));
 sg13g2_inv_1 _07925_ (.Y(_00283_),
    .A(net542));
 sg13g2_a22oi_1 _07926_ (.Y(_02014_),
    .B1(net1355),
    .B2(net442),
    .A2(net1378),
    .A1(net1666));
 sg13g2_inv_1 _07927_ (.Y(_00284_),
    .A(net443));
 sg13g2_a22oi_1 _07928_ (.Y(_02015_),
    .B1(net1354),
    .B2(net474),
    .A2(net1377),
    .A1(net1662));
 sg13g2_inv_1 _07929_ (.Y(_00285_),
    .A(_02015_));
 sg13g2_a22oi_1 _07930_ (.Y(_02016_),
    .B1(net1354),
    .B2(net507),
    .A2(net1377),
    .A1(net1658));
 sg13g2_inv_1 _07931_ (.Y(_00286_),
    .A(net508));
 sg13g2_a22oi_1 _07932_ (.Y(_02017_),
    .B1(net1354),
    .B2(net379),
    .A2(net1377),
    .A1(net1655));
 sg13g2_inv_1 _07933_ (.Y(_00287_),
    .A(_02017_));
 sg13g2_a22oi_1 _07934_ (.Y(_02018_),
    .B1(net1353),
    .B2(net444),
    .A2(net1376),
    .A1(net1654));
 sg13g2_inv_1 _07935_ (.Y(_00288_),
    .A(net445));
 sg13g2_a22oi_1 _07936_ (.Y(_02019_),
    .B1(net1354),
    .B2(net436),
    .A2(net1377),
    .A1(net1635));
 sg13g2_inv_1 _07937_ (.Y(_00289_),
    .A(net437));
 sg13g2_a22oi_1 _07938_ (.Y(_02020_),
    .B1(net1353),
    .B2(net609),
    .A2(net1380),
    .A1(net1628));
 sg13g2_inv_1 _07939_ (.Y(_00290_),
    .A(_02020_));
 sg13g2_a22oi_1 _07940_ (.Y(_02021_),
    .B1(net1352),
    .B2(net375),
    .A2(net1375),
    .A1(net1627));
 sg13g2_inv_1 _07941_ (.Y(_00291_),
    .A(net376));
 sg13g2_a22oi_1 _07942_ (.Y(_02022_),
    .B1(net1354),
    .B2(net612),
    .A2(net1377),
    .A1(net1616));
 sg13g2_inv_1 _07943_ (.Y(_00292_),
    .A(net613));
 sg13g2_a22oi_1 _07944_ (.Y(_02023_),
    .B1(net1352),
    .B2(net412),
    .A2(net1381),
    .A1(net1615));
 sg13g2_inv_1 _07945_ (.Y(_00293_),
    .A(net413));
 sg13g2_a22oi_1 _07946_ (.Y(_02024_),
    .B1(net1352),
    .B2(net494),
    .A2(net1375),
    .A1(net1611));
 sg13g2_inv_1 _07947_ (.Y(_00294_),
    .A(net495));
 sg13g2_a22oi_1 _07948_ (.Y(_02025_),
    .B1(net1353),
    .B2(net516),
    .A2(net1376),
    .A1(net1606));
 sg13g2_inv_1 _07949_ (.Y(_00295_),
    .A(net517));
 sg13g2_a22oi_1 _07950_ (.Y(_02026_),
    .B1(net1350),
    .B2(net414),
    .A2(net1373),
    .A1(net1602));
 sg13g2_inv_1 _07951_ (.Y(_00296_),
    .A(net415));
 sg13g2_a22oi_1 _07952_ (.Y(_02027_),
    .B1(net1350),
    .B2(net511),
    .A2(net1373),
    .A1(net1597));
 sg13g2_inv_1 _07953_ (.Y(_00297_),
    .A(net512));
 sg13g2_a22oi_1 _07954_ (.Y(_02028_),
    .B1(net1350),
    .B2(net449),
    .A2(net1373),
    .A1(net1590));
 sg13g2_inv_1 _07955_ (.Y(_00298_),
    .A(net450));
 sg13g2_a22oi_1 _07956_ (.Y(_02029_),
    .B1(net1351),
    .B2(net502),
    .A2(net1374),
    .A1(net1583));
 sg13g2_inv_1 _07957_ (.Y(_00299_),
    .A(net503));
 sg13g2_a22oi_1 _07958_ (.Y(_02030_),
    .B1(net1350),
    .B2(net464),
    .A2(net1373),
    .A1(net1578));
 sg13g2_inv_1 _07959_ (.Y(_00300_),
    .A(net465));
 sg13g2_a22oi_1 _07960_ (.Y(_02031_),
    .B1(net1350),
    .B2(net455),
    .A2(net1373),
    .A1(net1573));
 sg13g2_inv_1 _07961_ (.Y(_00301_),
    .A(net456));
 sg13g2_a22oi_1 _07962_ (.Y(_02032_),
    .B1(net1350),
    .B2(net391),
    .A2(net1373),
    .A1(net1569));
 sg13g2_inv_1 _07963_ (.Y(_00302_),
    .A(net392));
 sg13g2_a22oi_1 _07964_ (.Y(_02033_),
    .B1(net1352),
    .B2(net489),
    .A2(net1375),
    .A1(net1565));
 sg13g2_inv_1 _07965_ (.Y(_00303_),
    .A(net490));
 sg13g2_a22oi_1 _07966_ (.Y(_02034_),
    .B1(net1351),
    .B2(net513),
    .A2(net1374),
    .A1(net1513));
 sg13g2_inv_1 _07967_ (.Y(_00304_),
    .A(net514));
 sg13g2_a22oi_1 _07968_ (.Y(_02035_),
    .B1(net1353),
    .B2(net546),
    .A2(net1376),
    .A1(\cordic_inst.MUX_cordic_state$write_1__VAL_1[49] ));
 sg13g2_inv_1 _07969_ (.Y(_00305_),
    .A(net547));
 sg13g2_a22oi_1 _07970_ (.Y(_02036_),
    .B1(net1351),
    .B2(net457),
    .A2(net1374),
    .A1(net1506));
 sg13g2_inv_1 _07971_ (.Y(_00306_),
    .A(net458));
 sg13g2_a22oi_1 _07972_ (.Y(_02037_),
    .B1(net1352),
    .B2(net518),
    .A2(net1375),
    .A1(net1502));
 sg13g2_inv_1 _07973_ (.Y(_00307_),
    .A(net519));
 sg13g2_a22oi_1 _07974_ (.Y(_02038_),
    .B1(net1354),
    .B2(net555),
    .A2(net1377),
    .A1(net1499));
 sg13g2_inv_1 _07975_ (.Y(_00308_),
    .A(net556));
 sg13g2_a22oi_1 _07976_ (.Y(_02039_),
    .B1(net1354),
    .B2(net470),
    .A2(net1377),
    .A1(net1496));
 sg13g2_inv_1 _07977_ (.Y(_00309_),
    .A(net471));
 sg13g2_a22oi_1 _07978_ (.Y(_02040_),
    .B1(net1355),
    .B2(net422),
    .A2(net1378),
    .A1(net1492));
 sg13g2_inv_1 _07979_ (.Y(_00310_),
    .A(net423));
 sg13g2_a22oi_1 _07980_ (.Y(_02041_),
    .B1(net1355),
    .B2(net528),
    .A2(net1378),
    .A1(net1486));
 sg13g2_inv_1 _07981_ (.Y(_00311_),
    .A(net529));
 sg13g2_nand2_1 _07982_ (.Y(_02042_),
    .A(net1626),
    .B(net1535));
 sg13g2_nand2_1 _07983_ (.Y(_02043_),
    .A(net1617),
    .B(net1529));
 sg13g2_nand2_1 _07984_ (.Y(_02044_),
    .A(net1617),
    .B(net1535));
 sg13g2_nand2_1 _07985_ (.Y(_02045_),
    .A(net1626),
    .B(net1529));
 sg13g2_or2_1 _07986_ (.X(_02046_),
    .B(_02043_),
    .A(_02042_));
 sg13g2_nand2_1 _07987_ (.Y(_02047_),
    .A(net1613),
    .B(net1539));
 sg13g2_xnor2_1 _07988_ (.Y(_02048_),
    .A(_02044_),
    .B(_02045_));
 sg13g2_o21ai_1 _07989_ (.B1(_02046_),
    .Y(_02049_),
    .A1(_02047_),
    .A2(_02048_));
 sg13g2_nand2_1 _07990_ (.Y(_02050_),
    .A(net1601),
    .B(net1551));
 sg13g2_nand2_1 _07991_ (.Y(_02051_),
    .A(net1610),
    .B(net1546));
 sg13g2_nand2_1 _07992_ (.Y(_02052_),
    .A(net1604),
    .B(net1538));
 sg13g2_nand2_1 _07993_ (.Y(_02053_),
    .A(net1604),
    .B(net1545));
 sg13g2_nand2_1 _07994_ (.Y(_02054_),
    .A(net1609),
    .B(net1538));
 sg13g2_xor2_1 _07995_ (.B(_02054_),
    .A(_02053_),
    .X(_02055_));
 sg13g2_nand2b_1 _07996_ (.Y(_02056_),
    .B(_02055_),
    .A_N(_02050_));
 sg13g2_xnor2_1 _07997_ (.Y(_02057_),
    .A(_02050_),
    .B(_02055_));
 sg13g2_nand2_1 _07998_ (.Y(_02058_),
    .A(net1606),
    .B(net1552));
 sg13g2_nand2_1 _07999_ (.Y(_02059_),
    .A(net1601),
    .B(net1555));
 sg13g2_xor2_1 _08000_ (.B(_02058_),
    .A(_02051_),
    .X(_02060_));
 sg13g2_nand2b_1 _08001_ (.Y(_02061_),
    .B(_02060_),
    .A_N(_02059_));
 sg13g2_o21ai_1 _08002_ (.B1(_02061_),
    .Y(_02062_),
    .A1(_02051_),
    .A2(_02058_));
 sg13g2_xnor2_1 _08003_ (.Y(_02063_),
    .A(_02049_),
    .B(_02057_));
 sg13g2_nor2b_1 _08004_ (.A(_02063_),
    .B_N(_02062_),
    .Y(_02064_));
 sg13g2_a21o_1 _08005_ (.A2(_02057_),
    .A1(_02049_),
    .B1(_02064_),
    .X(_02065_));
 sg13g2_nand2_2 _08006_ (.Y(_02066_),
    .A(net1596),
    .B(net1555));
 sg13g2_nand2_2 _08007_ (.Y(_02067_),
    .A(net1587),
    .B(net1551));
 sg13g2_nor2_2 _08008_ (.A(_02066_),
    .B(_02067_),
    .Y(_02068_));
 sg13g2_a22oi_1 _08009_ (.Y(_02069_),
    .B1(net1555),
    .B2(net1589),
    .A2(net1551),
    .A1(net1596));
 sg13g2_nor2_1 _08010_ (.A(_02068_),
    .B(_02069_),
    .Y(_02070_));
 sg13g2_nand2_1 _08011_ (.Y(_02071_),
    .A(_02065_),
    .B(_02070_));
 sg13g2_and4_1 _08012_ (.A(net1634),
    .B(net1644),
    .C(net1518),
    .D(net1523),
    .X(_02072_));
 sg13g2_nand4_1 _08013_ (.B(net1645),
    .C(net1518),
    .A(net1634),
    .Y(_02073_),
    .D(net1523));
 sg13g2_nand2_1 _08014_ (.Y(_02074_),
    .A(net1628),
    .B(net1529));
 sg13g2_a22oi_1 _08015_ (.Y(_02075_),
    .B1(net1523),
    .B2(net1634),
    .A2(net1518),
    .A1(net1645));
 sg13g2_or3_1 _08016_ (.A(_02072_),
    .B(_02074_),
    .C(_02075_),
    .X(_02076_));
 sg13g2_o21ai_1 _08017_ (.B1(_02073_),
    .Y(_02077_),
    .A1(_02074_),
    .A2(_02075_));
 sg13g2_nand2_1 _08018_ (.Y(_02078_),
    .A(net1628),
    .B(net1523));
 sg13g2_and4_1 _08019_ (.A(net1634),
    .B(net1653),
    .C(net1732),
    .D(net1518),
    .X(_02079_));
 sg13g2_nand4_1 _08020_ (.B(net1653),
    .C(net1732),
    .A(net1634),
    .Y(_02080_),
    .D(net1516));
 sg13g2_a22oi_1 _08021_ (.Y(_02081_),
    .B1(net1516),
    .B2(net1634),
    .A2(net1732),
    .A1(net1653));
 sg13g2_or3_1 _08022_ (.A(_02078_),
    .B(_02079_),
    .C(_02081_),
    .X(_02082_));
 sg13g2_o21ai_1 _08023_ (.B1(_02078_),
    .Y(_02083_),
    .A1(_02079_),
    .A2(_02081_));
 sg13g2_and3_1 _08024_ (.X(_02084_),
    .A(_02077_),
    .B(_02082_),
    .C(_02083_));
 sg13g2_nand3_1 _08025_ (.B(_02082_),
    .C(_02083_),
    .A(_02077_),
    .Y(_02085_));
 sg13g2_a21o_1 _08026_ (.A2(_02083_),
    .A1(_02082_),
    .B1(_02077_),
    .X(_02086_));
 sg13g2_xor2_1 _08027_ (.B(_02048_),
    .A(_02047_),
    .X(_02087_));
 sg13g2_nand3_1 _08028_ (.B(_02086_),
    .C(_02087_),
    .A(_02085_),
    .Y(_02088_));
 sg13g2_a21o_1 _08029_ (.A2(_02087_),
    .A1(_02086_),
    .B1(_02084_),
    .X(_02089_));
 sg13g2_o21ai_1 _08030_ (.B1(_02080_),
    .Y(_02090_),
    .A1(_02078_),
    .A2(_02081_));
 sg13g2_nand2_1 _08031_ (.Y(_02091_),
    .A(net1630),
    .B(net1516));
 sg13g2_and4_1 _08032_ (.A(net1643),
    .B(net1653),
    .C(net1726),
    .D(net1732),
    .X(_02092_));
 sg13g2_nand4_1 _08033_ (.B(net1653),
    .C(net1723),
    .A(net1643),
    .Y(_02093_),
    .D(net1730));
 sg13g2_a22oi_1 _08034_ (.Y(_02094_),
    .B1(net1732),
    .B2(net1643),
    .A2(net1723),
    .A1(net1653));
 sg13g2_or3_1 _08035_ (.A(_02091_),
    .B(_02092_),
    .C(_02094_),
    .X(_02095_));
 sg13g2_o21ai_1 _08036_ (.B1(_02091_),
    .Y(_02096_),
    .A1(_02092_),
    .A2(_02094_));
 sg13g2_and3_1 _08037_ (.X(_02097_),
    .A(_02090_),
    .B(_02095_),
    .C(_02096_));
 sg13g2_nand3_1 _08038_ (.B(_02095_),
    .C(_02096_),
    .A(_02090_),
    .Y(_02098_));
 sg13g2_a21oi_1 _08039_ (.A1(_02095_),
    .A2(_02096_),
    .Y(_02099_),
    .B1(_02090_));
 sg13g2_nand2_1 _08040_ (.Y(_02100_),
    .A(net1613),
    .B(net1533));
 sg13g2_nand2_1 _08041_ (.Y(_02101_),
    .A(net1626),
    .B(net1523));
 sg13g2_or2_1 _08042_ (.X(_02102_),
    .B(_02101_),
    .A(_02043_));
 sg13g2_xnor2_1 _08043_ (.Y(_02103_),
    .A(_02043_),
    .B(_02101_));
 sg13g2_xnor2_1 _08044_ (.Y(_02104_),
    .A(_02100_),
    .B(_02103_));
 sg13g2_or3_1 _08045_ (.A(_02097_),
    .B(_02099_),
    .C(_02104_),
    .X(_02105_));
 sg13g2_o21ai_1 _08046_ (.B1(_02104_),
    .Y(_02106_),
    .A1(_02097_),
    .A2(_02099_));
 sg13g2_and3_1 _08047_ (.X(_02107_),
    .A(_02089_),
    .B(_02105_),
    .C(_02106_));
 sg13g2_nand3_1 _08048_ (.B(_02105_),
    .C(_02106_),
    .A(_02089_),
    .Y(_02108_));
 sg13g2_a21oi_1 _08049_ (.A1(_02105_),
    .A2(_02106_),
    .Y(_02109_),
    .B1(_02089_));
 sg13g2_xor2_1 _08050_ (.B(_02063_),
    .A(_02062_),
    .X(_02110_));
 sg13g2_or3_1 _08051_ (.A(_02107_),
    .B(_02109_),
    .C(_02110_),
    .X(_02111_));
 sg13g2_o21ai_1 _08052_ (.B1(_02108_),
    .Y(_02112_),
    .A1(_02109_),
    .A2(_02110_));
 sg13g2_o21ai_1 _08053_ (.B1(_02098_),
    .Y(_02113_),
    .A1(_02099_),
    .A2(_02104_));
 sg13g2_o21ai_1 _08054_ (.B1(_02093_),
    .Y(_02114_),
    .A1(_02091_),
    .A2(_02094_));
 sg13g2_nand2_1 _08055_ (.Y(_02115_),
    .A(net1630),
    .B(net1730));
 sg13g2_and4_1 _08056_ (.A(net1643),
    .B(net1653),
    .C(net1717),
    .D(net1723),
    .X(_02116_));
 sg13g2_nand4_1 _08057_ (.B(net1651),
    .C(net1717),
    .A(net1643),
    .Y(_02117_),
    .D(net1723));
 sg13g2_a22oi_1 _08058_ (.Y(_02118_),
    .B1(net1723),
    .B2(net1643),
    .A2(net1717),
    .A1(net1653));
 sg13g2_or3_1 _08059_ (.A(_02115_),
    .B(_02116_),
    .C(_02118_),
    .X(_02119_));
 sg13g2_o21ai_1 _08060_ (.B1(_02115_),
    .Y(_02120_),
    .A1(_02116_),
    .A2(_02118_));
 sg13g2_and3_1 _08061_ (.X(_02121_),
    .A(_02114_),
    .B(_02119_),
    .C(_02120_));
 sg13g2_nand3_1 _08062_ (.B(_02119_),
    .C(_02120_),
    .A(_02114_),
    .Y(_02122_));
 sg13g2_a21oi_1 _08063_ (.A1(_02119_),
    .A2(_02120_),
    .Y(_02123_),
    .B1(_02114_));
 sg13g2_nand2_1 _08064_ (.Y(_02124_),
    .A(net1613),
    .B(net1529));
 sg13g2_nand2_1 _08065_ (.Y(_02125_),
    .A(net1621),
    .B(net1516));
 sg13g2_and4_1 _08066_ (.A(net1621),
    .B(net1626),
    .C(net1516),
    .D(net1521),
    .X(_02126_));
 sg13g2_a22oi_1 _08067_ (.Y(_02127_),
    .B1(net1521),
    .B2(net1621),
    .A2(net1517),
    .A1(net1626));
 sg13g2_nor3_1 _08068_ (.A(_02124_),
    .B(_02126_),
    .C(_02127_),
    .Y(_02128_));
 sg13g2_o21ai_1 _08069_ (.B1(_02124_),
    .Y(_02129_),
    .A1(_02126_),
    .A2(_02127_));
 sg13g2_nand2b_1 _08070_ (.Y(_02130_),
    .B(_02129_),
    .A_N(_02128_));
 sg13g2_or3_1 _08071_ (.A(_02121_),
    .B(_02123_),
    .C(_02130_),
    .X(_02131_));
 sg13g2_o21ai_1 _08072_ (.B1(_02130_),
    .Y(_02132_),
    .A1(_02121_),
    .A2(_02123_));
 sg13g2_and3_1 _08073_ (.X(_02133_),
    .A(_02113_),
    .B(_02131_),
    .C(_02132_));
 sg13g2_nand3_1 _08074_ (.B(_02131_),
    .C(_02132_),
    .A(_02113_),
    .Y(_02134_));
 sg13g2_a21oi_1 _08075_ (.A1(_02131_),
    .A2(_02132_),
    .Y(_02135_),
    .B1(_02113_));
 sg13g2_o21ai_1 _08076_ (.B1(_02056_),
    .Y(_02136_),
    .A1(_02053_),
    .A2(_02054_));
 sg13g2_o21ai_1 _08077_ (.B1(_02102_),
    .Y(_02137_),
    .A1(_02100_),
    .A2(_02103_));
 sg13g2_nand2_1 _08078_ (.Y(_02138_),
    .A(net1599),
    .B(net1545));
 sg13g2_nand2_1 _08079_ (.Y(_02139_),
    .A(net1604),
    .B(net1534));
 sg13g2_nand2_1 _08080_ (.Y(_02140_),
    .A(net1609),
    .B(net1534));
 sg13g2_or2_1 _08081_ (.X(_02141_),
    .B(_02139_),
    .A(_02054_));
 sg13g2_xor2_1 _08082_ (.B(_02140_),
    .A(_02052_),
    .X(_02142_));
 sg13g2_nand2b_1 _08083_ (.Y(_02143_),
    .B(_02142_),
    .A_N(_02138_));
 sg13g2_xnor2_1 _08084_ (.Y(_02144_),
    .A(_02138_),
    .B(_02142_));
 sg13g2_xnor2_1 _08085_ (.Y(_02145_),
    .A(_02137_),
    .B(_02144_));
 sg13g2_nor2b_1 _08086_ (.A(_02145_),
    .B_N(_02136_),
    .Y(_02146_));
 sg13g2_xor2_1 _08087_ (.B(_02145_),
    .A(_02136_),
    .X(_02147_));
 sg13g2_or3_1 _08088_ (.A(_02133_),
    .B(_02135_),
    .C(_02147_),
    .X(_02148_));
 sg13g2_o21ai_1 _08089_ (.B1(_02147_),
    .Y(_02149_),
    .A1(_02133_),
    .A2(_02135_));
 sg13g2_and3_1 _08090_ (.X(_02150_),
    .A(_02112_),
    .B(_02148_),
    .C(_02149_));
 sg13g2_nand3_1 _08091_ (.B(_02148_),
    .C(_02149_),
    .A(_02112_),
    .Y(_02151_));
 sg13g2_xnor2_1 _08092_ (.Y(_02152_),
    .A(_02065_),
    .B(_02070_));
 sg13g2_a21oi_1 _08093_ (.A1(_02148_),
    .A2(_02149_),
    .Y(_02153_),
    .B1(_02112_));
 sg13g2_or3_1 _08094_ (.A(_02150_),
    .B(_02152_),
    .C(_02153_),
    .X(_02154_));
 sg13g2_o21ai_1 _08095_ (.B1(_02151_),
    .Y(_02155_),
    .A1(_02152_),
    .A2(_02153_));
 sg13g2_a21o_1 _08096_ (.A2(_02144_),
    .A1(_02137_),
    .B1(_02146_),
    .X(_02156_));
 sg13g2_and2_1 _08097_ (.A(net1581),
    .B(net1555),
    .X(_02157_));
 sg13g2_nand2_1 _08098_ (.Y(_02158_),
    .A(net1594),
    .B(net1545));
 sg13g2_nor2_1 _08099_ (.A(_02067_),
    .B(_02158_),
    .Y(_02159_));
 sg13g2_xor2_1 _08100_ (.B(_02158_),
    .A(_02067_),
    .X(_02160_));
 sg13g2_xor2_1 _08101_ (.B(_02160_),
    .A(_02157_),
    .X(_02161_));
 sg13g2_nand2_1 _08102_ (.Y(_02162_),
    .A(_02068_),
    .B(_02161_));
 sg13g2_xor2_1 _08103_ (.B(_02161_),
    .A(_02068_),
    .X(_02163_));
 sg13g2_nand2_1 _08104_ (.Y(_02164_),
    .A(_02156_),
    .B(_02163_));
 sg13g2_xnor2_1 _08105_ (.Y(_02165_),
    .A(_02156_),
    .B(_02163_));
 sg13g2_o21ai_1 _08106_ (.B1(_02134_),
    .Y(_02166_),
    .A1(_02135_),
    .A2(_02147_));
 sg13g2_o21ai_1 _08107_ (.B1(_02122_),
    .Y(_02167_),
    .A1(_02123_),
    .A2(_02130_));
 sg13g2_o21ai_1 _08108_ (.B1(_02117_),
    .Y(_02168_),
    .A1(_02115_),
    .A2(_02118_));
 sg13g2_nand2_1 _08109_ (.Y(_02169_),
    .A(net1630),
    .B(net1723));
 sg13g2_and4_1 _08110_ (.A(net1641),
    .B(net1651),
    .C(net1712),
    .D(net1717),
    .X(_02170_));
 sg13g2_nand4_1 _08111_ (.B(net1650),
    .C(net1712),
    .A(net1641),
    .Y(_02171_),
    .D(net1718));
 sg13g2_a22oi_1 _08112_ (.Y(_02172_),
    .B1(net1718),
    .B2(net1641),
    .A2(net1712),
    .A1(net1651));
 sg13g2_or3_1 _08113_ (.A(_02169_),
    .B(_02170_),
    .C(_02172_),
    .X(_02173_));
 sg13g2_o21ai_1 _08114_ (.B1(_02169_),
    .Y(_02174_),
    .A1(_02170_),
    .A2(_02172_));
 sg13g2_and3_1 _08115_ (.X(_02175_),
    .A(_02168_),
    .B(_02173_),
    .C(_02174_));
 sg13g2_nand3_1 _08116_ (.B(_02173_),
    .C(_02174_),
    .A(_02168_),
    .Y(_02176_));
 sg13g2_a21oi_1 _08117_ (.A1(_02173_),
    .A2(_02174_),
    .Y(_02177_),
    .B1(_02168_));
 sg13g2_nand2_1 _08118_ (.Y(_02178_),
    .A(net1614),
    .B(net1522));
 sg13g2_nand2_1 _08119_ (.Y(_02179_),
    .A(net1626),
    .B(net1730));
 sg13g2_or2_1 _08120_ (.X(_02180_),
    .B(_02179_),
    .A(_02125_));
 sg13g2_and2_1 _08121_ (.A(_02125_),
    .B(_02179_),
    .X(_02181_));
 sg13g2_xnor2_1 _08122_ (.Y(_02182_),
    .A(_02125_),
    .B(_02179_));
 sg13g2_xnor2_1 _08123_ (.Y(_02183_),
    .A(_02178_),
    .B(_02182_));
 sg13g2_or3_1 _08124_ (.A(_02175_),
    .B(_02177_),
    .C(_02183_),
    .X(_02184_));
 sg13g2_o21ai_1 _08125_ (.B1(_02183_),
    .Y(_02185_),
    .A1(_02175_),
    .A2(_02177_));
 sg13g2_and3_1 _08126_ (.X(_02186_),
    .A(_02167_),
    .B(_02184_),
    .C(_02185_));
 sg13g2_nand3_1 _08127_ (.B(_02184_),
    .C(_02185_),
    .A(_02167_),
    .Y(_02187_));
 sg13g2_a21oi_1 _08128_ (.A1(_02184_),
    .A2(_02185_),
    .Y(_02188_),
    .B1(_02167_));
 sg13g2_and2_1 _08129_ (.A(_02141_),
    .B(_02143_),
    .X(_02189_));
 sg13g2_or2_1 _08130_ (.X(_02190_),
    .B(_02128_),
    .A(_02126_));
 sg13g2_nand2_1 _08131_ (.Y(_02191_),
    .A(net1599),
    .B(net1538));
 sg13g2_nand2_1 _08132_ (.Y(_02192_),
    .A(net1604),
    .B(net1528));
 sg13g2_nand2_1 _08133_ (.Y(_02193_),
    .A(net1609),
    .B(net1528));
 sg13g2_or2_1 _08134_ (.X(_02194_),
    .B(_02192_),
    .A(_02140_));
 sg13g2_xnor2_1 _08135_ (.Y(_02195_),
    .A(_02139_),
    .B(_02193_));
 sg13g2_xor2_1 _08136_ (.B(_02195_),
    .A(_02191_),
    .X(_02196_));
 sg13g2_nand2_1 _08137_ (.Y(_02197_),
    .A(_02190_),
    .B(_02196_));
 sg13g2_xnor2_1 _08138_ (.Y(_02198_),
    .A(_02190_),
    .B(_02196_));
 sg13g2_xnor2_1 _08139_ (.Y(_02199_),
    .A(_02189_),
    .B(_02198_));
 sg13g2_or3_1 _08140_ (.A(_02186_),
    .B(_02188_),
    .C(_02199_),
    .X(_02200_));
 sg13g2_o21ai_1 _08141_ (.B1(_02199_),
    .Y(_02201_),
    .A1(_02186_),
    .A2(_02188_));
 sg13g2_and3_1 _08142_ (.X(_02202_),
    .A(_02166_),
    .B(_02200_),
    .C(_02201_));
 sg13g2_nand3_1 _08143_ (.B(_02200_),
    .C(_02201_),
    .A(_02166_),
    .Y(_02203_));
 sg13g2_a21oi_1 _08144_ (.A1(_02200_),
    .A2(_02201_),
    .Y(_02204_),
    .B1(_02166_));
 sg13g2_or3_1 _08145_ (.A(_02165_),
    .B(_02202_),
    .C(_02204_),
    .X(_02205_));
 sg13g2_o21ai_1 _08146_ (.B1(_02165_),
    .Y(_02206_),
    .A1(_02202_),
    .A2(_02204_));
 sg13g2_and3_1 _08147_ (.X(_02207_),
    .A(_02155_),
    .B(_02205_),
    .C(_02206_));
 sg13g2_nand3_1 _08148_ (.B(_02205_),
    .C(_02206_),
    .A(_02155_),
    .Y(_02208_));
 sg13g2_a21oi_1 _08149_ (.A1(_02205_),
    .A2(_02206_),
    .Y(_02209_),
    .B1(_02155_));
 sg13g2_o21ai_1 _08150_ (.B1(_02071_),
    .Y(_02210_),
    .A1(_02207_),
    .A2(_02209_));
 sg13g2_or3_1 _08151_ (.A(_02071_),
    .B(_02207_),
    .C(_02209_),
    .X(_02211_));
 sg13g2_and4_1 _08152_ (.A(net1633),
    .B(net1644),
    .C(net1523),
    .D(net1526),
    .X(_02212_));
 sg13g2_nand4_1 _08153_ (.B(net1644),
    .C(net1523),
    .A(net1633),
    .Y(_02213_),
    .D(net1526));
 sg13g2_nand2_1 _08154_ (.Y(_02214_),
    .A(net1628),
    .B(net1531));
 sg13g2_a22oi_1 _08155_ (.Y(_02215_),
    .B1(net1526),
    .B2(net1633),
    .A2(net1523),
    .A1(net1644));
 sg13g2_nor3_1 _08156_ (.A(_02212_),
    .B(_02214_),
    .C(_02215_),
    .Y(_02216_));
 sg13g2_o21ai_1 _08157_ (.B1(_02213_),
    .Y(_02217_),
    .A1(_02214_),
    .A2(_02215_));
 sg13g2_o21ai_1 _08158_ (.B1(_02074_),
    .Y(_02218_),
    .A1(_02072_),
    .A2(_02075_));
 sg13g2_and3_1 _08159_ (.X(_02219_),
    .A(_02076_),
    .B(_02217_),
    .C(_02218_));
 sg13g2_a21o_1 _08160_ (.A2(_02218_),
    .A1(_02076_),
    .B1(_02217_),
    .X(_02220_));
 sg13g2_nand2b_1 _08161_ (.Y(_02221_),
    .B(_02220_),
    .A_N(_02219_));
 sg13g2_nand2_1 _08162_ (.Y(_02222_),
    .A(net1615),
    .B(net1546));
 sg13g2_nand2_1 _08163_ (.Y(_02223_),
    .A(net1627),
    .B(net1539));
 sg13g2_nand2_1 _08164_ (.Y(_02224_),
    .A(net1616),
    .B(net1539));
 sg13g2_or2_1 _08165_ (.X(_02225_),
    .B(_02223_),
    .A(_02044_));
 sg13g2_xnor2_1 _08166_ (.Y(_02226_),
    .A(_02042_),
    .B(_02224_));
 sg13g2_xor2_1 _08167_ (.B(_02226_),
    .A(_02222_),
    .X(_02227_));
 sg13g2_a21o_1 _08168_ (.A2(_02227_),
    .A1(_02220_),
    .B1(_02219_),
    .X(_02228_));
 sg13g2_a21o_1 _08169_ (.A2(_02086_),
    .A1(_02085_),
    .B1(_02087_),
    .X(_02229_));
 sg13g2_and3_1 _08170_ (.X(_02230_),
    .A(_02088_),
    .B(_02228_),
    .C(_02229_));
 sg13g2_a21o_1 _08171_ (.A2(_02229_),
    .A1(_02088_),
    .B1(_02228_),
    .X(_02231_));
 sg13g2_nand2b_1 _08172_ (.Y(_02232_),
    .B(_02231_),
    .A_N(_02230_));
 sg13g2_nand2_2 _08173_ (.Y(_02233_),
    .A(net1610),
    .B(net1557));
 sg13g2_or2_1 _08174_ (.X(_02234_),
    .B(_02233_),
    .A(_02058_));
 sg13g2_inv_1 _08175_ (.Y(_02235_),
    .A(_02234_));
 sg13g2_o21ai_1 _08176_ (.B1(_02225_),
    .Y(_02236_),
    .A1(_02222_),
    .A2(_02226_));
 sg13g2_xnor2_1 _08177_ (.Y(_02237_),
    .A(_02059_),
    .B(_02060_));
 sg13g2_nand2_1 _08178_ (.Y(_02238_),
    .A(_02236_),
    .B(_02237_));
 sg13g2_xnor2_1 _08179_ (.Y(_02239_),
    .A(_02236_),
    .B(_02237_));
 sg13g2_xnor2_1 _08180_ (.Y(_02240_),
    .A(_02235_),
    .B(_02239_));
 sg13g2_a21o_1 _08181_ (.A2(_02240_),
    .A1(_02231_),
    .B1(_02230_),
    .X(_02241_));
 sg13g2_o21ai_1 _08182_ (.B1(_02110_),
    .Y(_02242_),
    .A1(_02107_),
    .A2(_02109_));
 sg13g2_and3_1 _08183_ (.X(_02243_),
    .A(_02111_),
    .B(_02241_),
    .C(_02242_));
 sg13g2_nand3_1 _08184_ (.B(_02241_),
    .C(_02242_),
    .A(_02111_),
    .Y(_02244_));
 sg13g2_o21ai_1 _08185_ (.B1(_02238_),
    .Y(_02245_),
    .A1(_02234_),
    .A2(_02239_));
 sg13g2_nand2b_1 _08186_ (.Y(_02246_),
    .B(_02245_),
    .A_N(_02066_));
 sg13g2_xor2_1 _08187_ (.B(_02245_),
    .A(_02066_),
    .X(_02247_));
 sg13g2_a21oi_1 _08188_ (.A1(_02111_),
    .A2(_02242_),
    .Y(_02248_),
    .B1(_02241_));
 sg13g2_nor2_1 _08189_ (.A(_02243_),
    .B(_02248_),
    .Y(_02249_));
 sg13g2_o21ai_1 _08190_ (.B1(_02244_),
    .Y(_02250_),
    .A1(_02247_),
    .A2(_02248_));
 sg13g2_o21ai_1 _08191_ (.B1(_02152_),
    .Y(_02251_),
    .A1(_02150_),
    .A2(_02153_));
 sg13g2_and3_1 _08192_ (.X(_02252_),
    .A(_02154_),
    .B(_02250_),
    .C(_02251_));
 sg13g2_nand3_1 _08193_ (.B(_02250_),
    .C(_02251_),
    .A(_02154_),
    .Y(_02253_));
 sg13g2_a21oi_1 _08194_ (.A1(_02154_),
    .A2(_02251_),
    .Y(_02254_),
    .B1(_02250_));
 sg13g2_nor3_1 _08195_ (.A(_02246_),
    .B(_02252_),
    .C(_02254_),
    .Y(_02255_));
 sg13g2_o21ai_1 _08196_ (.B1(_02253_),
    .Y(_02256_),
    .A1(_02246_),
    .A2(_02254_));
 sg13g2_and3_2 _08197_ (.X(_02257_),
    .A(_02210_),
    .B(_02211_),
    .C(_02256_));
 sg13g2_nand3_1 _08198_ (.B(_02211_),
    .C(_02256_),
    .A(_02210_),
    .Y(_02258_));
 sg13g2_a21oi_2 _08199_ (.B1(_02256_),
    .Y(_02259_),
    .A2(_02211_),
    .A1(_02210_));
 sg13g2_o21ai_1 _08200_ (.B1(_02246_),
    .Y(_02260_),
    .A1(_02252_),
    .A2(_02254_));
 sg13g2_nor2b_1 _08201_ (.A(_02255_),
    .B_N(_02260_),
    .Y(_02261_));
 sg13g2_nand2_1 _08202_ (.Y(_02262_),
    .A(net1645),
    .B(net1539));
 sg13g2_and4_1 _08203_ (.A(net1633),
    .B(net1644),
    .C(net1531),
    .D(net1541),
    .X(_02263_));
 sg13g2_nand2_1 _08204_ (.Y(_02264_),
    .A(net1628),
    .B(net1546));
 sg13g2_a22oi_1 _08205_ (.Y(_02265_),
    .B1(net1541),
    .B2(net1633),
    .A2(net1531),
    .A1(net1644));
 sg13g2_nor3_1 _08206_ (.A(_02263_),
    .B(_02264_),
    .C(_02265_),
    .Y(_02266_));
 sg13g2_or2_1 _08207_ (.X(_02267_),
    .B(_02266_),
    .A(_02263_));
 sg13g2_nand2_1 _08208_ (.Y(_02268_),
    .A(net1628),
    .B(net1541));
 sg13g2_and4_1 _08209_ (.A(net1633),
    .B(net1644),
    .C(net1526),
    .D(net1536),
    .X(_02269_));
 sg13g2_a22oi_1 _08210_ (.Y(_02270_),
    .B1(net1536),
    .B2(net1633),
    .A2(\cordic_inst.MUX_cordic_state$write_1__VAL_1[61] ),
    .A1(net1644));
 sg13g2_nor3_1 _08211_ (.A(_02268_),
    .B(_02269_),
    .C(_02270_),
    .Y(_02271_));
 sg13g2_o21ai_1 _08212_ (.B1(_02268_),
    .Y(_02272_),
    .A1(_02269_),
    .A2(_02270_));
 sg13g2_nor2b_1 _08213_ (.A(_02271_),
    .B_N(_02272_),
    .Y(_02273_));
 sg13g2_nand2_1 _08214_ (.Y(_02274_),
    .A(_02267_),
    .B(_02273_));
 sg13g2_nand2_1 _08215_ (.Y(_02275_),
    .A(net1615),
    .B(net1557));
 sg13g2_nand2_1 _08216_ (.Y(_02276_),
    .A(net1617),
    .B(net1546));
 sg13g2_nand2_1 _08217_ (.Y(_02277_),
    .A(net1627),
    .B(net1546));
 sg13g2_nand2_2 _08218_ (.Y(_02278_),
    .A(net1617),
    .B(net1554));
 sg13g2_xnor2_1 _08219_ (.Y(_02279_),
    .A(_02277_),
    .B(_02278_));
 sg13g2_or2_1 _08220_ (.X(_02280_),
    .B(_02279_),
    .A(_02275_));
 sg13g2_xnor2_1 _08221_ (.Y(_02281_),
    .A(_02275_),
    .B(_02279_));
 sg13g2_xnor2_1 _08222_ (.Y(_02282_),
    .A(_02267_),
    .B(_02273_));
 sg13g2_o21ai_1 _08223_ (.B1(_02274_),
    .Y(_02283_),
    .A1(_02281_),
    .A2(_02282_));
 sg13g2_nand2_1 _08224_ (.Y(_02284_),
    .A(net1615),
    .B(net1554));
 sg13g2_or2_1 _08225_ (.X(_02285_),
    .B(_02277_),
    .A(_02224_));
 sg13g2_xnor2_1 _08226_ (.Y(_02286_),
    .A(_02223_),
    .B(_02276_));
 sg13g2_xnor2_1 _08227_ (.Y(_02287_),
    .A(_02284_),
    .B(_02286_));
 sg13g2_or2_1 _08228_ (.X(_02288_),
    .B(_02271_),
    .A(_02269_));
 sg13g2_o21ai_1 _08229_ (.B1(_02214_),
    .Y(_02289_),
    .A1(_02212_),
    .A2(_02215_));
 sg13g2_nor2b_1 _08230_ (.A(_02216_),
    .B_N(_02289_),
    .Y(_02290_));
 sg13g2_nand2_1 _08231_ (.Y(_02291_),
    .A(_02288_),
    .B(_02290_));
 sg13g2_xnor2_1 _08232_ (.Y(_02292_),
    .A(_02288_),
    .B(_02290_));
 sg13g2_xnor2_1 _08233_ (.Y(_02293_),
    .A(_02287_),
    .B(_02292_));
 sg13g2_nand2b_1 _08234_ (.Y(_02294_),
    .B(_02283_),
    .A_N(_02293_));
 sg13g2_o21ai_1 _08235_ (.B1(_02280_),
    .Y(_02295_),
    .A1(_02277_),
    .A2(_02278_));
 sg13g2_nor2b_1 _08236_ (.A(_02233_),
    .B_N(_02295_),
    .Y(_02296_));
 sg13g2_xor2_1 _08237_ (.B(_02295_),
    .A(_02233_),
    .X(_02297_));
 sg13g2_xor2_1 _08238_ (.B(_02293_),
    .A(_02283_),
    .X(_02298_));
 sg13g2_o21ai_1 _08239_ (.B1(_02294_),
    .Y(_02299_),
    .A1(_02297_),
    .A2(_02298_));
 sg13g2_o21ai_1 _08240_ (.B1(_02285_),
    .Y(_02300_),
    .A1(_02284_),
    .A2(_02286_));
 sg13g2_a22oi_1 _08241_ (.Y(_02301_),
    .B1(net1557),
    .B2(net1606),
    .A2(net1552),
    .A1(net1610));
 sg13g2_nor2_1 _08242_ (.A(_02235_),
    .B(_02301_),
    .Y(_02302_));
 sg13g2_nand2_1 _08243_ (.Y(_02303_),
    .A(_02300_),
    .B(_02302_));
 sg13g2_xnor2_1 _08244_ (.Y(_02304_),
    .A(_02300_),
    .B(_02302_));
 sg13g2_o21ai_1 _08245_ (.B1(_02291_),
    .Y(_02305_),
    .A1(_02287_),
    .A2(_02292_));
 sg13g2_xnor2_1 _08246_ (.Y(_02306_),
    .A(_02221_),
    .B(_02227_));
 sg13g2_nand2_1 _08247_ (.Y(_02307_),
    .A(_02305_),
    .B(_02306_));
 sg13g2_xnor2_1 _08248_ (.Y(_02308_),
    .A(_02305_),
    .B(_02306_));
 sg13g2_xor2_1 _08249_ (.B(_02308_),
    .A(_02304_),
    .X(_02309_));
 sg13g2_nand2_1 _08250_ (.Y(_02310_),
    .A(_02299_),
    .B(_02309_));
 sg13g2_xor2_1 _08251_ (.B(_02309_),
    .A(_02299_),
    .X(_02311_));
 sg13g2_nand2_1 _08252_ (.Y(_02312_),
    .A(_02296_),
    .B(_02311_));
 sg13g2_o21ai_1 _08253_ (.B1(_02307_),
    .Y(_02313_),
    .A1(_02304_),
    .A2(_02308_));
 sg13g2_xnor2_1 _08254_ (.Y(_02314_),
    .A(_02232_),
    .B(_02240_));
 sg13g2_nand2_1 _08255_ (.Y(_02315_),
    .A(_02313_),
    .B(_02314_));
 sg13g2_xnor2_1 _08256_ (.Y(_02316_),
    .A(_02313_),
    .B(_02314_));
 sg13g2_xnor2_1 _08257_ (.Y(_02317_),
    .A(_02303_),
    .B(_02316_));
 sg13g2_a21o_1 _08258_ (.A2(_02312_),
    .A1(_02310_),
    .B1(_02317_),
    .X(_02318_));
 sg13g2_xnor2_1 _08259_ (.Y(_02319_),
    .A(_02247_),
    .B(_02249_));
 sg13g2_o21ai_1 _08260_ (.B1(_02315_),
    .Y(_02320_),
    .A1(_02303_),
    .A2(_02316_));
 sg13g2_and2_1 _08261_ (.A(_02319_),
    .B(_02320_),
    .X(_02321_));
 sg13g2_xnor2_1 _08262_ (.Y(_02322_),
    .A(_02319_),
    .B(_02320_));
 sg13g2_nor2_1 _08263_ (.A(_02318_),
    .B(_02322_),
    .Y(_02323_));
 sg13g2_nand2_1 _08264_ (.Y(_02324_),
    .A(_02261_),
    .B(_02323_));
 sg13g2_nor3_1 _08265_ (.A(_02257_),
    .B(_02259_),
    .C(_02324_),
    .Y(_02325_));
 sg13g2_nand3b_1 _08266_ (.B(_02260_),
    .C(_02321_),
    .Y(_02326_),
    .A_N(_02255_));
 sg13g2_o21ai_1 _08267_ (.B1(_02203_),
    .Y(_02327_),
    .A1(_02165_),
    .A2(_02204_));
 sg13g2_o21ai_1 _08268_ (.B1(_02197_),
    .Y(_02328_),
    .A1(_02189_),
    .A2(_02198_));
 sg13g2_nand2_1 _08269_ (.Y(_02329_),
    .A(net1575),
    .B(net1555));
 sg13g2_a21oi_1 _08270_ (.A1(_02157_),
    .A2(_02160_),
    .Y(_02330_),
    .B1(_02159_));
 sg13g2_nand2_1 _08271_ (.Y(_02331_),
    .A(net1581),
    .B(net1551));
 sg13g2_nand2_1 _08272_ (.Y(_02332_),
    .A(net1587),
    .B(net1538));
 sg13g2_and4_1 _08273_ (.A(net1587),
    .B(net1594),
    .C(net1538),
    .D(net1545),
    .X(_02333_));
 sg13g2_a22oi_1 _08274_ (.Y(_02334_),
    .B1(net1547),
    .B2(net1587),
    .A2(net1539),
    .A1(net1594));
 sg13g2_nor3_1 _08275_ (.A(_02331_),
    .B(_02333_),
    .C(_02334_),
    .Y(_02335_));
 sg13g2_o21ai_1 _08276_ (.B1(_02331_),
    .Y(_02336_),
    .A1(_02333_),
    .A2(_02334_));
 sg13g2_nor2b_1 _08277_ (.A(_02335_),
    .B_N(_02336_),
    .Y(_02337_));
 sg13g2_nand2b_1 _08278_ (.Y(_02338_),
    .B(_02337_),
    .A_N(_02330_));
 sg13g2_xnor2_1 _08279_ (.Y(_02339_),
    .A(_02330_),
    .B(_02337_));
 sg13g2_nand2b_1 _08280_ (.Y(_02340_),
    .B(_02339_),
    .A_N(_02329_));
 sg13g2_xnor2_1 _08281_ (.Y(_02341_),
    .A(_02329_),
    .B(_02339_));
 sg13g2_nand2_1 _08282_ (.Y(_02342_),
    .A(_02328_),
    .B(_02341_));
 sg13g2_xnor2_1 _08283_ (.Y(_02343_),
    .A(_02328_),
    .B(_02341_));
 sg13g2_xor2_1 _08284_ (.B(_02343_),
    .A(_02162_),
    .X(_02344_));
 sg13g2_o21ai_1 _08285_ (.B1(_02187_),
    .Y(_02345_),
    .A1(_02188_),
    .A2(_02199_));
 sg13g2_o21ai_1 _08286_ (.B1(_02194_),
    .Y(_02346_),
    .A1(_02191_),
    .A2(_02195_));
 sg13g2_inv_1 _08287_ (.Y(_02347_),
    .A(_02346_));
 sg13g2_o21ai_1 _08288_ (.B1(_02180_),
    .Y(_02348_),
    .A1(_02178_),
    .A2(_02181_));
 sg13g2_nand2_1 _08289_ (.Y(_02349_),
    .A(net1599),
    .B(net1533));
 sg13g2_nand2_1 _08290_ (.Y(_02350_),
    .A(net1604),
    .B(net1522));
 sg13g2_nand2_1 _08291_ (.Y(_02351_),
    .A(net1610),
    .B(net1522));
 sg13g2_or2_1 _08292_ (.X(_02352_),
    .B(_02350_),
    .A(_02193_));
 sg13g2_xnor2_1 _08293_ (.Y(_02353_),
    .A(_02192_),
    .B(_02351_));
 sg13g2_xor2_1 _08294_ (.B(_02353_),
    .A(_02349_),
    .X(_02354_));
 sg13g2_nand2_1 _08295_ (.Y(_02355_),
    .A(_02348_),
    .B(_02354_));
 sg13g2_xnor2_1 _08296_ (.Y(_02356_),
    .A(_02348_),
    .B(_02354_));
 sg13g2_xnor2_1 _08297_ (.Y(_02357_),
    .A(_02347_),
    .B(_02356_));
 sg13g2_o21ai_1 _08298_ (.B1(_02176_),
    .Y(_02358_),
    .A1(_02177_),
    .A2(_02183_));
 sg13g2_nand2_1 _08299_ (.Y(_02359_),
    .A(net1613),
    .B(net1516));
 sg13g2_nand2_1 _08300_ (.Y(_02360_),
    .A(net1620),
    .B(net1724));
 sg13g2_and4_1 _08301_ (.A(net1621),
    .B(net1625),
    .C(net1723),
    .D(net1730),
    .X(_02361_));
 sg13g2_a22oi_1 _08302_ (.Y(_02362_),
    .B1(net1730),
    .B2(net1620),
    .A2(net1724),
    .A1(net1625));
 sg13g2_nor3_1 _08303_ (.A(_02359_),
    .B(_02361_),
    .C(_02362_),
    .Y(_02363_));
 sg13g2_o21ai_1 _08304_ (.B1(_02359_),
    .Y(_02364_),
    .A1(_02361_),
    .A2(_02362_));
 sg13g2_nor2b_1 _08305_ (.A(_02363_),
    .B_N(_02364_),
    .Y(_02365_));
 sg13g2_o21ai_1 _08306_ (.B1(_02171_),
    .Y(_02366_),
    .A1(_02169_),
    .A2(_02172_));
 sg13g2_nand2_1 _08307_ (.Y(_02367_),
    .A(net1630),
    .B(net1718));
 sg13g2_and4_1 _08308_ (.A(net1640),
    .B(net1650),
    .C(net1706),
    .D(net1712),
    .X(_02368_));
 sg13g2_nand4_1 _08309_ (.B(net1650),
    .C(net1706),
    .A(net1640),
    .Y(_02369_),
    .D(net1712));
 sg13g2_a22oi_1 _08310_ (.Y(_02370_),
    .B1(net1712),
    .B2(net1640),
    .A2(net1706),
    .A1(net1650));
 sg13g2_or3_1 _08311_ (.A(_02367_),
    .B(_02368_),
    .C(_02370_),
    .X(_02371_));
 sg13g2_o21ai_1 _08312_ (.B1(_02367_),
    .Y(_02372_),
    .A1(_02368_),
    .A2(_02370_));
 sg13g2_and3_1 _08313_ (.X(_02373_),
    .A(_02366_),
    .B(_02371_),
    .C(_02372_));
 sg13g2_nand3_1 _08314_ (.B(_02371_),
    .C(_02372_),
    .A(_02366_),
    .Y(_02374_));
 sg13g2_a21o_1 _08315_ (.A2(_02372_),
    .A1(_02371_),
    .B1(_02366_),
    .X(_02375_));
 sg13g2_nand3_1 _08316_ (.B(_02374_),
    .C(_02375_),
    .A(_02365_),
    .Y(_02376_));
 sg13g2_a21o_1 _08317_ (.A2(_02375_),
    .A1(_02374_),
    .B1(_02365_),
    .X(_02377_));
 sg13g2_and3_1 _08318_ (.X(_02378_),
    .A(_02358_),
    .B(_02376_),
    .C(_02377_));
 sg13g2_nand3_1 _08319_ (.B(_02376_),
    .C(_02377_),
    .A(_02358_),
    .Y(_02379_));
 sg13g2_a21oi_1 _08320_ (.A1(_02376_),
    .A2(_02377_),
    .Y(_02380_),
    .B1(_02358_));
 sg13g2_or3_1 _08321_ (.A(_02357_),
    .B(_02378_),
    .C(_02380_),
    .X(_02381_));
 sg13g2_o21ai_1 _08322_ (.B1(_02357_),
    .Y(_02382_),
    .A1(_02378_),
    .A2(_02380_));
 sg13g2_and3_1 _08323_ (.X(_02383_),
    .A(_02345_),
    .B(_02381_),
    .C(_02382_));
 sg13g2_nand3_1 _08324_ (.B(_02381_),
    .C(_02382_),
    .A(_02345_),
    .Y(_02384_));
 sg13g2_a21o_1 _08325_ (.A2(_02382_),
    .A1(_02381_),
    .B1(_02345_),
    .X(_02385_));
 sg13g2_nand3_1 _08326_ (.B(_02384_),
    .C(_02385_),
    .A(_02344_),
    .Y(_02386_));
 sg13g2_a21o_1 _08327_ (.A2(_02385_),
    .A1(_02384_),
    .B1(_02344_),
    .X(_02387_));
 sg13g2_and3_1 _08328_ (.X(_02388_),
    .A(_02327_),
    .B(_02386_),
    .C(_02387_));
 sg13g2_a21oi_1 _08329_ (.A1(_02386_),
    .A2(_02387_),
    .Y(_02389_),
    .B1(_02327_));
 sg13g2_o21ai_1 _08330_ (.B1(_02164_),
    .Y(_02390_),
    .A1(_02388_),
    .A2(_02389_));
 sg13g2_or3_1 _08331_ (.A(_02164_),
    .B(_02388_),
    .C(_02389_),
    .X(_02391_));
 sg13g2_o21ai_1 _08332_ (.B1(_02208_),
    .Y(_02392_),
    .A1(_02071_),
    .A2(_02209_));
 sg13g2_nand3_1 _08333_ (.B(_02391_),
    .C(_02392_),
    .A(_02390_),
    .Y(_02393_));
 sg13g2_inv_1 _08334_ (.Y(_02394_),
    .A(_02393_));
 sg13g2_a21o_1 _08335_ (.A2(_02391_),
    .A1(_02390_),
    .B1(_02392_),
    .X(_02395_));
 sg13g2_nand2_1 _08336_ (.Y(_02396_),
    .A(_02393_),
    .B(_02395_));
 sg13g2_o21ai_1 _08337_ (.B1(_02258_),
    .Y(_02397_),
    .A1(_02259_),
    .A2(_02326_));
 sg13g2_nor4_2 _08338_ (.A(_02257_),
    .B(_02259_),
    .C(_02326_),
    .Y(_02398_),
    .D(_02396_));
 sg13g2_nand3_1 _08339_ (.B(_02393_),
    .C(_02395_),
    .A(_02257_),
    .Y(_02399_));
 sg13g2_xnor2_1 _08340_ (.Y(_02400_),
    .A(_02396_),
    .B(_02397_));
 sg13g2_and2_1 _08341_ (.A(_02325_),
    .B(_02400_),
    .X(_02401_));
 sg13g2_or2_1 _08342_ (.X(_02402_),
    .B(_02400_),
    .A(_02325_));
 sg13g2_nand2b_1 _08343_ (.Y(_02403_),
    .B(_02402_),
    .A_N(_02401_));
 sg13g2_o21ai_1 _08344_ (.B1(_02326_),
    .Y(_02404_),
    .A1(_02257_),
    .A2(_02259_));
 sg13g2_nand2_1 _08345_ (.Y(_02405_),
    .A(_02310_),
    .B(_02317_));
 sg13g2_nor2_1 _08346_ (.A(_02296_),
    .B(_02311_),
    .Y(_02406_));
 sg13g2_xnor2_1 _08347_ (.Y(_02407_),
    .A(_02281_),
    .B(_02282_));
 sg13g2_nand2_1 _08348_ (.Y(_02408_),
    .A(net1645),
    .B(net1546));
 sg13g2_nand2_1 _08349_ (.Y(_02409_),
    .A(net1634),
    .B(net1546));
 sg13g2_or2_1 _08350_ (.X(_02410_),
    .B(_02409_),
    .A(_02262_));
 sg13g2_nand2_1 _08351_ (.Y(_02411_),
    .A(net1629),
    .B(net1554));
 sg13g2_xnor2_1 _08352_ (.Y(_02412_),
    .A(_02262_),
    .B(_02409_));
 sg13g2_o21ai_1 _08353_ (.B1(_02410_),
    .Y(_02413_),
    .A1(_02411_),
    .A2(_02412_));
 sg13g2_o21ai_1 _08354_ (.B1(_02264_),
    .Y(_02414_),
    .A1(_02263_),
    .A2(_02265_));
 sg13g2_nor2b_1 _08355_ (.A(_02266_),
    .B_N(_02414_),
    .Y(_02415_));
 sg13g2_a22oi_1 _08356_ (.Y(_02416_),
    .B1(net1557),
    .B2(net1616),
    .A2(net1554),
    .A1(net1627));
 sg13g2_and2_1 _08357_ (.A(net1627),
    .B(net1557),
    .X(_02417_));
 sg13g2_nor2b_2 _08358_ (.A(_02278_),
    .B_N(_02417_),
    .Y(_02418_));
 sg13g2_xnor2_1 _08359_ (.Y(_02419_),
    .A(_02413_),
    .B(_02415_));
 sg13g2_nor3_1 _08360_ (.A(_02416_),
    .B(_02418_),
    .C(_02419_),
    .Y(_02420_));
 sg13g2_a21o_1 _08361_ (.A2(_02415_),
    .A1(_02413_),
    .B1(_02420_),
    .X(_02421_));
 sg13g2_nand2b_1 _08362_ (.Y(_02422_),
    .B(_02421_),
    .A_N(_02407_));
 sg13g2_xnor2_1 _08363_ (.Y(_02423_),
    .A(_02407_),
    .B(_02421_));
 sg13g2_nand2_1 _08364_ (.Y(_02424_),
    .A(_02418_),
    .B(_02423_));
 sg13g2_xnor2_1 _08365_ (.Y(_02425_),
    .A(_02297_),
    .B(_02298_));
 sg13g2_a21oi_1 _08366_ (.A1(_02422_),
    .A2(_02424_),
    .Y(_02426_),
    .B1(_02425_));
 sg13g2_xor2_1 _08367_ (.B(_02412_),
    .A(_02411_),
    .X(_02427_));
 sg13g2_o21ai_1 _08368_ (.B1(_02419_),
    .Y(_02428_),
    .A1(_02416_),
    .A2(_02418_));
 sg13g2_nor2b_1 _08369_ (.A(_02420_),
    .B_N(_02428_),
    .Y(_02429_));
 sg13g2_nand2_1 _08370_ (.Y(_02430_),
    .A(net1634),
    .B(net1554));
 sg13g2_nand2_1 _08371_ (.Y(_02431_),
    .A(net1628),
    .B(net1557));
 sg13g2_or2_1 _08372_ (.X(_02432_),
    .B(_02431_),
    .A(_02408_));
 sg13g2_o21ai_1 _08373_ (.B1(net1557),
    .Y(_02433_),
    .A1(net1628),
    .A2(net1645));
 sg13g2_a22oi_1 _08374_ (.Y(_02434_),
    .B1(_02433_),
    .B2(_02408_),
    .A2(_02432_),
    .A1(_02430_));
 sg13g2_a22oi_1 _08375_ (.Y(_02435_),
    .B1(_02429_),
    .B2(_02434_),
    .A2(_02427_),
    .A1(_02417_));
 sg13g2_o21ai_1 _08376_ (.B1(_02429_),
    .Y(_02436_),
    .A1(_02417_),
    .A2(_02427_));
 sg13g2_or4_1 _08377_ (.A(_05559_),
    .B(_05573_),
    .C(_02430_),
    .D(_02431_),
    .X(_02437_));
 sg13g2_a221oi_1 _08378_ (.B2(_02437_),
    .C1(_02435_),
    .B1(_02436_),
    .A1(_02418_),
    .Y(_02438_),
    .A2(_02423_));
 sg13g2_o21ai_1 _08379_ (.B1(_02438_),
    .Y(_02439_),
    .A1(_02418_),
    .A2(_02423_));
 sg13g2_a21oi_1 _08380_ (.A1(_02422_),
    .A2(_02425_),
    .Y(_02440_),
    .B1(_02439_));
 sg13g2_o21ai_1 _08381_ (.B1(_02312_),
    .Y(_02441_),
    .A1(_02426_),
    .A2(_02440_));
 sg13g2_nand2_1 _08382_ (.Y(_02442_),
    .A(_02318_),
    .B(_02405_));
 sg13g2_nor4_1 _08383_ (.A(_02322_),
    .B(_02406_),
    .C(_02441_),
    .D(_02442_),
    .Y(_02443_));
 sg13g2_or2_1 _08384_ (.X(_02444_),
    .B(_02321_),
    .A(_02261_));
 sg13g2_a21o_1 _08385_ (.A2(_02444_),
    .A1(_02326_),
    .B1(_02323_),
    .X(_02445_));
 sg13g2_and3_2 _08386_ (.X(_02446_),
    .A(_02404_),
    .B(_02443_),
    .C(_02445_));
 sg13g2_xnor2_1 _08387_ (.Y(_02447_),
    .A(_02403_),
    .B(_02446_));
 sg13g2_o21ai_1 _08388_ (.B1(net1760),
    .Y(_02448_),
    .A1(net1400),
    .A2(_02447_));
 sg13g2_a21oi_1 _08389_ (.A1(net1400),
    .A2(_05551_),
    .Y(_00312_),
    .B1(_02448_));
 sg13g2_a21o_1 _08390_ (.A2(_02446_),
    .A1(_02402_),
    .B1(_02401_),
    .X(_02449_));
 sg13g2_o21ai_1 _08391_ (.B1(_02342_),
    .Y(_02450_),
    .A1(_02162_),
    .A2(_02343_));
 sg13g2_a21o_1 _08392_ (.A2(_02385_),
    .A1(_02344_),
    .B1(_02383_),
    .X(_02451_));
 sg13g2_o21ai_1 _08393_ (.B1(_02379_),
    .Y(_02452_),
    .A1(_02357_),
    .A2(_02380_));
 sg13g2_o21ai_1 _08394_ (.B1(_02352_),
    .Y(_02453_),
    .A1(_02349_),
    .A2(_02353_));
 sg13g2_inv_1 _08395_ (.Y(_02454_),
    .A(_02453_));
 sg13g2_or2_1 _08396_ (.X(_02455_),
    .B(_02363_),
    .A(_02361_));
 sg13g2_nand2_1 _08397_ (.Y(_02456_),
    .A(net1599),
    .B(net1528));
 sg13g2_nand2_1 _08398_ (.Y(_02457_),
    .A(net1604),
    .B(net1516));
 sg13g2_nand2_1 _08399_ (.Y(_02458_),
    .A(net1609),
    .B(net1516));
 sg13g2_or2_1 _08400_ (.X(_02459_),
    .B(_02457_),
    .A(_02351_));
 sg13g2_xnor2_1 _08401_ (.Y(_02460_),
    .A(_02350_),
    .B(_02458_));
 sg13g2_xor2_1 _08402_ (.B(_02460_),
    .A(_02456_),
    .X(_02461_));
 sg13g2_nand2_1 _08403_ (.Y(_02462_),
    .A(_02455_),
    .B(_02461_));
 sg13g2_xnor2_1 _08404_ (.Y(_02463_),
    .A(_02455_),
    .B(_02461_));
 sg13g2_xnor2_1 _08405_ (.Y(_02464_),
    .A(_02454_),
    .B(_02463_));
 sg13g2_a21o_1 _08406_ (.A2(_02375_),
    .A1(_02365_),
    .B1(_02373_),
    .X(_02465_));
 sg13g2_nand2_1 _08407_ (.Y(_02466_),
    .A(net1613),
    .B(net1730));
 sg13g2_nand2_1 _08408_ (.Y(_02467_),
    .A(net1625),
    .B(net1717));
 sg13g2_or2_1 _08409_ (.X(_02468_),
    .B(_02467_),
    .A(_02360_));
 sg13g2_and2_1 _08410_ (.A(_02360_),
    .B(_02467_),
    .X(_02469_));
 sg13g2_xnor2_1 _08411_ (.Y(_02470_),
    .A(_02360_),
    .B(_02467_));
 sg13g2_xnor2_1 _08412_ (.Y(_02471_),
    .A(_02466_),
    .B(_02470_));
 sg13g2_o21ai_1 _08413_ (.B1(_02369_),
    .Y(_02472_),
    .A1(_02367_),
    .A2(_02370_));
 sg13g2_nand2_1 _08414_ (.Y(_02473_),
    .A(net1630),
    .B(net1712));
 sg13g2_and4_1 _08415_ (.A(net1641),
    .B(net1650),
    .C(net1699),
    .D(net1706),
    .X(_02474_));
 sg13g2_nand4_1 _08416_ (.B(net1651),
    .C(net1699),
    .A(net1640),
    .Y(_02475_),
    .D(net1706));
 sg13g2_a22oi_1 _08417_ (.Y(_02476_),
    .B1(net1706),
    .B2(net1640),
    .A2(net1699),
    .A1(net1651));
 sg13g2_or3_1 _08418_ (.A(_02473_),
    .B(_02474_),
    .C(_02476_),
    .X(_02477_));
 sg13g2_o21ai_1 _08419_ (.B1(_02473_),
    .Y(_02478_),
    .A1(_02474_),
    .A2(_02476_));
 sg13g2_and3_1 _08420_ (.X(_02479_),
    .A(_02472_),
    .B(_02477_),
    .C(_02478_));
 sg13g2_nand3_1 _08421_ (.B(_02477_),
    .C(_02478_),
    .A(_02472_),
    .Y(_02480_));
 sg13g2_a21oi_1 _08422_ (.A1(_02477_),
    .A2(_02478_),
    .Y(_02481_),
    .B1(_02472_));
 sg13g2_or3_1 _08423_ (.A(_02471_),
    .B(_02479_),
    .C(_02481_),
    .X(_02482_));
 sg13g2_o21ai_1 _08424_ (.B1(_02471_),
    .Y(_02483_),
    .A1(_02479_),
    .A2(_02481_));
 sg13g2_and3_1 _08425_ (.X(_02484_),
    .A(_02465_),
    .B(_02482_),
    .C(_02483_));
 sg13g2_nand3_1 _08426_ (.B(_02482_),
    .C(_02483_),
    .A(_02465_),
    .Y(_02485_));
 sg13g2_a21oi_1 _08427_ (.A1(_02482_),
    .A2(_02483_),
    .Y(_02486_),
    .B1(_02465_));
 sg13g2_or3_1 _08428_ (.A(_02464_),
    .B(_02484_),
    .C(_02486_),
    .X(_02487_));
 sg13g2_o21ai_1 _08429_ (.B1(_02464_),
    .Y(_02488_),
    .A1(_02484_),
    .A2(_02486_));
 sg13g2_and3_1 _08430_ (.X(_02489_),
    .A(_02452_),
    .B(_02487_),
    .C(_02488_));
 sg13g2_nand3_1 _08431_ (.B(_02487_),
    .C(_02488_),
    .A(_02452_),
    .Y(_02490_));
 sg13g2_a21oi_1 _08432_ (.A1(_02487_),
    .A2(_02488_),
    .Y(_02491_),
    .B1(_02452_));
 sg13g2_nand2_1 _08433_ (.Y(_02492_),
    .A(_02338_),
    .B(_02340_));
 sg13g2_o21ai_1 _08434_ (.B1(_02355_),
    .Y(_02493_),
    .A1(_02347_),
    .A2(_02356_));
 sg13g2_inv_1 _08435_ (.Y(_02494_),
    .A(_02493_));
 sg13g2_a22oi_1 _08436_ (.Y(_02495_),
    .B1(net1555),
    .B2(net1571),
    .A2(net1551),
    .A1(net1577));
 sg13g2_nand2_1 _08437_ (.Y(_02496_),
    .A(net1571),
    .B(net1552));
 sg13g2_or2_1 _08438_ (.X(_02497_),
    .B(_02496_),
    .A(_02329_));
 sg13g2_nand2b_1 _08439_ (.Y(_02498_),
    .B(_02497_),
    .A_N(_02495_));
 sg13g2_or2_1 _08440_ (.X(_02499_),
    .B(_02335_),
    .A(_02333_));
 sg13g2_nand2_1 _08441_ (.Y(_02500_),
    .A(net1581),
    .B(net1545));
 sg13g2_nand2_1 _08442_ (.Y(_02501_),
    .A(net1594),
    .B(net1533));
 sg13g2_or2_1 _08443_ (.X(_02502_),
    .B(_02501_),
    .A(_02332_));
 sg13g2_and2_1 _08444_ (.A(_02332_),
    .B(_02501_),
    .X(_02503_));
 sg13g2_xor2_1 _08445_ (.B(_02501_),
    .A(_02332_),
    .X(_02504_));
 sg13g2_xnor2_1 _08446_ (.Y(_02505_),
    .A(_02500_),
    .B(_02504_));
 sg13g2_nand2_1 _08447_ (.Y(_02506_),
    .A(_02499_),
    .B(_02505_));
 sg13g2_xnor2_1 _08448_ (.Y(_02507_),
    .A(_02499_),
    .B(_02505_));
 sg13g2_xnor2_1 _08449_ (.Y(_02508_),
    .A(_02498_),
    .B(_02507_));
 sg13g2_xor2_1 _08450_ (.B(_02508_),
    .A(_02493_),
    .X(_02509_));
 sg13g2_nand2b_1 _08451_ (.Y(_02510_),
    .B(_02492_),
    .A_N(_02509_));
 sg13g2_xor2_1 _08452_ (.B(_02509_),
    .A(_02492_),
    .X(_02511_));
 sg13g2_or3_1 _08453_ (.A(_02489_),
    .B(_02491_),
    .C(_02511_),
    .X(_02512_));
 sg13g2_o21ai_1 _08454_ (.B1(_02511_),
    .Y(_02513_),
    .A1(_02489_),
    .A2(_02491_));
 sg13g2_and3_1 _08455_ (.X(_02514_),
    .A(_02451_),
    .B(_02512_),
    .C(_02513_));
 sg13g2_a21o_1 _08456_ (.A2(_02513_),
    .A1(_02512_),
    .B1(_02451_),
    .X(_02515_));
 sg13g2_nand2b_1 _08457_ (.Y(_02516_),
    .B(_02515_),
    .A_N(_02514_));
 sg13g2_xnor2_1 _08458_ (.Y(_02517_),
    .A(_02450_),
    .B(_02516_));
 sg13g2_nand2b_2 _08459_ (.Y(_02518_),
    .B(_02391_),
    .A_N(_02388_));
 sg13g2_nand2_2 _08460_ (.Y(_02519_),
    .A(_02517_),
    .B(_02518_));
 sg13g2_or2_1 _08461_ (.X(_02520_),
    .B(_02518_),
    .A(_02517_));
 sg13g2_xor2_1 _08462_ (.B(_02518_),
    .A(_02517_),
    .X(_02521_));
 sg13g2_nand2_1 _08463_ (.Y(_02522_),
    .A(_02394_),
    .B(_02521_));
 sg13g2_xnor2_1 _08464_ (.Y(_02523_),
    .A(_02394_),
    .B(_02521_));
 sg13g2_xor2_1 _08465_ (.B(_02523_),
    .A(_02399_),
    .X(_02524_));
 sg13g2_nor2_1 _08466_ (.A(_02398_),
    .B(_02524_),
    .Y(_02525_));
 sg13g2_xor2_1 _08467_ (.B(_02524_),
    .A(_02398_),
    .X(_02526_));
 sg13g2_xnor2_1 _08468_ (.Y(_02527_),
    .A(_02449_),
    .B(_02526_));
 sg13g2_o21ai_1 _08469_ (.B1(net1760),
    .Y(_02528_),
    .A1(net1473),
    .A2(net615));
 sg13g2_a21oi_1 _08470_ (.A1(net1472),
    .A2(_02527_),
    .Y(_00313_),
    .B1(net616));
 sg13g2_a221oi_1 _08471_ (.B2(_02398_),
    .C1(_02401_),
    .B1(_02524_),
    .A1(_02402_),
    .Y(_02529_),
    .A2(_02446_));
 sg13g2_o21ai_1 _08472_ (.B1(_02510_),
    .Y(_02530_),
    .A1(_02494_),
    .A2(_02508_));
 sg13g2_nand2b_1 _08473_ (.Y(_02531_),
    .B(_02530_),
    .A_N(_02497_));
 sg13g2_xnor2_1 _08474_ (.Y(_02532_),
    .A(_02497_),
    .B(_02530_));
 sg13g2_o21ai_1 _08475_ (.B1(_02490_),
    .Y(_02533_),
    .A1(_02491_),
    .A2(_02511_));
 sg13g2_o21ai_1 _08476_ (.B1(_02506_),
    .Y(_02534_),
    .A1(_02498_),
    .A2(_02507_));
 sg13g2_inv_1 _08477_ (.Y(_02535_),
    .A(_02534_));
 sg13g2_o21ai_1 _08478_ (.B1(_02462_),
    .Y(_02536_),
    .A1(_02454_),
    .A2(_02463_));
 sg13g2_nand2_1 _08479_ (.Y(_02537_),
    .A(net1567),
    .B(net1555));
 sg13g2_nand2_1 _08480_ (.Y(_02538_),
    .A(net1571),
    .B(net1545));
 sg13g2_nand2_1 _08481_ (.Y(_02539_),
    .A(net1577),
    .B(net1545));
 sg13g2_xor2_1 _08482_ (.B(_02539_),
    .A(_02496_),
    .X(_02540_));
 sg13g2_nand2b_1 _08483_ (.Y(_02541_),
    .B(_02540_),
    .A_N(_02537_));
 sg13g2_xnor2_1 _08484_ (.Y(_02542_),
    .A(_02537_),
    .B(_02540_));
 sg13g2_inv_1 _08485_ (.Y(_02543_),
    .A(_02542_));
 sg13g2_o21ai_1 _08486_ (.B1(_02502_),
    .Y(_02544_),
    .A1(_02500_),
    .A2(_02503_));
 sg13g2_nand2_1 _08487_ (.Y(_02545_),
    .A(net1581),
    .B(net1538));
 sg13g2_nand2_1 _08488_ (.Y(_02546_),
    .A(net1588),
    .B(net1528));
 sg13g2_and4_1 _08489_ (.A(net1587),
    .B(net1594),
    .C(net1529),
    .D(net1534),
    .X(_02547_));
 sg13g2_a22oi_1 _08490_ (.Y(_02548_),
    .B1(net1534),
    .B2(net1588),
    .A2(net1529),
    .A1(net1595));
 sg13g2_nor3_1 _08491_ (.A(_02545_),
    .B(_02547_),
    .C(_02548_),
    .Y(_02549_));
 sg13g2_o21ai_1 _08492_ (.B1(_02545_),
    .Y(_02550_),
    .A1(_02547_),
    .A2(_02548_));
 sg13g2_nor2b_1 _08493_ (.A(_02549_),
    .B_N(_02550_),
    .Y(_02551_));
 sg13g2_nand2_1 _08494_ (.Y(_02552_),
    .A(_02544_),
    .B(_02551_));
 sg13g2_xnor2_1 _08495_ (.Y(_02553_),
    .A(_02544_),
    .B(_02551_));
 sg13g2_xnor2_1 _08496_ (.Y(_02554_),
    .A(_02543_),
    .B(_02553_));
 sg13g2_nand2b_1 _08497_ (.Y(_02555_),
    .B(_02536_),
    .A_N(_02554_));
 sg13g2_xor2_1 _08498_ (.B(_02554_),
    .A(_02536_),
    .X(_02556_));
 sg13g2_xnor2_1 _08499_ (.Y(_02557_),
    .A(_02535_),
    .B(_02556_));
 sg13g2_o21ai_1 _08500_ (.B1(_02485_),
    .Y(_02558_),
    .A1(_02464_),
    .A2(_02486_));
 sg13g2_o21ai_1 _08501_ (.B1(_02459_),
    .Y(_02559_),
    .A1(_02456_),
    .A2(_02460_));
 sg13g2_inv_1 _08502_ (.Y(_02560_),
    .A(_02559_));
 sg13g2_o21ai_1 _08503_ (.B1(_02468_),
    .Y(_02561_),
    .A1(_02466_),
    .A2(_02469_));
 sg13g2_nand2_1 _08504_ (.Y(_02562_),
    .A(net1599),
    .B(net1522));
 sg13g2_nand2_1 _08505_ (.Y(_02563_),
    .A(net1604),
    .B(net1730));
 sg13g2_nand2_1 _08506_ (.Y(_02564_),
    .A(net1609),
    .B(net1730));
 sg13g2_or2_1 _08507_ (.X(_02565_),
    .B(_02563_),
    .A(_02458_));
 sg13g2_xnor2_1 _08508_ (.Y(_02566_),
    .A(_02457_),
    .B(_02564_));
 sg13g2_xor2_1 _08509_ (.B(_02566_),
    .A(_02562_),
    .X(_02567_));
 sg13g2_nand2_1 _08510_ (.Y(_02568_),
    .A(_02561_),
    .B(_02567_));
 sg13g2_xnor2_1 _08511_ (.Y(_02569_),
    .A(_02561_),
    .B(_02567_));
 sg13g2_xnor2_1 _08512_ (.Y(_02570_),
    .A(_02560_),
    .B(_02569_));
 sg13g2_o21ai_1 _08513_ (.B1(_02480_),
    .Y(_02571_),
    .A1(_02471_),
    .A2(_02481_));
 sg13g2_nand2_1 _08514_ (.Y(_02572_),
    .A(net1613),
    .B(net1723));
 sg13g2_nand2_1 _08515_ (.Y(_02573_),
    .A(net1620),
    .B(net1713));
 sg13g2_and4_1 _08516_ (.A(net1620),
    .B(net1625),
    .C(net1712),
    .D(net1717),
    .X(_02574_));
 sg13g2_a22oi_1 _08517_ (.Y(_02575_),
    .B1(net1717),
    .B2(net1620),
    .A2(net1713),
    .A1(net1626));
 sg13g2_nor3_1 _08518_ (.A(_02572_),
    .B(_02574_),
    .C(_02575_),
    .Y(_02576_));
 sg13g2_o21ai_1 _08519_ (.B1(_02572_),
    .Y(_02577_),
    .A1(_02574_),
    .A2(_02575_));
 sg13g2_nand2b_1 _08520_ (.Y(_02578_),
    .B(_02577_),
    .A_N(_02576_));
 sg13g2_o21ai_1 _08521_ (.B1(_02475_),
    .Y(_02579_),
    .A1(_02473_),
    .A2(_02476_));
 sg13g2_nand2_1 _08522_ (.Y(_02580_),
    .A(net1630),
    .B(net1707));
 sg13g2_and4_1 _08523_ (.A(net1640),
    .B(net1650),
    .C(net1694),
    .D(net1699),
    .X(_02581_));
 sg13g2_nand4_1 _08524_ (.B(net1650),
    .C(net1694),
    .A(net1640),
    .Y(_02582_),
    .D(net1699));
 sg13g2_a22oi_1 _08525_ (.Y(_02583_),
    .B1(net1700),
    .B2(net1640),
    .A2(net1694),
    .A1(net1650));
 sg13g2_or3_1 _08526_ (.A(_02580_),
    .B(_02581_),
    .C(_02583_),
    .X(_02584_));
 sg13g2_o21ai_1 _08527_ (.B1(_02580_),
    .Y(_02585_),
    .A1(_02581_),
    .A2(_02583_));
 sg13g2_and3_1 _08528_ (.X(_02586_),
    .A(_02579_),
    .B(_02584_),
    .C(_02585_));
 sg13g2_nand3_1 _08529_ (.B(_02584_),
    .C(_02585_),
    .A(_02579_),
    .Y(_02587_));
 sg13g2_a21oi_1 _08530_ (.A1(_02584_),
    .A2(_02585_),
    .Y(_02588_),
    .B1(_02579_));
 sg13g2_or3_1 _08531_ (.A(_02578_),
    .B(_02586_),
    .C(_02588_),
    .X(_02589_));
 sg13g2_o21ai_1 _08532_ (.B1(_02578_),
    .Y(_02590_),
    .A1(_02586_),
    .A2(_02588_));
 sg13g2_and3_1 _08533_ (.X(_02591_),
    .A(_02571_),
    .B(_02589_),
    .C(_02590_));
 sg13g2_nand3_1 _08534_ (.B(_02589_),
    .C(_02590_),
    .A(_02571_),
    .Y(_02592_));
 sg13g2_a21oi_1 _08535_ (.A1(_02589_),
    .A2(_02590_),
    .Y(_02593_),
    .B1(_02571_));
 sg13g2_or3_1 _08536_ (.A(_02570_),
    .B(_02591_),
    .C(_02593_),
    .X(_02594_));
 sg13g2_o21ai_1 _08537_ (.B1(_02570_),
    .Y(_02595_),
    .A1(_02591_),
    .A2(_02593_));
 sg13g2_and3_1 _08538_ (.X(_02596_),
    .A(_02558_),
    .B(_02594_),
    .C(_02595_));
 sg13g2_nand3_1 _08539_ (.B(_02594_),
    .C(_02595_),
    .A(_02558_),
    .Y(_02597_));
 sg13g2_a21oi_1 _08540_ (.A1(_02594_),
    .A2(_02595_),
    .Y(_02598_),
    .B1(_02558_));
 sg13g2_or3_1 _08541_ (.A(_02557_),
    .B(_02596_),
    .C(_02598_),
    .X(_02599_));
 sg13g2_o21ai_1 _08542_ (.B1(_02557_),
    .Y(_02600_),
    .A1(_02596_),
    .A2(_02598_));
 sg13g2_and3_1 _08543_ (.X(_02601_),
    .A(_02533_),
    .B(_02599_),
    .C(_02600_));
 sg13g2_nand3_1 _08544_ (.B(_02599_),
    .C(_02600_),
    .A(_02533_),
    .Y(_02602_));
 sg13g2_a21o_1 _08545_ (.A2(_02600_),
    .A1(_02599_),
    .B1(_02533_),
    .X(_02603_));
 sg13g2_a21oi_1 _08546_ (.A1(_02602_),
    .A2(_02603_),
    .Y(_02604_),
    .B1(_02532_));
 sg13g2_and3_1 _08547_ (.X(_02605_),
    .A(_02532_),
    .B(_02602_),
    .C(_02603_));
 sg13g2_a21oi_1 _08548_ (.A1(_02450_),
    .A2(_02515_),
    .Y(_02606_),
    .B1(_02514_));
 sg13g2_or3_1 _08549_ (.A(_02604_),
    .B(_02605_),
    .C(_02606_),
    .X(_02607_));
 sg13g2_o21ai_1 _08550_ (.B1(_02606_),
    .Y(_02608_),
    .A1(_02604_),
    .A2(_02605_));
 sg13g2_and2_1 _08551_ (.A(_02607_),
    .B(_02608_),
    .X(_02609_));
 sg13g2_nor2b_2 _08552_ (.A(_02519_),
    .B_N(_02609_),
    .Y(_02610_));
 sg13g2_xor2_1 _08553_ (.B(_02609_),
    .A(_02519_),
    .X(_02611_));
 sg13g2_o21ai_1 _08554_ (.B1(_02522_),
    .Y(_02612_),
    .A1(_02399_),
    .A2(_02523_));
 sg13g2_and4_1 _08555_ (.A(_02394_),
    .B(_02519_),
    .C(_02520_),
    .D(_02609_),
    .X(_02613_));
 sg13g2_nor3_1 _08556_ (.A(_02399_),
    .B(_02523_),
    .C(_02611_),
    .Y(_02614_));
 sg13g2_inv_1 _08557_ (.Y(_02615_),
    .A(_02614_));
 sg13g2_xor2_1 _08558_ (.B(_02612_),
    .A(_02611_),
    .X(_02616_));
 sg13g2_nor3_1 _08559_ (.A(_02525_),
    .B(_02529_),
    .C(_02616_),
    .Y(_02617_));
 sg13g2_o21ai_1 _08560_ (.B1(_02616_),
    .Y(_02618_),
    .A1(_02525_),
    .A2(_02529_));
 sg13g2_nor2b_2 _08561_ (.A(_02617_),
    .B_N(_02618_),
    .Y(_02619_));
 sg13g2_o21ai_1 _08562_ (.B1(net1758),
    .Y(_02620_),
    .A1(net1399),
    .A2(_02619_));
 sg13g2_a21oi_1 _08563_ (.A1(net1399),
    .A2(_05550_),
    .Y(_00314_),
    .B1(_02620_));
 sg13g2_a21o_1 _08564_ (.A2(_02603_),
    .A1(_02532_),
    .B1(_02601_),
    .X(_02621_));
 sg13g2_o21ai_1 _08565_ (.B1(_02555_),
    .Y(_02622_),
    .A1(_02535_),
    .A2(_02556_));
 sg13g2_o21ai_1 _08566_ (.B1(_02541_),
    .Y(_02623_),
    .A1(_02496_),
    .A2(_02539_));
 sg13g2_nand2_2 _08567_ (.Y(_02624_),
    .A(net1563),
    .B(net1555));
 sg13g2_nand2b_1 _08568_ (.Y(_02625_),
    .B(_02623_),
    .A_N(_02624_));
 sg13g2_xnor2_1 _08569_ (.Y(_02626_),
    .A(_02623_),
    .B(_02624_));
 sg13g2_nand2_1 _08570_ (.Y(_02627_),
    .A(_02622_),
    .B(_02626_));
 sg13g2_xnor2_1 _08571_ (.Y(_02628_),
    .A(_02622_),
    .B(_02626_));
 sg13g2_o21ai_1 _08572_ (.B1(_02597_),
    .Y(_02629_),
    .A1(_02557_),
    .A2(_02598_));
 sg13g2_o21ai_1 _08573_ (.B1(_02552_),
    .Y(_02630_),
    .A1(_02543_),
    .A2(_02553_));
 sg13g2_inv_1 _08574_ (.Y(_02631_),
    .A(_02630_));
 sg13g2_o21ai_1 _08575_ (.B1(_02568_),
    .Y(_02632_),
    .A1(_02560_),
    .A2(_02569_));
 sg13g2_nand2_2 _08576_ (.Y(_02633_),
    .A(net1575),
    .B(net1538));
 sg13g2_xor2_1 _08577_ (.B(_02633_),
    .A(_02538_),
    .X(_02634_));
 sg13g2_nand3_1 _08578_ (.B(net1551),
    .C(_02634_),
    .A(net1567),
    .Y(_02635_));
 sg13g2_a21o_1 _08579_ (.A2(net1551),
    .A1(net1567),
    .B1(_02634_),
    .X(_02636_));
 sg13g2_nand2_1 _08580_ (.Y(_02637_),
    .A(_02635_),
    .B(_02636_));
 sg13g2_or2_1 _08581_ (.X(_02638_),
    .B(_02549_),
    .A(_02547_));
 sg13g2_nand2_1 _08582_ (.Y(_02639_),
    .A(net1581),
    .B(net1534));
 sg13g2_nand2_1 _08583_ (.Y(_02640_),
    .A(net1594),
    .B(net1521));
 sg13g2_or2_1 _08584_ (.X(_02641_),
    .B(_02640_),
    .A(_02546_));
 sg13g2_and2_1 _08585_ (.A(_02546_),
    .B(_02640_),
    .X(_02642_));
 sg13g2_xor2_1 _08586_ (.B(_02640_),
    .A(_02546_),
    .X(_02643_));
 sg13g2_xnor2_1 _08587_ (.Y(_02644_),
    .A(_02639_),
    .B(_02643_));
 sg13g2_nand2_1 _08588_ (.Y(_02645_),
    .A(_02638_),
    .B(_02644_));
 sg13g2_xnor2_1 _08589_ (.Y(_02646_),
    .A(_02638_),
    .B(_02644_));
 sg13g2_xnor2_1 _08590_ (.Y(_02647_),
    .A(_02637_),
    .B(_02646_));
 sg13g2_nand2b_1 _08591_ (.Y(_02648_),
    .B(_02632_),
    .A_N(_02647_));
 sg13g2_xor2_1 _08592_ (.B(_02647_),
    .A(_02632_),
    .X(_02649_));
 sg13g2_xnor2_1 _08593_ (.Y(_02650_),
    .A(_02631_),
    .B(_02649_));
 sg13g2_o21ai_1 _08594_ (.B1(_02592_),
    .Y(_02651_),
    .A1(_02570_),
    .A2(_02593_));
 sg13g2_o21ai_1 _08595_ (.B1(_02565_),
    .Y(_02652_),
    .A1(_02562_),
    .A2(_02566_));
 sg13g2_inv_1 _08596_ (.Y(_02653_),
    .A(_02652_));
 sg13g2_or2_1 _08597_ (.X(_02654_),
    .B(_02576_),
    .A(_02574_));
 sg13g2_nand2_1 _08598_ (.Y(_02655_),
    .A(net1599),
    .B(net1517));
 sg13g2_nand2_1 _08599_ (.Y(_02656_),
    .A(net1604),
    .B(net1724));
 sg13g2_nand2_1 _08600_ (.Y(_02657_),
    .A(net1609),
    .B(net1724));
 sg13g2_or2_1 _08601_ (.X(_02658_),
    .B(_02656_),
    .A(_02564_));
 sg13g2_xnor2_1 _08602_ (.Y(_02659_),
    .A(_02563_),
    .B(_02657_));
 sg13g2_xor2_1 _08603_ (.B(_02659_),
    .A(_02655_),
    .X(_02660_));
 sg13g2_nand2_1 _08604_ (.Y(_02661_),
    .A(_02654_),
    .B(_02660_));
 sg13g2_xnor2_1 _08605_ (.Y(_02662_),
    .A(_02654_),
    .B(_02660_));
 sg13g2_xnor2_1 _08606_ (.Y(_02663_),
    .A(_02652_),
    .B(_02662_));
 sg13g2_xnor2_1 _08607_ (.Y(_02664_),
    .A(_02653_),
    .B(_02662_));
 sg13g2_o21ai_1 _08608_ (.B1(_02587_),
    .Y(_02665_),
    .A1(_02578_),
    .A2(_02588_));
 sg13g2_nand2_1 _08609_ (.Y(_02666_),
    .A(net1613),
    .B(net1717));
 sg13g2_nand2_1 _08610_ (.Y(_02667_),
    .A(net1625),
    .B(net1706));
 sg13g2_or2_1 _08611_ (.X(_02668_),
    .B(_02667_),
    .A(_02573_));
 sg13g2_and2_1 _08612_ (.A(_02573_),
    .B(_02667_),
    .X(_02669_));
 sg13g2_xor2_1 _08613_ (.B(_02667_),
    .A(_02573_),
    .X(_02670_));
 sg13g2_xnor2_1 _08614_ (.Y(_02671_),
    .A(_02666_),
    .B(_02670_));
 sg13g2_o21ai_1 _08615_ (.B1(_02582_),
    .Y(_02672_),
    .A1(_02580_),
    .A2(_02583_));
 sg13g2_nand2_1 _08616_ (.Y(_02673_),
    .A(net1630),
    .B(net1699));
 sg13g2_and4_1 _08617_ (.A(net1642),
    .B(net1652),
    .C(net1689),
    .D(net1694),
    .X(_02674_));
 sg13g2_nand4_1 _08618_ (.B(net1652),
    .C(net1689),
    .A(net1642),
    .Y(_02675_),
    .D(net1694));
 sg13g2_a22oi_1 _08619_ (.Y(_02676_),
    .B1(net1695),
    .B2(net1642),
    .A2(net1689),
    .A1(net1652));
 sg13g2_or3_1 _08620_ (.A(_02673_),
    .B(_02674_),
    .C(_02676_),
    .X(_02677_));
 sg13g2_o21ai_1 _08621_ (.B1(_02673_),
    .Y(_02678_),
    .A1(_02674_),
    .A2(_02676_));
 sg13g2_and3_1 _08622_ (.X(_02679_),
    .A(_02672_),
    .B(_02677_),
    .C(_02678_));
 sg13g2_nand3_1 _08623_ (.B(_02677_),
    .C(_02678_),
    .A(_02672_),
    .Y(_02680_));
 sg13g2_a21o_1 _08624_ (.A2(_02678_),
    .A1(_02677_),
    .B1(_02672_),
    .X(_02681_));
 sg13g2_nand3_1 _08625_ (.B(_02680_),
    .C(_02681_),
    .A(_02671_),
    .Y(_02682_));
 sg13g2_a21o_1 _08626_ (.A2(_02681_),
    .A1(_02680_),
    .B1(_02671_),
    .X(_02683_));
 sg13g2_nand3_1 _08627_ (.B(_02682_),
    .C(_02683_),
    .A(_02665_),
    .Y(_02684_));
 sg13g2_a21oi_1 _08628_ (.A1(_02682_),
    .A2(_02683_),
    .Y(_02685_),
    .B1(_02665_));
 sg13g2_a21o_1 _08629_ (.A2(_02683_),
    .A1(_02682_),
    .B1(_02665_),
    .X(_02686_));
 sg13g2_nand3_1 _08630_ (.B(_02684_),
    .C(_02686_),
    .A(_02663_),
    .Y(_02687_));
 sg13g2_a21o_1 _08631_ (.A2(_02686_),
    .A1(_02684_),
    .B1(_02663_),
    .X(_02688_));
 sg13g2_and3_1 _08632_ (.X(_02689_),
    .A(_02651_),
    .B(_02687_),
    .C(_02688_));
 sg13g2_nand3_1 _08633_ (.B(_02687_),
    .C(_02688_),
    .A(_02651_),
    .Y(_02690_));
 sg13g2_a21oi_1 _08634_ (.A1(_02687_),
    .A2(_02688_),
    .Y(_02691_),
    .B1(_02651_));
 sg13g2_or3_1 _08635_ (.A(_02650_),
    .B(_02689_),
    .C(_02691_),
    .X(_02692_));
 sg13g2_o21ai_1 _08636_ (.B1(_02650_),
    .Y(_02693_),
    .A1(_02689_),
    .A2(_02691_));
 sg13g2_and3_1 _08637_ (.X(_02694_),
    .A(_02629_),
    .B(_02692_),
    .C(_02693_));
 sg13g2_nand3_1 _08638_ (.B(_02692_),
    .C(_02693_),
    .A(_02629_),
    .Y(_02695_));
 sg13g2_a21oi_1 _08639_ (.A1(_02692_),
    .A2(_02693_),
    .Y(_02696_),
    .B1(_02629_));
 sg13g2_or3_1 _08640_ (.A(_02628_),
    .B(_02694_),
    .C(_02696_),
    .X(_02697_));
 sg13g2_o21ai_1 _08641_ (.B1(_02628_),
    .Y(_02698_),
    .A1(_02694_),
    .A2(_02696_));
 sg13g2_and3_1 _08642_ (.X(_02699_),
    .A(_02621_),
    .B(_02697_),
    .C(_02698_));
 sg13g2_nand3_1 _08643_ (.B(_02697_),
    .C(_02698_),
    .A(_02621_),
    .Y(_02700_));
 sg13g2_a21oi_1 _08644_ (.A1(_02697_),
    .A2(_02698_),
    .Y(_02701_),
    .B1(_02621_));
 sg13g2_o21ai_1 _08645_ (.B1(_02531_),
    .Y(_02702_),
    .A1(_02699_),
    .A2(_02701_));
 sg13g2_or3_1 _08646_ (.A(_02531_),
    .B(_02699_),
    .C(_02701_),
    .X(_02703_));
 sg13g2_nand2_1 _08647_ (.Y(_02704_),
    .A(_02702_),
    .B(_02703_));
 sg13g2_nand3b_1 _08648_ (.B(_02702_),
    .C(_02703_),
    .Y(_02705_),
    .A_N(_02607_));
 sg13g2_xor2_1 _08649_ (.B(_02704_),
    .A(_02607_),
    .X(_02706_));
 sg13g2_nor2_1 _08650_ (.A(_02610_),
    .B(_02613_),
    .Y(_02707_));
 sg13g2_xor2_1 _08651_ (.B(_02707_),
    .A(_02706_),
    .X(_02708_));
 sg13g2_nor2_1 _08652_ (.A(_02614_),
    .B(_02617_),
    .Y(_02709_));
 sg13g2_nor4_1 _08653_ (.A(_02525_),
    .B(_02529_),
    .C(_02616_),
    .D(_02708_),
    .Y(_02710_));
 sg13g2_xnor2_1 _08654_ (.Y(_02711_),
    .A(_02708_),
    .B(_02709_));
 sg13g2_o21ai_1 _08655_ (.B1(net1761),
    .Y(_02712_),
    .A1(net1469),
    .A2(net594));
 sg13g2_a21oi_1 _08656_ (.A1(net1469),
    .A2(_02711_),
    .Y(_00315_),
    .B1(_02712_));
 sg13g2_nand2_1 _08657_ (.Y(_02713_),
    .A(_02613_),
    .B(_02706_));
 sg13g2_o21ai_1 _08658_ (.B1(_02713_),
    .Y(_02714_),
    .A1(_02615_),
    .A2(_02708_));
 sg13g2_or2_1 _08659_ (.X(_02715_),
    .B(_02714_),
    .A(_02710_));
 sg13g2_o21ai_1 _08660_ (.B1(_02700_),
    .Y(_02716_),
    .A1(_02531_),
    .A2(_02701_));
 sg13g2_o21ai_1 _08661_ (.B1(_02695_),
    .Y(_02717_),
    .A1(_02628_),
    .A2(_02696_));
 sg13g2_o21ai_1 _08662_ (.B1(_02648_),
    .Y(_02718_),
    .A1(_02631_),
    .A2(_02649_));
 sg13g2_o21ai_1 _08663_ (.B1(_02635_),
    .Y(_02719_),
    .A1(_02538_),
    .A2(_02633_));
 sg13g2_a22oi_1 _08664_ (.Y(_02720_),
    .B1(net1556),
    .B2(net1511),
    .A2(net1551),
    .A1(net1563));
 sg13g2_nand2_2 _08665_ (.Y(_02721_),
    .A(net1511),
    .B(net1553));
 sg13g2_nor2_1 _08666_ (.A(_02624_),
    .B(_02721_),
    .Y(_02722_));
 sg13g2_or2_1 _08667_ (.X(_02723_),
    .B(_02721_),
    .A(_02624_));
 sg13g2_nor2_1 _08668_ (.A(_02720_),
    .B(_02722_),
    .Y(_02724_));
 sg13g2_and2_1 _08669_ (.A(_02719_),
    .B(_02724_),
    .X(_02725_));
 sg13g2_xnor2_1 _08670_ (.Y(_02726_),
    .A(_02719_),
    .B(_02724_));
 sg13g2_nor2_1 _08671_ (.A(_02625_),
    .B(_02726_),
    .Y(_02727_));
 sg13g2_inv_1 _08672_ (.Y(_02728_),
    .A(_02727_));
 sg13g2_xor2_1 _08673_ (.B(_02726_),
    .A(_02625_),
    .X(_02729_));
 sg13g2_nand2_1 _08674_ (.Y(_02730_),
    .A(_02718_),
    .B(_02729_));
 sg13g2_xnor2_1 _08675_ (.Y(_02731_),
    .A(_02718_),
    .B(_02729_));
 sg13g2_o21ai_1 _08676_ (.B1(_02690_),
    .Y(_02732_),
    .A1(_02650_),
    .A2(_02691_));
 sg13g2_o21ai_1 _08677_ (.B1(_02645_),
    .Y(_02733_),
    .A1(_02637_),
    .A2(_02646_));
 sg13g2_inv_1 _08678_ (.Y(_02734_),
    .A(_02733_));
 sg13g2_o21ai_1 _08679_ (.B1(_02661_),
    .Y(_02735_),
    .A1(_02653_),
    .A2(_02662_));
 sg13g2_nand2_1 _08680_ (.Y(_02736_),
    .A(net1567),
    .B(net1545));
 sg13g2_nand2_2 _08681_ (.Y(_02737_),
    .A(net1571),
    .B(net1533));
 sg13g2_nor2_2 _08682_ (.A(_02633_),
    .B(_02737_),
    .Y(_02738_));
 sg13g2_a22oi_1 _08683_ (.Y(_02739_),
    .B1(net1538),
    .B2(net1573),
    .A2(net1533),
    .A1(net1575));
 sg13g2_nor2_1 _08684_ (.A(_02738_),
    .B(_02739_),
    .Y(_02740_));
 sg13g2_nor3_1 _08685_ (.A(_02736_),
    .B(_02738_),
    .C(_02739_),
    .Y(_02741_));
 sg13g2_xor2_1 _08686_ (.B(_02740_),
    .A(_02736_),
    .X(_02742_));
 sg13g2_o21ai_1 _08687_ (.B1(_02641_),
    .Y(_02743_),
    .A1(_02639_),
    .A2(_02642_));
 sg13g2_nand2_1 _08688_ (.Y(_02744_),
    .A(net1581),
    .B(net1528));
 sg13g2_nand2_1 _08689_ (.Y(_02745_),
    .A(net1588),
    .B(net1517));
 sg13g2_and4_1 _08690_ (.A(net1588),
    .B(net1595),
    .C(net1517),
    .D(net1521),
    .X(_02746_));
 sg13g2_a22oi_1 _08691_ (.Y(_02747_),
    .B1(net1521),
    .B2(net1587),
    .A2(net1517),
    .A1(net1595));
 sg13g2_nor3_1 _08692_ (.A(_02744_),
    .B(_02746_),
    .C(_02747_),
    .Y(_02748_));
 sg13g2_o21ai_1 _08693_ (.B1(_02744_),
    .Y(_02749_),
    .A1(_02746_),
    .A2(_02747_));
 sg13g2_nor2b_1 _08694_ (.A(_02748_),
    .B_N(_02749_),
    .Y(_02750_));
 sg13g2_nand2_1 _08695_ (.Y(_02751_),
    .A(_02743_),
    .B(_02750_));
 sg13g2_xnor2_1 _08696_ (.Y(_02752_),
    .A(_02743_),
    .B(_02750_));
 sg13g2_xnor2_1 _08697_ (.Y(_02753_),
    .A(_02742_),
    .B(_02752_));
 sg13g2_nand2b_1 _08698_ (.Y(_02754_),
    .B(_02735_),
    .A_N(_02753_));
 sg13g2_xor2_1 _08699_ (.B(_02753_),
    .A(_02735_),
    .X(_02755_));
 sg13g2_xnor2_1 _08700_ (.Y(_02756_),
    .A(_02734_),
    .B(_02755_));
 sg13g2_o21ai_1 _08701_ (.B1(_02684_),
    .Y(_02757_),
    .A1(_02664_),
    .A2(_02685_));
 sg13g2_o21ai_1 _08702_ (.B1(_02658_),
    .Y(_02758_),
    .A1(_02655_),
    .A2(_02659_));
 sg13g2_inv_1 _08703_ (.Y(_02759_),
    .A(_02758_));
 sg13g2_o21ai_1 _08704_ (.B1(_02668_),
    .Y(_02760_),
    .A1(_02666_),
    .A2(_02669_));
 sg13g2_nand2_1 _08705_ (.Y(_02761_),
    .A(net1599),
    .B(net1731));
 sg13g2_nand2_1 _08706_ (.Y(_02762_),
    .A(net1605),
    .B(net1718));
 sg13g2_nand2_1 _08707_ (.Y(_02763_),
    .A(net1609),
    .B(net1718));
 sg13g2_or2_1 _08708_ (.X(_02764_),
    .B(_02762_),
    .A(_02657_));
 sg13g2_xnor2_1 _08709_ (.Y(_02765_),
    .A(_02656_),
    .B(_02763_));
 sg13g2_xor2_1 _08710_ (.B(_02765_),
    .A(_02761_),
    .X(_02766_));
 sg13g2_nand2_1 _08711_ (.Y(_02767_),
    .A(_02760_),
    .B(_02766_));
 sg13g2_xnor2_1 _08712_ (.Y(_02768_),
    .A(_02760_),
    .B(_02766_));
 sg13g2_xnor2_1 _08713_ (.Y(_02769_),
    .A(_02758_),
    .B(_02768_));
 sg13g2_xnor2_1 _08714_ (.Y(_02770_),
    .A(_02759_),
    .B(_02768_));
 sg13g2_a21o_1 _08715_ (.A2(_02681_),
    .A1(_02671_),
    .B1(_02679_),
    .X(_02771_));
 sg13g2_nand2_1 _08716_ (.Y(_02772_),
    .A(net1613),
    .B(net1713));
 sg13g2_nand2_2 _08717_ (.Y(_02773_),
    .A(net1620),
    .B(net1700));
 sg13g2_and4_1 _08718_ (.A(net1620),
    .B(net1625),
    .C(net1699),
    .D(net1706),
    .X(_02774_));
 sg13g2_or2_1 _08719_ (.X(_02775_),
    .B(_02773_),
    .A(_02667_));
 sg13g2_a22oi_1 _08720_ (.Y(_02776_),
    .B1(net1707),
    .B2(net1620),
    .A2(net1699),
    .A1(net1625));
 sg13g2_nor2_1 _08721_ (.A(_02774_),
    .B(_02776_),
    .Y(_02777_));
 sg13g2_xnor2_1 _08722_ (.Y(_02778_),
    .A(_02772_),
    .B(_02777_));
 sg13g2_o21ai_1 _08723_ (.B1(_02675_),
    .Y(_02779_),
    .A1(_02673_),
    .A2(_02676_));
 sg13g2_nand2_1 _08724_ (.Y(_02780_),
    .A(net1630),
    .B(net1695));
 sg13g2_and4_1 _08725_ (.A(net1642),
    .B(net1652),
    .C(net1686),
    .D(net1689),
    .X(_02781_));
 sg13g2_nand4_1 _08726_ (.B(net1652),
    .C(net1686),
    .A(net1642),
    .Y(_02782_),
    .D(net1690));
 sg13g2_a22oi_1 _08727_ (.Y(_02783_),
    .B1(net1690),
    .B2(net1642),
    .A2(net1686),
    .A1(net1652));
 sg13g2_or3_1 _08728_ (.A(_02780_),
    .B(_02781_),
    .C(_02783_),
    .X(_02784_));
 sg13g2_o21ai_1 _08729_ (.B1(_02780_),
    .Y(_02785_),
    .A1(_02781_),
    .A2(_02783_));
 sg13g2_and3_1 _08730_ (.X(_02786_),
    .A(_02779_),
    .B(_02784_),
    .C(_02785_));
 sg13g2_nand3_1 _08731_ (.B(_02784_),
    .C(_02785_),
    .A(_02779_),
    .Y(_02787_));
 sg13g2_a21o_1 _08732_ (.A2(_02785_),
    .A1(_02784_),
    .B1(_02779_),
    .X(_02788_));
 sg13g2_nand3_1 _08733_ (.B(_02787_),
    .C(_02788_),
    .A(_02778_),
    .Y(_02789_));
 sg13g2_a21o_1 _08734_ (.A2(_02788_),
    .A1(_02787_),
    .B1(_02778_),
    .X(_02790_));
 sg13g2_nand3_1 _08735_ (.B(_02789_),
    .C(_02790_),
    .A(_02771_),
    .Y(_02791_));
 sg13g2_a21oi_1 _08736_ (.A1(_02789_),
    .A2(_02790_),
    .Y(_02792_),
    .B1(_02771_));
 sg13g2_a21o_1 _08737_ (.A2(_02790_),
    .A1(_02789_),
    .B1(_02771_),
    .X(_02793_));
 sg13g2_nand3_1 _08738_ (.B(_02791_),
    .C(_02793_),
    .A(_02769_),
    .Y(_02794_));
 sg13g2_a21o_1 _08739_ (.A2(_02793_),
    .A1(_02791_),
    .B1(_02769_),
    .X(_02795_));
 sg13g2_and3_1 _08740_ (.X(_02796_),
    .A(_02757_),
    .B(_02794_),
    .C(_02795_));
 sg13g2_nand3_1 _08741_ (.B(_02794_),
    .C(_02795_),
    .A(_02757_),
    .Y(_02797_));
 sg13g2_a21oi_1 _08742_ (.A1(_02794_),
    .A2(_02795_),
    .Y(_02798_),
    .B1(_02757_));
 sg13g2_or3_1 _08743_ (.A(_02756_),
    .B(_02796_),
    .C(_02798_),
    .X(_02799_));
 sg13g2_o21ai_1 _08744_ (.B1(_02756_),
    .Y(_02800_),
    .A1(_02796_),
    .A2(_02798_));
 sg13g2_and3_1 _08745_ (.X(_02801_),
    .A(_02732_),
    .B(_02799_),
    .C(_02800_));
 sg13g2_nand3_1 _08746_ (.B(_02799_),
    .C(_02800_),
    .A(_02732_),
    .Y(_02802_));
 sg13g2_a21oi_1 _08747_ (.A1(_02799_),
    .A2(_02800_),
    .Y(_02803_),
    .B1(_02732_));
 sg13g2_or3_1 _08748_ (.A(_02731_),
    .B(_02801_),
    .C(_02803_),
    .X(_02804_));
 sg13g2_o21ai_1 _08749_ (.B1(_02731_),
    .Y(_02805_),
    .A1(_02801_),
    .A2(_02803_));
 sg13g2_and3_1 _08750_ (.X(_02806_),
    .A(_02717_),
    .B(_02804_),
    .C(_02805_));
 sg13g2_nand3_1 _08751_ (.B(_02804_),
    .C(_02805_),
    .A(_02717_),
    .Y(_02807_));
 sg13g2_a21oi_1 _08752_ (.A1(_02804_),
    .A2(_02805_),
    .Y(_02808_),
    .B1(_02717_));
 sg13g2_o21ai_1 _08753_ (.B1(_02627_),
    .Y(_02809_),
    .A1(_02806_),
    .A2(_02808_));
 sg13g2_or3_1 _08754_ (.A(_02627_),
    .B(_02806_),
    .C(_02808_),
    .X(_02810_));
 sg13g2_and3_2 _08755_ (.X(_02811_),
    .A(_02716_),
    .B(_02809_),
    .C(_02810_));
 sg13g2_a21oi_2 _08756_ (.B1(_02716_),
    .Y(_02812_),
    .A2(_02810_),
    .A1(_02809_));
 sg13g2_nor3_1 _08757_ (.A(_02705_),
    .B(_02811_),
    .C(_02812_),
    .Y(_02813_));
 sg13g2_or3_1 _08758_ (.A(_02705_),
    .B(_02811_),
    .C(_02812_),
    .X(_02814_));
 sg13g2_o21ai_1 _08759_ (.B1(_02705_),
    .Y(_02815_),
    .A1(_02811_),
    .A2(_02812_));
 sg13g2_and4_1 _08760_ (.A(_02610_),
    .B(_02706_),
    .C(_02814_),
    .D(_02815_),
    .X(_02816_));
 sg13g2_nand4_1 _08761_ (.B(_02706_),
    .C(_02814_),
    .A(_02610_),
    .Y(_02817_),
    .D(_02815_));
 sg13g2_a22oi_1 _08762_ (.Y(_02818_),
    .B1(_02814_),
    .B2(_02815_),
    .A2(_02706_),
    .A1(_02610_));
 sg13g2_nor2_1 _08763_ (.A(_02816_),
    .B(_02818_),
    .Y(_02819_));
 sg13g2_xnor2_1 _08764_ (.Y(_02820_),
    .A(_02715_),
    .B(_02819_));
 sg13g2_o21ai_1 _08765_ (.B1(net1755),
    .Y(_02821_),
    .A1(net1471),
    .A2(net603));
 sg13g2_a21oi_1 _08766_ (.A1(net1471),
    .A2(_02820_),
    .Y(_00316_),
    .B1(_02821_));
 sg13g2_o21ai_1 _08767_ (.B1(_02802_),
    .Y(_02822_),
    .A1(_02731_),
    .A2(_02803_));
 sg13g2_o21ai_1 _08768_ (.B1(_02754_),
    .Y(_02823_),
    .A1(_02734_),
    .A2(_02755_));
 sg13g2_nand2_1 _08769_ (.Y(_02824_),
    .A(net1509),
    .B(net1556));
 sg13g2_nand2_1 _08770_ (.Y(_02825_),
    .A(net1511),
    .B(net1547));
 sg13g2_nand2_1 _08771_ (.Y(_02826_),
    .A(net1563),
    .B(net1547));
 sg13g2_or2_1 _08772_ (.X(_02827_),
    .B(_02826_),
    .A(_02721_));
 sg13g2_xor2_1 _08773_ (.B(_02826_),
    .A(_02721_),
    .X(_02828_));
 sg13g2_nand2b_1 _08774_ (.Y(_02829_),
    .B(_02828_),
    .A_N(_02824_));
 sg13g2_xnor2_1 _08775_ (.Y(_02830_),
    .A(_02824_),
    .B(_02828_));
 sg13g2_o21ai_1 _08776_ (.B1(_02830_),
    .Y(_02831_),
    .A1(_02738_),
    .A2(_02741_));
 sg13g2_nor3_1 _08777_ (.A(_02738_),
    .B(_02741_),
    .C(_02830_),
    .Y(_02832_));
 sg13g2_or3_1 _08778_ (.A(_02738_),
    .B(_02741_),
    .C(_02830_),
    .X(_02833_));
 sg13g2_and2_1 _08779_ (.A(_02831_),
    .B(_02833_),
    .X(_02834_));
 sg13g2_nor2_1 _08780_ (.A(_02722_),
    .B(_02725_),
    .Y(_02835_));
 sg13g2_xnor2_1 _08781_ (.Y(_02836_),
    .A(_02834_),
    .B(_02835_));
 sg13g2_nand2_1 _08782_ (.Y(_02837_),
    .A(_02823_),
    .B(_02836_));
 sg13g2_xnor2_1 _08783_ (.Y(_02838_),
    .A(_02823_),
    .B(_02836_));
 sg13g2_xnor2_1 _08784_ (.Y(_02839_),
    .A(_02728_),
    .B(_02838_));
 sg13g2_o21ai_1 _08785_ (.B1(_02797_),
    .Y(_02840_),
    .A1(_02756_),
    .A2(_02798_));
 sg13g2_o21ai_1 _08786_ (.B1(_02751_),
    .Y(_02841_),
    .A1(_02742_),
    .A2(_02752_));
 sg13g2_inv_1 _08787_ (.Y(_02842_),
    .A(_02841_));
 sg13g2_o21ai_1 _08788_ (.B1(_02767_),
    .Y(_02843_),
    .A1(_02759_),
    .A2(_02768_));
 sg13g2_nand2_1 _08789_ (.Y(_02844_),
    .A(net1567),
    .B(net1540));
 sg13g2_nand2_2 _08790_ (.Y(_02845_),
    .A(net1575),
    .B(net1528));
 sg13g2_or2_1 _08791_ (.X(_02846_),
    .B(_02845_),
    .A(_02737_));
 sg13g2_and2_1 _08792_ (.A(_02737_),
    .B(_02845_),
    .X(_02847_));
 sg13g2_xnor2_1 _08793_ (.Y(_02848_),
    .A(_02737_),
    .B(_02845_));
 sg13g2_xnor2_1 _08794_ (.Y(_02849_),
    .A(_02844_),
    .B(_02848_));
 sg13g2_or2_1 _08795_ (.X(_02850_),
    .B(_02748_),
    .A(_02746_));
 sg13g2_nand2_1 _08796_ (.Y(_02851_),
    .A(net1582),
    .B(net1521));
 sg13g2_nand2_1 _08797_ (.Y(_02852_),
    .A(net1595),
    .B(net1731));
 sg13g2_or2_1 _08798_ (.X(_02853_),
    .B(_02852_),
    .A(_02745_));
 sg13g2_and2_1 _08799_ (.A(_02745_),
    .B(_02852_),
    .X(_02854_));
 sg13g2_xor2_1 _08800_ (.B(_02852_),
    .A(_02745_),
    .X(_02855_));
 sg13g2_xnor2_1 _08801_ (.Y(_02856_),
    .A(_02851_),
    .B(_02855_));
 sg13g2_nand2_1 _08802_ (.Y(_02857_),
    .A(_02850_),
    .B(_02856_));
 sg13g2_xnor2_1 _08803_ (.Y(_02858_),
    .A(_02850_),
    .B(_02856_));
 sg13g2_xnor2_1 _08804_ (.Y(_02859_),
    .A(_02849_),
    .B(_02858_));
 sg13g2_nand2b_1 _08805_ (.Y(_02860_),
    .B(_02843_),
    .A_N(_02859_));
 sg13g2_xor2_1 _08806_ (.B(_02859_),
    .A(_02843_),
    .X(_02861_));
 sg13g2_xnor2_1 _08807_ (.Y(_02862_),
    .A(_02842_),
    .B(_02861_));
 sg13g2_o21ai_1 _08808_ (.B1(_02791_),
    .Y(_02863_),
    .A1(_02770_),
    .A2(_02792_));
 sg13g2_o21ai_1 _08809_ (.B1(_02764_),
    .Y(_02864_),
    .A1(_02761_),
    .A2(_02765_));
 sg13g2_inv_1 _08810_ (.Y(_02865_),
    .A(_02864_));
 sg13g2_o21ai_1 _08811_ (.B1(_02775_),
    .Y(_02866_),
    .A1(_02772_),
    .A2(_02776_));
 sg13g2_nand2_1 _08812_ (.Y(_02867_),
    .A(net1599),
    .B(net1725));
 sg13g2_nand2_1 _08813_ (.Y(_02868_),
    .A(net1605),
    .B(net1713));
 sg13g2_nand2_1 _08814_ (.Y(_02869_),
    .A(net1609),
    .B(net1713));
 sg13g2_or2_1 _08815_ (.X(_02870_),
    .B(_02868_),
    .A(_02763_));
 sg13g2_xnor2_1 _08816_ (.Y(_02871_),
    .A(_02762_),
    .B(_02869_));
 sg13g2_xor2_1 _08817_ (.B(_02871_),
    .A(_02867_),
    .X(_02872_));
 sg13g2_nand2_1 _08818_ (.Y(_02873_),
    .A(_02866_),
    .B(_02872_));
 sg13g2_xnor2_1 _08819_ (.Y(_02874_),
    .A(_02866_),
    .B(_02872_));
 sg13g2_xnor2_1 _08820_ (.Y(_02875_),
    .A(_02865_),
    .B(_02874_));
 sg13g2_a21o_1 _08821_ (.A2(_02788_),
    .A1(_02778_),
    .B1(_02786_),
    .X(_02876_));
 sg13g2_nand2_1 _08822_ (.Y(_02877_),
    .A(net1614),
    .B(net1707));
 sg13g2_nand2_1 _08823_ (.Y(_02878_),
    .A(net1625),
    .B(net1695));
 sg13g2_or2_1 _08824_ (.X(_02879_),
    .B(_02878_),
    .A(_02773_));
 sg13g2_and2_1 _08825_ (.A(_02773_),
    .B(_02878_),
    .X(_02880_));
 sg13g2_xnor2_1 _08826_ (.Y(_02881_),
    .A(_02773_),
    .B(_02878_));
 sg13g2_xnor2_1 _08827_ (.Y(_02882_),
    .A(_02877_),
    .B(_02881_));
 sg13g2_o21ai_1 _08828_ (.B1(_02782_),
    .Y(_02883_),
    .A1(_02780_),
    .A2(_02783_));
 sg13g2_nand2_1 _08829_ (.Y(_02884_),
    .A(net1632),
    .B(net1690));
 sg13g2_and4_1 _08830_ (.A(net1638),
    .B(net1648),
    .C(net1680),
    .D(net1686),
    .X(_02885_));
 sg13g2_nand4_1 _08831_ (.B(net1648),
    .C(net1680),
    .A(net1638),
    .Y(_02886_),
    .D(net1688));
 sg13g2_a22oi_1 _08832_ (.Y(_02887_),
    .B1(net1688),
    .B2(net1638),
    .A2(net1680),
    .A1(net1648));
 sg13g2_or3_1 _08833_ (.A(_02884_),
    .B(_02885_),
    .C(_02887_),
    .X(_02888_));
 sg13g2_o21ai_1 _08834_ (.B1(_02884_),
    .Y(_02889_),
    .A1(_02885_),
    .A2(_02887_));
 sg13g2_and3_1 _08835_ (.X(_02890_),
    .A(_02883_),
    .B(_02888_),
    .C(_02889_));
 sg13g2_nand3_1 _08836_ (.B(_02888_),
    .C(_02889_),
    .A(_02883_),
    .Y(_02891_));
 sg13g2_a21oi_1 _08837_ (.A1(_02888_),
    .A2(_02889_),
    .Y(_02892_),
    .B1(_02883_));
 sg13g2_or3_1 _08838_ (.A(_02882_),
    .B(_02890_),
    .C(_02892_),
    .X(_02893_));
 sg13g2_o21ai_1 _08839_ (.B1(_02882_),
    .Y(_02894_),
    .A1(_02890_),
    .A2(_02892_));
 sg13g2_and3_1 _08840_ (.X(_02895_),
    .A(_02876_),
    .B(_02893_),
    .C(_02894_));
 sg13g2_nand3_1 _08841_ (.B(_02893_),
    .C(_02894_),
    .A(_02876_),
    .Y(_02896_));
 sg13g2_a21oi_1 _08842_ (.A1(_02893_),
    .A2(_02894_),
    .Y(_02897_),
    .B1(_02876_));
 sg13g2_or3_1 _08843_ (.A(_02875_),
    .B(_02895_),
    .C(_02897_),
    .X(_02898_));
 sg13g2_o21ai_1 _08844_ (.B1(_02875_),
    .Y(_02899_),
    .A1(_02895_),
    .A2(_02897_));
 sg13g2_and3_1 _08845_ (.X(_02900_),
    .A(_02863_),
    .B(_02898_),
    .C(_02899_));
 sg13g2_nand3_1 _08846_ (.B(_02898_),
    .C(_02899_),
    .A(_02863_),
    .Y(_02901_));
 sg13g2_a21oi_1 _08847_ (.A1(_02898_),
    .A2(_02899_),
    .Y(_02902_),
    .B1(_02863_));
 sg13g2_or3_1 _08848_ (.A(_02862_),
    .B(_02900_),
    .C(_02902_),
    .X(_02903_));
 sg13g2_o21ai_1 _08849_ (.B1(_02862_),
    .Y(_02904_),
    .A1(_02900_),
    .A2(_02902_));
 sg13g2_and3_1 _08850_ (.X(_02905_),
    .A(_02840_),
    .B(_02903_),
    .C(_02904_));
 sg13g2_nand3_1 _08851_ (.B(_02903_),
    .C(_02904_),
    .A(_02840_),
    .Y(_02906_));
 sg13g2_a21oi_1 _08852_ (.A1(_02903_),
    .A2(_02904_),
    .Y(_02907_),
    .B1(_02840_));
 sg13g2_or3_1 _08853_ (.A(_02839_),
    .B(_02905_),
    .C(_02907_),
    .X(_02908_));
 sg13g2_o21ai_1 _08854_ (.B1(_02839_),
    .Y(_02909_),
    .A1(_02905_),
    .A2(_02907_));
 sg13g2_and3_1 _08855_ (.X(_02910_),
    .A(_02822_),
    .B(_02908_),
    .C(_02909_));
 sg13g2_nand3_1 _08856_ (.B(_02908_),
    .C(_02909_),
    .A(_02822_),
    .Y(_02911_));
 sg13g2_a21oi_1 _08857_ (.A1(_02908_),
    .A2(_02909_),
    .Y(_02912_),
    .B1(_02822_));
 sg13g2_o21ai_1 _08858_ (.B1(_02730_),
    .Y(_02913_),
    .A1(_02910_),
    .A2(_02912_));
 sg13g2_or3_1 _08859_ (.A(_02730_),
    .B(_02910_),
    .C(_02912_),
    .X(_02914_));
 sg13g2_o21ai_1 _08860_ (.B1(_02807_),
    .Y(_02915_),
    .A1(_02627_),
    .A2(_02808_));
 sg13g2_nand3_1 _08861_ (.B(_02914_),
    .C(_02915_),
    .A(_02913_),
    .Y(_02916_));
 sg13g2_a21o_2 _08862_ (.A2(_02914_),
    .A1(_02913_),
    .B1(_02915_),
    .X(_02917_));
 sg13g2_and3_1 _08863_ (.X(_02918_),
    .A(_02811_),
    .B(_02916_),
    .C(_02917_));
 sg13g2_nand3_1 _08864_ (.B(_02916_),
    .C(_02917_),
    .A(_02811_),
    .Y(_02919_));
 sg13g2_a21o_1 _08865_ (.A2(_02917_),
    .A1(_02916_),
    .B1(_02811_),
    .X(_02920_));
 sg13g2_a21oi_1 _08866_ (.A1(_02919_),
    .A2(_02920_),
    .Y(_02921_),
    .B1(_02813_));
 sg13g2_and3_1 _08867_ (.X(_02922_),
    .A(_02813_),
    .B(_02919_),
    .C(_02920_));
 sg13g2_nand3_1 _08868_ (.B(_02919_),
    .C(_02920_),
    .A(_02813_),
    .Y(_02923_));
 sg13g2_nor2_1 _08869_ (.A(_02921_),
    .B(_02922_),
    .Y(_02924_));
 sg13g2_a21oi_1 _08870_ (.A1(_02715_),
    .A2(_02819_),
    .Y(_02925_),
    .B1(_02816_));
 sg13g2_xor2_1 _08871_ (.B(_02925_),
    .A(_02924_),
    .X(_02926_));
 sg13g2_o21ai_1 _08872_ (.B1(net1755),
    .Y(_02927_),
    .A1(net1469),
    .A2(net597));
 sg13g2_a21oi_1 _08873_ (.A1(net1469),
    .A2(_02926_),
    .Y(_00317_),
    .B1(_02927_));
 sg13g2_o21ai_1 _08874_ (.B1(_02911_),
    .Y(_02928_),
    .A1(_02730_),
    .A2(_02912_));
 sg13g2_o21ai_1 _08875_ (.B1(_02837_),
    .Y(_02929_),
    .A1(_02728_),
    .A2(_02838_));
 sg13g2_o21ai_1 _08876_ (.B1(_02906_),
    .Y(_02930_),
    .A1(_02839_),
    .A2(_02907_));
 sg13g2_and2_1 _08877_ (.A(_02725_),
    .B(_02834_),
    .X(_02931_));
 sg13g2_inv_1 _08878_ (.Y(_02932_),
    .A(_02931_));
 sg13g2_o21ai_1 _08879_ (.B1(_02860_),
    .Y(_02933_),
    .A1(_02842_),
    .A2(_02861_));
 sg13g2_nand2_2 _08880_ (.Y(_02934_),
    .A(net1505),
    .B(net1556));
 sg13g2_and2_1 _08881_ (.A(_02827_),
    .B(_02829_),
    .X(_02935_));
 sg13g2_o21ai_1 _08882_ (.B1(_02846_),
    .Y(_02936_),
    .A1(_02844_),
    .A2(_02847_));
 sg13g2_nand2_1 _08883_ (.Y(_02937_),
    .A(net1509),
    .B(net1553));
 sg13g2_nand2_1 _08884_ (.Y(_02938_),
    .A(net1511),
    .B(net1540));
 sg13g2_nand2_1 _08885_ (.Y(_02939_),
    .A(net1563),
    .B(net1540));
 sg13g2_or2_1 _08886_ (.X(_02940_),
    .B(_02938_),
    .A(_02826_));
 sg13g2_xnor2_1 _08887_ (.Y(_02941_),
    .A(_02825_),
    .B(_02939_));
 sg13g2_xor2_1 _08888_ (.B(_02941_),
    .A(_02937_),
    .X(_02942_));
 sg13g2_nand2_1 _08889_ (.Y(_02943_),
    .A(_02936_),
    .B(_02942_));
 sg13g2_xnor2_1 _08890_ (.Y(_02944_),
    .A(_02936_),
    .B(_02942_));
 sg13g2_xor2_1 _08891_ (.B(_02944_),
    .A(_02935_),
    .X(_02945_));
 sg13g2_a21oi_1 _08892_ (.A1(_02723_),
    .A2(_02831_),
    .Y(_02946_),
    .B1(_02832_));
 sg13g2_xor2_1 _08893_ (.B(_02946_),
    .A(_02945_),
    .X(_02947_));
 sg13g2_nor2b_1 _08894_ (.A(_02934_),
    .B_N(_02947_),
    .Y(_02948_));
 sg13g2_xnor2_1 _08895_ (.Y(_02949_),
    .A(_02934_),
    .B(_02947_));
 sg13g2_nand2_1 _08896_ (.Y(_02950_),
    .A(_02933_),
    .B(_02949_));
 sg13g2_xnor2_1 _08897_ (.Y(_02951_),
    .A(_02933_),
    .B(_02949_));
 sg13g2_xnor2_1 _08898_ (.Y(_02952_),
    .A(_02932_),
    .B(_02951_));
 sg13g2_o21ai_1 _08899_ (.B1(_02901_),
    .Y(_02953_),
    .A1(_02862_),
    .A2(_02902_));
 sg13g2_o21ai_1 _08900_ (.B1(_02857_),
    .Y(_02954_),
    .A1(_02849_),
    .A2(_02858_));
 sg13g2_inv_1 _08901_ (.Y(_02955_),
    .A(_02954_));
 sg13g2_o21ai_1 _08902_ (.B1(_02873_),
    .Y(_02956_),
    .A1(_02865_),
    .A2(_02874_));
 sg13g2_nand2_1 _08903_ (.Y(_02957_),
    .A(net1567),
    .B(net1533));
 sg13g2_nand2_2 _08904_ (.Y(_02958_),
    .A(net1573),
    .B(net1521));
 sg13g2_nor2_1 _08905_ (.A(_02845_),
    .B(_02958_),
    .Y(_02959_));
 sg13g2_or2_1 _08906_ (.X(_02960_),
    .B(_02958_),
    .A(_02845_));
 sg13g2_a22oi_1 _08907_ (.Y(_02961_),
    .B1(net1528),
    .B2(net1571),
    .A2(net1521),
    .A1(net1575));
 sg13g2_nor3_1 _08908_ (.A(_02957_),
    .B(_02959_),
    .C(_02961_),
    .Y(_02962_));
 sg13g2_o21ai_1 _08909_ (.B1(_02957_),
    .Y(_02963_),
    .A1(_02959_),
    .A2(_02961_));
 sg13g2_nand2b_1 _08910_ (.Y(_02964_),
    .B(_02963_),
    .A_N(_02962_));
 sg13g2_o21ai_1 _08911_ (.B1(_02853_),
    .Y(_02965_),
    .A1(_02851_),
    .A2(_02854_));
 sg13g2_nand2_1 _08912_ (.Y(_02966_),
    .A(net1582),
    .B(net1517));
 sg13g2_nand2_1 _08913_ (.Y(_02967_),
    .A(net1585),
    .B(net1725));
 sg13g2_and4_1 _08914_ (.A(net1587),
    .B(net1594),
    .C(net1725),
    .D(net1731),
    .X(_02968_));
 sg13g2_a22oi_1 _08915_ (.Y(_02969_),
    .B1(net1731),
    .B2(net1587),
    .A2(net1725),
    .A1(net1594));
 sg13g2_nor3_1 _08916_ (.A(_02966_),
    .B(_02968_),
    .C(_02969_),
    .Y(_02970_));
 sg13g2_o21ai_1 _08917_ (.B1(_02966_),
    .Y(_02971_),
    .A1(_02968_),
    .A2(_02969_));
 sg13g2_nor2b_1 _08918_ (.A(_02970_),
    .B_N(_02971_),
    .Y(_02972_));
 sg13g2_nand2_1 _08919_ (.Y(_02973_),
    .A(_02965_),
    .B(_02972_));
 sg13g2_xnor2_1 _08920_ (.Y(_02974_),
    .A(_02965_),
    .B(_02972_));
 sg13g2_xnor2_1 _08921_ (.Y(_02975_),
    .A(_02964_),
    .B(_02974_));
 sg13g2_nand2b_1 _08922_ (.Y(_02976_),
    .B(_02956_),
    .A_N(_02975_));
 sg13g2_xor2_1 _08923_ (.B(_02975_),
    .A(_02956_),
    .X(_02977_));
 sg13g2_xnor2_1 _08924_ (.Y(_02978_),
    .A(_02955_),
    .B(_02977_));
 sg13g2_o21ai_1 _08925_ (.B1(_02896_),
    .Y(_02979_),
    .A1(_02875_),
    .A2(_02897_));
 sg13g2_o21ai_1 _08926_ (.B1(_02870_),
    .Y(_02980_),
    .A1(_02867_),
    .A2(_02871_));
 sg13g2_inv_1 _08927_ (.Y(_02981_),
    .A(_02980_));
 sg13g2_o21ai_1 _08928_ (.B1(_02879_),
    .Y(_02982_),
    .A1(_02877_),
    .A2(_02880_));
 sg13g2_nand2_1 _08929_ (.Y(_02983_),
    .A(net1600),
    .B(net1718));
 sg13g2_nand2_1 _08930_ (.Y(_02984_),
    .A(net1603),
    .B(net1707));
 sg13g2_nand2_1 _08931_ (.Y(_02985_),
    .A(net1608),
    .B(net1707));
 sg13g2_or2_1 _08932_ (.X(_02986_),
    .B(_02984_),
    .A(_02869_));
 sg13g2_xnor2_1 _08933_ (.Y(_02987_),
    .A(_02868_),
    .B(_02985_));
 sg13g2_xor2_1 _08934_ (.B(_02987_),
    .A(_02983_),
    .X(_02988_));
 sg13g2_nand2_1 _08935_ (.Y(_02989_),
    .A(_02982_),
    .B(_02988_));
 sg13g2_xnor2_1 _08936_ (.Y(_02990_),
    .A(_02982_),
    .B(_02988_));
 sg13g2_xnor2_1 _08937_ (.Y(_02991_),
    .A(_02981_),
    .B(_02990_));
 sg13g2_o21ai_1 _08938_ (.B1(_02891_),
    .Y(_02992_),
    .A1(_02882_),
    .A2(_02892_));
 sg13g2_nand2_1 _08939_ (.Y(_02993_),
    .A(net1612),
    .B(net1700));
 sg13g2_nand2_1 _08940_ (.Y(_02994_),
    .A(net1618),
    .B(net1689));
 sg13g2_and4_1 _08941_ (.A(net1618),
    .B(net1623),
    .C(net1689),
    .D(net1694),
    .X(_02995_));
 sg13g2_a22oi_1 _08942_ (.Y(_02996_),
    .B1(net1694),
    .B2(net1618),
    .A2(net1689),
    .A1(net1624));
 sg13g2_nor3_1 _08943_ (.A(_02993_),
    .B(_02995_),
    .C(_02996_),
    .Y(_02997_));
 sg13g2_o21ai_1 _08944_ (.B1(_02993_),
    .Y(_02998_),
    .A1(_02995_),
    .A2(_02996_));
 sg13g2_nand2b_1 _08945_ (.Y(_02999_),
    .B(_02998_),
    .A_N(_02997_));
 sg13g2_o21ai_1 _08946_ (.B1(_02886_),
    .Y(_03000_),
    .A1(_02884_),
    .A2(_02887_));
 sg13g2_nand2_1 _08947_ (.Y(_03001_),
    .A(net1631),
    .B(net1686));
 sg13g2_and4_1 _08948_ (.A(net1638),
    .B(net1649),
    .C(net1675),
    .D(net1680),
    .X(_03002_));
 sg13g2_nand4_1 _08949_ (.B(net1648),
    .C(net1675),
    .A(net1638),
    .Y(_03003_),
    .D(net1680));
 sg13g2_a22oi_1 _08950_ (.Y(_03004_),
    .B1(net1681),
    .B2(net1639),
    .A2(net1676),
    .A1(net1648));
 sg13g2_or3_1 _08951_ (.A(_03001_),
    .B(_03002_),
    .C(_03004_),
    .X(_03005_));
 sg13g2_o21ai_1 _08952_ (.B1(_03001_),
    .Y(_03006_),
    .A1(_03002_),
    .A2(_03004_));
 sg13g2_and3_1 _08953_ (.X(_03007_),
    .A(_03000_),
    .B(_03005_),
    .C(_03006_));
 sg13g2_nand3_1 _08954_ (.B(_03005_),
    .C(_03006_),
    .A(_03000_),
    .Y(_03008_));
 sg13g2_a21oi_1 _08955_ (.A1(_03005_),
    .A2(_03006_),
    .Y(_03009_),
    .B1(_03000_));
 sg13g2_or3_1 _08956_ (.A(_02999_),
    .B(_03007_),
    .C(_03009_),
    .X(_03010_));
 sg13g2_o21ai_1 _08957_ (.B1(_02999_),
    .Y(_03011_),
    .A1(_03007_),
    .A2(_03009_));
 sg13g2_and3_1 _08958_ (.X(_03012_),
    .A(_02992_),
    .B(_03010_),
    .C(_03011_));
 sg13g2_nand3_1 _08959_ (.B(_03010_),
    .C(_03011_),
    .A(_02992_),
    .Y(_03013_));
 sg13g2_a21oi_1 _08960_ (.A1(_03010_),
    .A2(_03011_),
    .Y(_03014_),
    .B1(_02992_));
 sg13g2_or3_1 _08961_ (.A(_02991_),
    .B(_03012_),
    .C(_03014_),
    .X(_03015_));
 sg13g2_o21ai_1 _08962_ (.B1(_02991_),
    .Y(_03016_),
    .A1(_03012_),
    .A2(_03014_));
 sg13g2_and3_1 _08963_ (.X(_03017_),
    .A(_02979_),
    .B(_03015_),
    .C(_03016_));
 sg13g2_nand3_1 _08964_ (.B(_03015_),
    .C(_03016_),
    .A(_02979_),
    .Y(_03018_));
 sg13g2_a21oi_1 _08965_ (.A1(_03015_),
    .A2(_03016_),
    .Y(_03019_),
    .B1(_02979_));
 sg13g2_or3_1 _08966_ (.A(_02978_),
    .B(_03017_),
    .C(_03019_),
    .X(_03020_));
 sg13g2_o21ai_1 _08967_ (.B1(_02978_),
    .Y(_03021_),
    .A1(_03017_),
    .A2(_03019_));
 sg13g2_and3_1 _08968_ (.X(_03022_),
    .A(_02953_),
    .B(_03020_),
    .C(_03021_));
 sg13g2_a21oi_1 _08969_ (.A1(_03020_),
    .A2(_03021_),
    .Y(_03023_),
    .B1(_02953_));
 sg13g2_or3_1 _08970_ (.A(_02952_),
    .B(_03022_),
    .C(_03023_),
    .X(_03024_));
 sg13g2_o21ai_1 _08971_ (.B1(_02952_),
    .Y(_03025_),
    .A1(_03022_),
    .A2(_03023_));
 sg13g2_nand3_1 _08972_ (.B(_03024_),
    .C(_03025_),
    .A(_02930_),
    .Y(_03026_));
 sg13g2_a21o_1 _08973_ (.A2(_03025_),
    .A1(_03024_),
    .B1(_02930_),
    .X(_03027_));
 sg13g2_a21o_1 _08974_ (.A2(_03027_),
    .A1(_03026_),
    .B1(_02929_),
    .X(_03028_));
 sg13g2_nand3_1 _08975_ (.B(_03026_),
    .C(_03027_),
    .A(_02929_),
    .Y(_03029_));
 sg13g2_and3_1 _08976_ (.X(_03030_),
    .A(_02928_),
    .B(_03028_),
    .C(_03029_));
 sg13g2_nand3_1 _08977_ (.B(_03028_),
    .C(_03029_),
    .A(_02928_),
    .Y(_03031_));
 sg13g2_a21oi_1 _08978_ (.A1(_03028_),
    .A2(_03029_),
    .Y(_03032_),
    .B1(_02928_));
 sg13g2_or3_1 _08979_ (.A(_02916_),
    .B(_03030_),
    .C(_03032_),
    .X(_03033_));
 sg13g2_o21ai_1 _08980_ (.B1(_02916_),
    .Y(_03034_),
    .A1(_03030_),
    .A2(_03032_));
 sg13g2_nand3_1 _08981_ (.B(_03033_),
    .C(_03034_),
    .A(_02918_),
    .Y(_03035_));
 sg13g2_a21o_1 _08982_ (.A2(_03034_),
    .A1(_03033_),
    .B1(_02918_),
    .X(_03036_));
 sg13g2_and2_1 _08983_ (.A(_03035_),
    .B(_03036_),
    .X(_03037_));
 sg13g2_nor4_1 _08984_ (.A(_02816_),
    .B(_02818_),
    .C(_02921_),
    .D(_02922_),
    .Y(_03038_));
 sg13g2_o21ai_1 _08985_ (.B1(_03038_),
    .Y(_03039_),
    .A1(_02710_),
    .A2(_02714_));
 sg13g2_o21ai_1 _08986_ (.B1(_02923_),
    .Y(_03040_),
    .A1(_02817_),
    .A2(_02921_));
 sg13g2_a21oi_1 _08987_ (.A1(_02715_),
    .A2(_03038_),
    .Y(_03041_),
    .B1(_03040_));
 sg13g2_nand2b_1 _08988_ (.Y(_03042_),
    .B(_03037_),
    .A_N(_03041_));
 sg13g2_xnor2_1 _08989_ (.Y(_03043_),
    .A(_03037_),
    .B(_03041_));
 sg13g2_o21ai_1 _08990_ (.B1(net1751),
    .Y(_03044_),
    .A1(net1398),
    .A2(_03043_));
 sg13g2_a21oi_1 _08991_ (.A1(net1398),
    .A2(_05549_),
    .Y(_00318_),
    .B1(_03044_));
 sg13g2_nand2_1 _08992_ (.Y(_03045_),
    .A(_03035_),
    .B(_03042_));
 sg13g2_o21ai_1 _08993_ (.B1(_02950_),
    .Y(_03046_),
    .A1(_02932_),
    .A2(_02951_));
 sg13g2_inv_1 _08994_ (.Y(_03047_),
    .A(_03046_));
 sg13g2_nand2b_1 _08995_ (.Y(_03048_),
    .B(_03024_),
    .A_N(_03022_));
 sg13g2_o21ai_1 _08996_ (.B1(_03018_),
    .Y(_03049_),
    .A1(_02978_),
    .A2(_03019_));
 sg13g2_o21ai_1 _08997_ (.B1(_02973_),
    .Y(_03050_),
    .A1(_02964_),
    .A2(_02974_));
 sg13g2_inv_1 _08998_ (.Y(_03051_),
    .A(_03050_));
 sg13g2_o21ai_1 _08999_ (.B1(_02989_),
    .Y(_03052_),
    .A1(_02981_),
    .A2(_02990_));
 sg13g2_nand2_1 _09000_ (.Y(_03053_),
    .A(net1569),
    .B(net1528));
 sg13g2_nand2_2 _09001_ (.Y(_03054_),
    .A(net1577),
    .B(net1514));
 sg13g2_or2_1 _09002_ (.X(_03055_),
    .B(_03054_),
    .A(_02958_));
 sg13g2_and2_1 _09003_ (.A(_02958_),
    .B(_03054_),
    .X(_03056_));
 sg13g2_xnor2_1 _09004_ (.Y(_03057_),
    .A(_02958_),
    .B(_03054_));
 sg13g2_xnor2_1 _09005_ (.Y(_03058_),
    .A(_03053_),
    .B(_03057_));
 sg13g2_or2_1 _09006_ (.X(_03059_),
    .B(_02970_),
    .A(_02968_));
 sg13g2_nand2_1 _09007_ (.Y(_03060_),
    .A(net1580),
    .B(net1731));
 sg13g2_nand2_1 _09008_ (.Y(_03061_),
    .A(net1592),
    .B(net1718));
 sg13g2_or2_1 _09009_ (.X(_03062_),
    .B(_03061_),
    .A(_02967_));
 sg13g2_and2_1 _09010_ (.A(_02967_),
    .B(_03061_),
    .X(_03063_));
 sg13g2_xor2_1 _09011_ (.B(_03061_),
    .A(_02967_),
    .X(_03064_));
 sg13g2_xnor2_1 _09012_ (.Y(_03065_),
    .A(_03060_),
    .B(_03064_));
 sg13g2_nand2_1 _09013_ (.Y(_03066_),
    .A(_03059_),
    .B(_03065_));
 sg13g2_xnor2_1 _09014_ (.Y(_03067_),
    .A(_03059_),
    .B(_03065_));
 sg13g2_xnor2_1 _09015_ (.Y(_03068_),
    .A(_03058_),
    .B(_03067_));
 sg13g2_nand2b_1 _09016_ (.Y(_03069_),
    .B(_03052_),
    .A_N(_03068_));
 sg13g2_xor2_1 _09017_ (.B(_03068_),
    .A(_03052_),
    .X(_03070_));
 sg13g2_xnor2_1 _09018_ (.Y(_03071_),
    .A(_03051_),
    .B(_03070_));
 sg13g2_o21ai_1 _09019_ (.B1(_03013_),
    .Y(_03072_),
    .A1(_02991_),
    .A2(_03014_));
 sg13g2_o21ai_1 _09020_ (.B1(_02986_),
    .Y(_03073_),
    .A1(_02983_),
    .A2(_02987_));
 sg13g2_inv_1 _09021_ (.Y(_03074_),
    .A(_03073_));
 sg13g2_or2_1 _09022_ (.X(_03075_),
    .B(_02997_),
    .A(_02995_));
 sg13g2_nand2_1 _09023_ (.Y(_03076_),
    .A(net1598),
    .B(net1713));
 sg13g2_nand2_1 _09024_ (.Y(_03077_),
    .A(net1603),
    .B(net1700));
 sg13g2_nand2_1 _09025_ (.Y(_03078_),
    .A(net1607),
    .B(net1700));
 sg13g2_or2_1 _09026_ (.X(_03079_),
    .B(_03077_),
    .A(_02985_));
 sg13g2_xnor2_1 _09027_ (.Y(_03080_),
    .A(_02984_),
    .B(_03078_));
 sg13g2_xor2_1 _09028_ (.B(_03080_),
    .A(_03076_),
    .X(_03081_));
 sg13g2_nand2_1 _09029_ (.Y(_03082_),
    .A(_03075_),
    .B(_03081_));
 sg13g2_xnor2_1 _09030_ (.Y(_03083_),
    .A(_03075_),
    .B(_03081_));
 sg13g2_xnor2_1 _09031_ (.Y(_03084_),
    .A(_03074_),
    .B(_03083_));
 sg13g2_o21ai_1 _09032_ (.B1(_03008_),
    .Y(_03085_),
    .A1(_02999_),
    .A2(_03009_));
 sg13g2_nand2_1 _09033_ (.Y(_03086_),
    .A(net1612),
    .B(net1694));
 sg13g2_nand2_1 _09034_ (.Y(_03087_),
    .A(net1624),
    .B(net1686));
 sg13g2_or2_1 _09035_ (.X(_03088_),
    .B(_03087_),
    .A(_02994_));
 sg13g2_and2_1 _09036_ (.A(_02994_),
    .B(_03087_),
    .X(_03089_));
 sg13g2_xnor2_1 _09037_ (.Y(_03090_),
    .A(_02994_),
    .B(_03087_));
 sg13g2_xnor2_1 _09038_ (.Y(_03091_),
    .A(_03086_),
    .B(_03090_));
 sg13g2_o21ai_1 _09039_ (.B1(_03003_),
    .Y(_03092_),
    .A1(_03001_),
    .A2(_03004_));
 sg13g2_nand2_1 _09040_ (.Y(_03093_),
    .A(net1631),
    .B(net1681));
 sg13g2_and4_1 _09041_ (.A(net1638),
    .B(net1648),
    .C(net1672),
    .D(net1676),
    .X(_03094_));
 sg13g2_nand4_1 _09042_ (.B(net1648),
    .C(net1671),
    .A(net1638),
    .Y(_03095_),
    .D(net1676));
 sg13g2_a22oi_1 _09043_ (.Y(_03096_),
    .B1(net1676),
    .B2(net1638),
    .A2(net1672),
    .A1(net1648));
 sg13g2_or3_1 _09044_ (.A(_03093_),
    .B(_03094_),
    .C(_03096_),
    .X(_03097_));
 sg13g2_o21ai_1 _09045_ (.B1(_03093_),
    .Y(_03098_),
    .A1(_03094_),
    .A2(_03096_));
 sg13g2_and3_1 _09046_ (.X(_03099_),
    .A(_03092_),
    .B(_03097_),
    .C(_03098_));
 sg13g2_nand3_1 _09047_ (.B(_03097_),
    .C(_03098_),
    .A(_03092_),
    .Y(_03100_));
 sg13g2_a21oi_1 _09048_ (.A1(_03097_),
    .A2(_03098_),
    .Y(_03101_),
    .B1(_03092_));
 sg13g2_or3_1 _09049_ (.A(_03091_),
    .B(_03099_),
    .C(_03101_),
    .X(_03102_));
 sg13g2_o21ai_1 _09050_ (.B1(_03091_),
    .Y(_03103_),
    .A1(_03099_),
    .A2(_03101_));
 sg13g2_and3_1 _09051_ (.X(_03104_),
    .A(_03085_),
    .B(_03102_),
    .C(_03103_));
 sg13g2_nand3_1 _09052_ (.B(_03102_),
    .C(_03103_),
    .A(_03085_),
    .Y(_03105_));
 sg13g2_a21oi_1 _09053_ (.A1(_03102_),
    .A2(_03103_),
    .Y(_03106_),
    .B1(_03085_));
 sg13g2_or3_1 _09054_ (.A(_03084_),
    .B(_03104_),
    .C(_03106_),
    .X(_03107_));
 sg13g2_o21ai_1 _09055_ (.B1(_03084_),
    .Y(_03108_),
    .A1(_03104_),
    .A2(_03106_));
 sg13g2_and3_1 _09056_ (.X(_03109_),
    .A(_03072_),
    .B(_03107_),
    .C(_03108_));
 sg13g2_nand3_1 _09057_ (.B(_03107_),
    .C(_03108_),
    .A(_03072_),
    .Y(_03110_));
 sg13g2_a21oi_1 _09058_ (.A1(_03107_),
    .A2(_03108_),
    .Y(_03111_),
    .B1(_03072_));
 sg13g2_or3_1 _09059_ (.A(_03071_),
    .B(_03109_),
    .C(_03111_),
    .X(_03112_));
 sg13g2_o21ai_1 _09060_ (.B1(_03071_),
    .Y(_03113_),
    .A1(_03109_),
    .A2(_03111_));
 sg13g2_nand3_1 _09061_ (.B(_03112_),
    .C(_03113_),
    .A(_03049_),
    .Y(_03114_));
 sg13g2_a21o_1 _09062_ (.A2(_03113_),
    .A1(_03112_),
    .B1(_03049_),
    .X(_03115_));
 sg13g2_nand2_1 _09063_ (.Y(_03116_),
    .A(_03114_),
    .B(_03115_));
 sg13g2_a21o_1 _09064_ (.A2(_02946_),
    .A1(_02945_),
    .B1(_02948_),
    .X(_03117_));
 sg13g2_o21ai_1 _09065_ (.B1(_02976_),
    .Y(_03118_),
    .A1(_02955_),
    .A2(_02977_));
 sg13g2_a22oi_1 _09066_ (.Y(_03119_),
    .B1(net1556),
    .B2(net1501),
    .A2(net1553),
    .A1(net1505));
 sg13g2_nand2_2 _09067_ (.Y(_03120_),
    .A(net1501),
    .B(net1553));
 sg13g2_nor2_2 _09068_ (.A(_02934_),
    .B(_03120_),
    .Y(_03121_));
 sg13g2_o21ai_1 _09069_ (.B1(_02943_),
    .Y(_03122_),
    .A1(_02935_),
    .A2(_02944_));
 sg13g2_o21ai_1 _09070_ (.B1(_02940_),
    .Y(_03123_),
    .A1(_02937_),
    .A2(_02941_));
 sg13g2_inv_1 _09071_ (.Y(_03124_),
    .A(_03123_));
 sg13g2_o21ai_1 _09072_ (.B1(_02960_),
    .Y(_03125_),
    .A1(_02957_),
    .A2(_02961_));
 sg13g2_nand2_1 _09073_ (.Y(_03126_),
    .A(net1509),
    .B(net1547));
 sg13g2_nand2_1 _09074_ (.Y(_03127_),
    .A(net1511),
    .B(net1533));
 sg13g2_nand2_1 _09075_ (.Y(_03128_),
    .A(net1563),
    .B(net1533));
 sg13g2_or2_1 _09076_ (.X(_03129_),
    .B(_03127_),
    .A(_02939_));
 sg13g2_xnor2_1 _09077_ (.Y(_03130_),
    .A(_02938_),
    .B(_03128_));
 sg13g2_xor2_1 _09078_ (.B(_03130_),
    .A(_03126_),
    .X(_03131_));
 sg13g2_nand2_1 _09079_ (.Y(_03132_),
    .A(_03125_),
    .B(_03131_));
 sg13g2_xnor2_1 _09080_ (.Y(_03133_),
    .A(_03125_),
    .B(_03131_));
 sg13g2_xnor2_1 _09081_ (.Y(_03134_),
    .A(_03123_),
    .B(_03133_));
 sg13g2_xnor2_1 _09082_ (.Y(_03135_),
    .A(_03122_),
    .B(_03134_));
 sg13g2_nor3_1 _09083_ (.A(_03119_),
    .B(_03121_),
    .C(_03135_),
    .Y(_03136_));
 sg13g2_o21ai_1 _09084_ (.B1(_03135_),
    .Y(_03137_),
    .A1(_03119_),
    .A2(_03121_));
 sg13g2_nand2b_1 _09085_ (.Y(_03138_),
    .B(_03137_),
    .A_N(_03136_));
 sg13g2_nand2b_1 _09086_ (.Y(_03139_),
    .B(_03118_),
    .A_N(_03138_));
 sg13g2_xor2_1 _09087_ (.B(_03138_),
    .A(_03118_),
    .X(_03140_));
 sg13g2_nand2b_1 _09088_ (.Y(_03141_),
    .B(_03117_),
    .A_N(_03140_));
 sg13g2_xor2_1 _09089_ (.B(_03140_),
    .A(_03117_),
    .X(_03142_));
 sg13g2_xor2_1 _09090_ (.B(_03142_),
    .A(_03116_),
    .X(_03143_));
 sg13g2_nand2_1 _09091_ (.Y(_03144_),
    .A(_03048_),
    .B(_03143_));
 sg13g2_xnor2_1 _09092_ (.Y(_03145_),
    .A(_03048_),
    .B(_03143_));
 sg13g2_xnor2_1 _09093_ (.Y(_03146_),
    .A(_03047_),
    .B(_03145_));
 sg13g2_nand2_1 _09094_ (.Y(_03147_),
    .A(_03026_),
    .B(_03029_));
 sg13g2_nand2b_1 _09095_ (.Y(_03148_),
    .B(_03147_),
    .A_N(_03146_));
 sg13g2_xor2_1 _09096_ (.B(_03147_),
    .A(_03146_),
    .X(_03149_));
 sg13g2_nor2_1 _09097_ (.A(_03031_),
    .B(_03149_),
    .Y(_03150_));
 sg13g2_xnor2_1 _09098_ (.Y(_03151_),
    .A(_03031_),
    .B(_03149_));
 sg13g2_xor2_1 _09099_ (.B(_03151_),
    .A(_03033_),
    .X(_03152_));
 sg13g2_xnor2_1 _09100_ (.Y(_03153_),
    .A(_03045_),
    .B(_03152_));
 sg13g2_inv_1 _09101_ (.Y(_03154_),
    .A(_03153_));
 sg13g2_o21ai_1 _09102_ (.B1(net1751),
    .Y(_03155_),
    .A1(net1470),
    .A2(net580));
 sg13g2_a21oi_1 _09103_ (.A1(net1470),
    .A2(_03153_),
    .Y(_00319_),
    .B1(_03155_));
 sg13g2_nand2_1 _09104_ (.Y(_03156_),
    .A(_03139_),
    .B(_03141_));
 sg13g2_inv_1 _09105_ (.Y(_03157_),
    .A(_03156_));
 sg13g2_o21ai_1 _09106_ (.B1(_03114_),
    .Y(_03158_),
    .A1(_03116_),
    .A2(_03142_));
 sg13g2_o21ai_1 _09107_ (.B1(_03110_),
    .Y(_03159_),
    .A1(_03071_),
    .A2(_03111_));
 sg13g2_o21ai_1 _09108_ (.B1(_03066_),
    .Y(_03160_),
    .A1(_03058_),
    .A2(_03067_));
 sg13g2_inv_1 _09109_ (.Y(_03161_),
    .A(_03160_));
 sg13g2_o21ai_1 _09110_ (.B1(_03082_),
    .Y(_03162_),
    .A1(_03074_),
    .A2(_03083_));
 sg13g2_nand2_1 _09111_ (.Y(_03163_),
    .A(net1566),
    .B(net1520));
 sg13g2_nand2_2 _09112_ (.Y(_03164_),
    .A(net1570),
    .B(net1728));
 sg13g2_nor2_1 _09113_ (.A(_03054_),
    .B(_03164_),
    .Y(_03165_));
 sg13g2_or2_1 _09114_ (.X(_03166_),
    .B(_03164_),
    .A(_03054_));
 sg13g2_a22oi_1 _09115_ (.Y(_03167_),
    .B1(net1514),
    .B2(net1570),
    .A2(net1729),
    .A1(net1574));
 sg13g2_nor3_1 _09116_ (.A(_03163_),
    .B(_03165_),
    .C(_03167_),
    .Y(_03168_));
 sg13g2_o21ai_1 _09117_ (.B1(_03163_),
    .Y(_03169_),
    .A1(_03165_),
    .A2(_03167_));
 sg13g2_nand2b_1 _09118_ (.Y(_03170_),
    .B(_03169_),
    .A_N(_03168_));
 sg13g2_o21ai_1 _09119_ (.B1(_03062_),
    .Y(_03171_),
    .A1(_03060_),
    .A2(_03063_));
 sg13g2_nand2_1 _09120_ (.Y(_03172_),
    .A(net1580),
    .B(net1722));
 sg13g2_nand2_1 _09121_ (.Y(_03173_),
    .A(net1585),
    .B(net1710));
 sg13g2_and4_1 _09122_ (.A(net1585),
    .B(net1592),
    .C(net1710),
    .D(net1715),
    .X(_03174_));
 sg13g2_a22oi_1 _09123_ (.Y(_03175_),
    .B1(net1715),
    .B2(net1586),
    .A2(net1714),
    .A1(net1593));
 sg13g2_nor3_1 _09124_ (.A(_03172_),
    .B(_03174_),
    .C(_03175_),
    .Y(_03176_));
 sg13g2_o21ai_1 _09125_ (.B1(_03172_),
    .Y(_03177_),
    .A1(_03174_),
    .A2(_03175_));
 sg13g2_nor2b_1 _09126_ (.A(_03176_),
    .B_N(_03177_),
    .Y(_03178_));
 sg13g2_nand2_1 _09127_ (.Y(_03179_),
    .A(_03171_),
    .B(_03178_));
 sg13g2_xnor2_1 _09128_ (.Y(_03180_),
    .A(_03171_),
    .B(_03178_));
 sg13g2_xnor2_1 _09129_ (.Y(_03181_),
    .A(_03170_),
    .B(_03180_));
 sg13g2_nand2b_1 _09130_ (.Y(_03182_),
    .B(_03162_),
    .A_N(_03181_));
 sg13g2_xor2_1 _09131_ (.B(_03181_),
    .A(_03162_),
    .X(_03183_));
 sg13g2_xnor2_1 _09132_ (.Y(_03184_),
    .A(_03161_),
    .B(_03183_));
 sg13g2_o21ai_1 _09133_ (.B1(_03105_),
    .Y(_03185_),
    .A1(_03084_),
    .A2(_03106_));
 sg13g2_o21ai_1 _09134_ (.B1(_03079_),
    .Y(_03186_),
    .A1(_03076_),
    .A2(_03080_));
 sg13g2_inv_1 _09135_ (.Y(_03187_),
    .A(_03186_));
 sg13g2_o21ai_1 _09136_ (.B1(_03088_),
    .Y(_03188_),
    .A1(_03086_),
    .A2(_03089_));
 sg13g2_nand2_1 _09137_ (.Y(_03189_),
    .A(net1598),
    .B(net1708));
 sg13g2_nand2_1 _09138_ (.Y(_03190_),
    .A(net1605),
    .B(net1696));
 sg13g2_nand2_1 _09139_ (.Y(_03191_),
    .A(net1608),
    .B(net1696));
 sg13g2_or2_1 _09140_ (.X(_03192_),
    .B(_03190_),
    .A(_03078_));
 sg13g2_xnor2_1 _09141_ (.Y(_03193_),
    .A(_03077_),
    .B(_03191_));
 sg13g2_xor2_1 _09142_ (.B(_03193_),
    .A(_03189_),
    .X(_03194_));
 sg13g2_nand2_1 _09143_ (.Y(_03195_),
    .A(_03188_),
    .B(_03194_));
 sg13g2_xnor2_1 _09144_ (.Y(_03196_),
    .A(_03188_),
    .B(_03194_));
 sg13g2_xnor2_1 _09145_ (.Y(_03197_),
    .A(_03187_),
    .B(_03196_));
 sg13g2_o21ai_1 _09146_ (.B1(_03100_),
    .Y(_03198_),
    .A1(_03091_),
    .A2(_03101_));
 sg13g2_nand2_1 _09147_ (.Y(_03199_),
    .A(net1612),
    .B(net1689));
 sg13g2_nand2_1 _09148_ (.Y(_03200_),
    .A(net1618),
    .B(net1680));
 sg13g2_and4_1 _09149_ (.A(net1619),
    .B(net1624),
    .C(net1680),
    .D(net1686),
    .X(_03201_));
 sg13g2_a22oi_1 _09150_ (.Y(_03202_),
    .B1(net1686),
    .B2(net1619),
    .A2(net1680),
    .A1(net1623));
 sg13g2_nor3_1 _09151_ (.A(_03199_),
    .B(_03201_),
    .C(_03202_),
    .Y(_03203_));
 sg13g2_o21ai_1 _09152_ (.B1(_03199_),
    .Y(_03204_),
    .A1(_03201_),
    .A2(_03202_));
 sg13g2_nand2b_1 _09153_ (.Y(_03205_),
    .B(_03204_),
    .A_N(_03203_));
 sg13g2_o21ai_1 _09154_ (.B1(_03095_),
    .Y(_03206_),
    .A1(_03093_),
    .A2(_03096_));
 sg13g2_nand2_1 _09155_ (.Y(_03207_),
    .A(net1631),
    .B(net1676));
 sg13g2_and4_1 _09156_ (.A(net1636),
    .B(net1646),
    .C(net1668),
    .D(net1672),
    .X(_03208_));
 sg13g2_nand4_1 _09157_ (.B(net1647),
    .C(net1668),
    .A(net1637),
    .Y(_03209_),
    .D(net1672));
 sg13g2_a22oi_1 _09158_ (.Y(_03210_),
    .B1(net1671),
    .B2(net1637),
    .A2(net1668),
    .A1(net1646));
 sg13g2_or3_1 _09159_ (.A(_03207_),
    .B(_03208_),
    .C(_03210_),
    .X(_03211_));
 sg13g2_o21ai_1 _09160_ (.B1(_03207_),
    .Y(_03212_),
    .A1(_03208_),
    .A2(_03210_));
 sg13g2_and3_1 _09161_ (.X(_03213_),
    .A(_03206_),
    .B(_03211_),
    .C(_03212_));
 sg13g2_nand3_1 _09162_ (.B(_03211_),
    .C(_03212_),
    .A(_03206_),
    .Y(_03214_));
 sg13g2_a21oi_1 _09163_ (.A1(_03211_),
    .A2(_03212_),
    .Y(_03215_),
    .B1(_03206_));
 sg13g2_or3_1 _09164_ (.A(_03205_),
    .B(_03213_),
    .C(_03215_),
    .X(_03216_));
 sg13g2_o21ai_1 _09165_ (.B1(_03205_),
    .Y(_03217_),
    .A1(_03213_),
    .A2(_03215_));
 sg13g2_and3_1 _09166_ (.X(_03218_),
    .A(_03198_),
    .B(_03216_),
    .C(_03217_));
 sg13g2_nand3_1 _09167_ (.B(_03216_),
    .C(_03217_),
    .A(_03198_),
    .Y(_03219_));
 sg13g2_a21oi_1 _09168_ (.A1(_03216_),
    .A2(_03217_),
    .Y(_03220_),
    .B1(_03198_));
 sg13g2_or3_1 _09169_ (.A(_03197_),
    .B(_03218_),
    .C(_03220_),
    .X(_03221_));
 sg13g2_o21ai_1 _09170_ (.B1(_03197_),
    .Y(_03222_),
    .A1(_03218_),
    .A2(_03220_));
 sg13g2_and3_1 _09171_ (.X(_03223_),
    .A(_03185_),
    .B(_03221_),
    .C(_03222_));
 sg13g2_nand3_1 _09172_ (.B(_03221_),
    .C(_03222_),
    .A(_03185_),
    .Y(_03224_));
 sg13g2_a21oi_1 _09173_ (.A1(_03221_),
    .A2(_03222_),
    .Y(_03225_),
    .B1(_03185_));
 sg13g2_or3_1 _09174_ (.A(_03184_),
    .B(_03223_),
    .C(_03225_),
    .X(_03226_));
 sg13g2_o21ai_1 _09175_ (.B1(_03184_),
    .Y(_03227_),
    .A1(_03223_),
    .A2(_03225_));
 sg13g2_and3_1 _09176_ (.X(_03228_),
    .A(_03159_),
    .B(_03226_),
    .C(_03227_));
 sg13g2_nand3_1 _09177_ (.B(_03226_),
    .C(_03227_),
    .A(_03159_),
    .Y(_03229_));
 sg13g2_a21oi_1 _09178_ (.A1(_03226_),
    .A2(_03227_),
    .Y(_03230_),
    .B1(_03159_));
 sg13g2_nor2_1 _09179_ (.A(_03228_),
    .B(_03230_),
    .Y(_03231_));
 sg13g2_a21o_1 _09180_ (.A2(_03134_),
    .A1(_03122_),
    .B1(_03136_),
    .X(_03232_));
 sg13g2_o21ai_1 _09181_ (.B1(_03069_),
    .Y(_03233_),
    .A1(_03051_),
    .A2(_03070_));
 sg13g2_nand2_1 _09182_ (.Y(_03234_),
    .A(net1499),
    .B(net1556));
 sg13g2_nand2_1 _09183_ (.Y(_03235_),
    .A(net1501),
    .B(net1544));
 sg13g2_nand2_1 _09184_ (.Y(_03236_),
    .A(net1505),
    .B(net1547));
 sg13g2_xor2_1 _09185_ (.B(_03236_),
    .A(_03120_),
    .X(_03237_));
 sg13g2_nand2b_1 _09186_ (.Y(_03238_),
    .B(_03237_),
    .A_N(_03234_));
 sg13g2_xnor2_1 _09187_ (.Y(_03239_),
    .A(_03234_),
    .B(_03237_));
 sg13g2_nand2_1 _09188_ (.Y(_03240_),
    .A(_03121_),
    .B(_03239_));
 sg13g2_xor2_1 _09189_ (.B(_03239_),
    .A(_03121_),
    .X(_03241_));
 sg13g2_inv_1 _09190_ (.Y(_03242_),
    .A(_03241_));
 sg13g2_o21ai_1 _09191_ (.B1(_03132_),
    .Y(_03243_),
    .A1(_03124_),
    .A2(_03133_));
 sg13g2_o21ai_1 _09192_ (.B1(_03129_),
    .Y(_03244_),
    .A1(_03126_),
    .A2(_03130_));
 sg13g2_inv_1 _09193_ (.Y(_03245_),
    .A(_03244_));
 sg13g2_o21ai_1 _09194_ (.B1(_03055_),
    .Y(_03246_),
    .A1(_03053_),
    .A2(_03056_));
 sg13g2_nand2_1 _09195_ (.Y(_03247_),
    .A(net1509),
    .B(net1537));
 sg13g2_nand2_1 _09196_ (.Y(_03248_),
    .A(net1511),
    .B(net1527));
 sg13g2_nand2_2 _09197_ (.Y(_03249_),
    .A(net1563),
    .B(net1530));
 sg13g2_or2_1 _09198_ (.X(_03250_),
    .B(_03248_),
    .A(_03128_));
 sg13g2_xnor2_1 _09199_ (.Y(_03251_),
    .A(_03127_),
    .B(_03249_));
 sg13g2_xor2_1 _09200_ (.B(_03251_),
    .A(_03247_),
    .X(_03252_));
 sg13g2_nand2_1 _09201_ (.Y(_03253_),
    .A(_03246_),
    .B(_03252_));
 sg13g2_xnor2_1 _09202_ (.Y(_03254_),
    .A(_03246_),
    .B(_03252_));
 sg13g2_xnor2_1 _09203_ (.Y(_03255_),
    .A(_03245_),
    .B(_03254_));
 sg13g2_nand2b_1 _09204_ (.Y(_03256_),
    .B(_03243_),
    .A_N(_03255_));
 sg13g2_xor2_1 _09205_ (.B(_03255_),
    .A(_03243_),
    .X(_03257_));
 sg13g2_xnor2_1 _09206_ (.Y(_03258_),
    .A(_03242_),
    .B(_03257_));
 sg13g2_nor2b_1 _09207_ (.A(_03258_),
    .B_N(_03233_),
    .Y(_03259_));
 sg13g2_xor2_1 _09208_ (.B(_03258_),
    .A(_03233_),
    .X(_03260_));
 sg13g2_nor2b_1 _09209_ (.A(_03260_),
    .B_N(_03232_),
    .Y(_03261_));
 sg13g2_xor2_1 _09210_ (.B(_03260_),
    .A(_03232_),
    .X(_03262_));
 sg13g2_xnor2_1 _09211_ (.Y(_03263_),
    .A(_03231_),
    .B(_03262_));
 sg13g2_nand2_1 _09212_ (.Y(_03264_),
    .A(_03158_),
    .B(_03263_));
 sg13g2_xnor2_1 _09213_ (.Y(_03265_),
    .A(_03158_),
    .B(_03263_));
 sg13g2_xnor2_1 _09214_ (.Y(_03266_),
    .A(_03157_),
    .B(_03265_));
 sg13g2_o21ai_1 _09215_ (.B1(_03144_),
    .Y(_03267_),
    .A1(_03047_),
    .A2(_03145_));
 sg13g2_nand2b_1 _09216_ (.Y(_03268_),
    .B(_03267_),
    .A_N(_03266_));
 sg13g2_xnor2_1 _09217_ (.Y(_03269_),
    .A(_03266_),
    .B(_03267_));
 sg13g2_nor2b_1 _09218_ (.A(_03148_),
    .B_N(_03269_),
    .Y(_03270_));
 sg13g2_xor2_1 _09219_ (.B(_03269_),
    .A(_03148_),
    .X(_03271_));
 sg13g2_inv_1 _09220_ (.Y(_03272_),
    .A(_03271_));
 sg13g2_or3_1 _09221_ (.A(_03031_),
    .B(_03149_),
    .C(_03271_),
    .X(_03273_));
 sg13g2_xor2_1 _09222_ (.B(_03271_),
    .A(_03150_),
    .X(_03274_));
 sg13g2_nand2_1 _09223_ (.Y(_03275_),
    .A(_03037_),
    .B(_03152_));
 sg13g2_a21oi_1 _09224_ (.A1(_03033_),
    .A2(_03035_),
    .Y(_03276_),
    .B1(_03151_));
 sg13g2_inv_1 _09225_ (.Y(_03277_),
    .A(_03276_));
 sg13g2_a21oi_1 _09226_ (.A1(_03037_),
    .A2(_03152_),
    .Y(_03278_),
    .B1(_03276_));
 sg13g2_nor2_1 _09227_ (.A(_03040_),
    .B(_03276_),
    .Y(_03279_));
 sg13g2_a21o_1 _09228_ (.A2(_03279_),
    .A1(_03039_),
    .B1(_03278_),
    .X(_03280_));
 sg13g2_a221oi_1 _09229_ (.B2(_03039_),
    .C1(_03274_),
    .B1(_03279_),
    .A1(_03275_),
    .Y(_03281_),
    .A2(_03277_));
 sg13g2_xnor2_1 _09230_ (.Y(_03282_),
    .A(_03274_),
    .B(_03280_));
 sg13g2_inv_1 _09231_ (.Y(_03283_),
    .A(_03282_));
 sg13g2_o21ai_1 _09232_ (.B1(net1751),
    .Y(_03284_),
    .A1(net1469),
    .A2(net638));
 sg13g2_a21oi_1 _09233_ (.A1(net1469),
    .A2(_03282_),
    .Y(_00320_),
    .B1(_03284_));
 sg13g2_a21oi_1 _09234_ (.A1(_03150_),
    .A2(_03272_),
    .Y(_03285_),
    .B1(_03281_));
 sg13g2_nor2_1 _09235_ (.A(_03259_),
    .B(_03261_),
    .Y(_03286_));
 sg13g2_nor2_1 _09236_ (.A(_03240_),
    .B(_03286_),
    .Y(_03287_));
 sg13g2_inv_1 _09237_ (.Y(_03288_),
    .A(_03287_));
 sg13g2_xnor2_1 _09238_ (.Y(_03289_),
    .A(_03240_),
    .B(_03286_));
 sg13g2_o21ai_1 _09239_ (.B1(_03229_),
    .Y(_03290_),
    .A1(_03230_),
    .A2(_03262_));
 sg13g2_o21ai_1 _09240_ (.B1(_03256_),
    .Y(_03291_),
    .A1(_03242_),
    .A2(_03257_));
 sg13g2_inv_1 _09241_ (.Y(_03292_),
    .A(_03291_));
 sg13g2_o21ai_1 _09242_ (.B1(_03182_),
    .Y(_03293_),
    .A1(_03161_),
    .A2(_03183_));
 sg13g2_nand2_1 _09243_ (.Y(_03294_),
    .A(net1495),
    .B(net1556));
 sg13g2_o21ai_1 _09244_ (.B1(_03238_),
    .Y(_03295_),
    .A1(_03120_),
    .A2(_03236_));
 sg13g2_nand2_1 _09245_ (.Y(_03296_),
    .A(net1499),
    .B(net1549));
 sg13g2_nand2_2 _09246_ (.Y(_03297_),
    .A(net1505),
    .B(net1542));
 sg13g2_or2_1 _09247_ (.X(_03298_),
    .B(_03297_),
    .A(_03235_));
 sg13g2_xnor2_1 _09248_ (.Y(_03299_),
    .A(_03235_),
    .B(_03297_));
 sg13g2_xor2_1 _09249_ (.B(_03299_),
    .A(_03296_),
    .X(_03300_));
 sg13g2_nand2_1 _09250_ (.Y(_03301_),
    .A(_03295_),
    .B(_03300_));
 sg13g2_xnor2_1 _09251_ (.Y(_03302_),
    .A(_03295_),
    .B(_03300_));
 sg13g2_xor2_1 _09252_ (.B(_03302_),
    .A(_03294_),
    .X(_03303_));
 sg13g2_inv_1 _09253_ (.Y(_03304_),
    .A(_03303_));
 sg13g2_o21ai_1 _09254_ (.B1(_03253_),
    .Y(_03305_),
    .A1(_03245_),
    .A2(_03254_));
 sg13g2_o21ai_1 _09255_ (.B1(_03250_),
    .Y(_03306_),
    .A1(_03247_),
    .A2(_03251_));
 sg13g2_inv_1 _09256_ (.Y(_03307_),
    .A(_03306_));
 sg13g2_o21ai_1 _09257_ (.B1(_03166_),
    .Y(_03308_),
    .A1(_03163_),
    .A2(_03167_));
 sg13g2_nand2_1 _09258_ (.Y(_03309_),
    .A(net1509),
    .B(net1532));
 sg13g2_nand2_1 _09259_ (.Y(_03310_),
    .A(net1510),
    .B(net1520));
 sg13g2_nand2_1 _09260_ (.Y(_03311_),
    .A(net1562),
    .B(net1520));
 sg13g2_or2_1 _09261_ (.X(_03312_),
    .B(_03310_),
    .A(_03249_));
 sg13g2_xnor2_1 _09262_ (.Y(_03313_),
    .A(_03248_),
    .B(_03311_));
 sg13g2_xor2_1 _09263_ (.B(_03313_),
    .A(_03309_),
    .X(_03314_));
 sg13g2_nand2_1 _09264_ (.Y(_03315_),
    .A(_03308_),
    .B(_03314_));
 sg13g2_xnor2_1 _09265_ (.Y(_03316_),
    .A(_03308_),
    .B(_03314_));
 sg13g2_xnor2_1 _09266_ (.Y(_03317_),
    .A(_03307_),
    .B(_03316_));
 sg13g2_nand2b_1 _09267_ (.Y(_03318_),
    .B(_03305_),
    .A_N(_03317_));
 sg13g2_xor2_1 _09268_ (.B(_03317_),
    .A(_03305_),
    .X(_03319_));
 sg13g2_xor2_1 _09269_ (.B(_03319_),
    .A(_03303_),
    .X(_03320_));
 sg13g2_nand2b_1 _09270_ (.Y(_03321_),
    .B(_03293_),
    .A_N(_03320_));
 sg13g2_xor2_1 _09271_ (.B(_03320_),
    .A(_03293_),
    .X(_03322_));
 sg13g2_xnor2_1 _09272_ (.Y(_03323_),
    .A(_03292_),
    .B(_03322_));
 sg13g2_o21ai_1 _09273_ (.B1(_03224_),
    .Y(_03324_),
    .A1(_03184_),
    .A2(_03225_));
 sg13g2_o21ai_1 _09274_ (.B1(_03179_),
    .Y(_03325_),
    .A1(_03170_),
    .A2(_03180_));
 sg13g2_inv_1 _09275_ (.Y(_03326_),
    .A(_03325_));
 sg13g2_o21ai_1 _09276_ (.B1(_03195_),
    .Y(_03327_),
    .A1(_03187_),
    .A2(_03196_));
 sg13g2_nand2_1 _09277_ (.Y(_03328_),
    .A(net1566),
    .B(net1514));
 sg13g2_nand2_1 _09278_ (.Y(_03329_),
    .A(net1574),
    .B(net1726));
 sg13g2_or2_1 _09279_ (.X(_03330_),
    .B(_03329_),
    .A(_03164_));
 sg13g2_and2_1 _09280_ (.A(_03164_),
    .B(_03329_),
    .X(_03331_));
 sg13g2_xnor2_1 _09281_ (.Y(_03332_),
    .A(_03164_),
    .B(_03329_));
 sg13g2_xnor2_1 _09282_ (.Y(_03333_),
    .A(_03328_),
    .B(_03332_));
 sg13g2_or2_1 _09283_ (.X(_03334_),
    .B(_03176_),
    .A(_03174_));
 sg13g2_nand2_1 _09284_ (.Y(_03335_),
    .A(net1580),
    .B(net1719));
 sg13g2_nand2_1 _09285_ (.Y(_03336_),
    .A(net1592),
    .B(net1708));
 sg13g2_or2_1 _09286_ (.X(_03337_),
    .B(_03336_),
    .A(_03173_));
 sg13g2_and2_1 _09287_ (.A(_03173_),
    .B(_03336_),
    .X(_03338_));
 sg13g2_xor2_1 _09288_ (.B(_03336_),
    .A(_03173_),
    .X(_03339_));
 sg13g2_xnor2_1 _09289_ (.Y(_03340_),
    .A(_03335_),
    .B(_03339_));
 sg13g2_nand2_1 _09290_ (.Y(_03341_),
    .A(_03334_),
    .B(_03340_));
 sg13g2_xnor2_1 _09291_ (.Y(_03342_),
    .A(_03334_),
    .B(_03340_));
 sg13g2_xor2_1 _09292_ (.B(_03342_),
    .A(_03333_),
    .X(_03343_));
 sg13g2_nand2_1 _09293_ (.Y(_03344_),
    .A(_03327_),
    .B(_03343_));
 sg13g2_xnor2_1 _09294_ (.Y(_03345_),
    .A(_03327_),
    .B(_03343_));
 sg13g2_xnor2_1 _09295_ (.Y(_03346_),
    .A(_03326_),
    .B(_03345_));
 sg13g2_o21ai_1 _09296_ (.B1(_03219_),
    .Y(_03347_),
    .A1(_03197_),
    .A2(_03220_));
 sg13g2_o21ai_1 _09297_ (.B1(_03192_),
    .Y(_03348_),
    .A1(_03189_),
    .A2(_03193_));
 sg13g2_inv_1 _09298_ (.Y(_03349_),
    .A(_03348_));
 sg13g2_or2_1 _09299_ (.X(_03350_),
    .B(_03203_),
    .A(_03201_));
 sg13g2_nand2_1 _09300_ (.Y(_03351_),
    .A(net1598),
    .B(net1701));
 sg13g2_nand2_1 _09301_ (.Y(_03352_),
    .A(net1603),
    .B(net1691));
 sg13g2_nand2_1 _09302_ (.Y(_03353_),
    .A(net1607),
    .B(net1691));
 sg13g2_or2_1 _09303_ (.X(_03354_),
    .B(_03352_),
    .A(_03191_));
 sg13g2_xnor2_1 _09304_ (.Y(_03355_),
    .A(_03190_),
    .B(_03353_));
 sg13g2_xor2_1 _09305_ (.B(_03355_),
    .A(_03351_),
    .X(_03356_));
 sg13g2_nand2_1 _09306_ (.Y(_03357_),
    .A(_03350_),
    .B(_03356_));
 sg13g2_xnor2_1 _09307_ (.Y(_03358_),
    .A(_03350_),
    .B(_03356_));
 sg13g2_xnor2_1 _09308_ (.Y(_03359_),
    .A(_03349_),
    .B(_03358_));
 sg13g2_o21ai_1 _09309_ (.B1(_03214_),
    .Y(_03360_),
    .A1(_03205_),
    .A2(_03215_));
 sg13g2_nand2_1 _09310_ (.Y(_03361_),
    .A(net1612),
    .B(net1687));
 sg13g2_nand2_1 _09311_ (.Y(_03362_),
    .A(net1623),
    .B(net1676));
 sg13g2_or2_1 _09312_ (.X(_03363_),
    .B(_03362_),
    .A(_03200_));
 sg13g2_and2_1 _09313_ (.A(_03200_),
    .B(_03362_),
    .X(_03364_));
 sg13g2_xnor2_1 _09314_ (.Y(_03365_),
    .A(_03200_),
    .B(_03362_));
 sg13g2_xnor2_1 _09315_ (.Y(_03366_),
    .A(_03361_),
    .B(_03365_));
 sg13g2_o21ai_1 _09316_ (.B1(_03209_),
    .Y(_03367_),
    .A1(_03207_),
    .A2(_03210_));
 sg13g2_nand2_1 _09317_ (.Y(_03368_),
    .A(net1631),
    .B(net1672));
 sg13g2_and4_1 _09318_ (.A(net1636),
    .B(net1647),
    .C(net1664),
    .D(net1668),
    .X(_03369_));
 sg13g2_nand4_1 _09319_ (.B(net1646),
    .C(net1664),
    .A(net1636),
    .Y(_03370_),
    .D(net1668));
 sg13g2_a22oi_1 _09320_ (.Y(_03371_),
    .B1(net1669),
    .B2(net1637),
    .A2(net1664),
    .A1(net1647));
 sg13g2_or3_1 _09321_ (.A(_03368_),
    .B(_03369_),
    .C(_03371_),
    .X(_03372_));
 sg13g2_o21ai_1 _09322_ (.B1(_03368_),
    .Y(_03373_),
    .A1(_03369_),
    .A2(_03371_));
 sg13g2_and3_1 _09323_ (.X(_03374_),
    .A(_03367_),
    .B(_03372_),
    .C(_03373_));
 sg13g2_nand3_1 _09324_ (.B(_03372_),
    .C(_03373_),
    .A(_03367_),
    .Y(_03375_));
 sg13g2_a21oi_1 _09325_ (.A1(_03372_),
    .A2(_03373_),
    .Y(_03376_),
    .B1(_03367_));
 sg13g2_or3_1 _09326_ (.A(_03366_),
    .B(_03374_),
    .C(_03376_),
    .X(_03377_));
 sg13g2_o21ai_1 _09327_ (.B1(_03366_),
    .Y(_03378_),
    .A1(_03374_),
    .A2(_03376_));
 sg13g2_and3_1 _09328_ (.X(_03379_),
    .A(_03360_),
    .B(_03377_),
    .C(_03378_));
 sg13g2_nand3_1 _09329_ (.B(_03377_),
    .C(_03378_),
    .A(_03360_),
    .Y(_03380_));
 sg13g2_a21oi_1 _09330_ (.A1(_03377_),
    .A2(_03378_),
    .Y(_03381_),
    .B1(_03360_));
 sg13g2_or3_1 _09331_ (.A(_03359_),
    .B(_03379_),
    .C(_03381_),
    .X(_03382_));
 sg13g2_o21ai_1 _09332_ (.B1(_03359_),
    .Y(_03383_),
    .A1(_03379_),
    .A2(_03381_));
 sg13g2_and3_1 _09333_ (.X(_03384_),
    .A(_03347_),
    .B(_03382_),
    .C(_03383_));
 sg13g2_nand3_1 _09334_ (.B(_03382_),
    .C(_03383_),
    .A(_03347_),
    .Y(_03385_));
 sg13g2_a21oi_1 _09335_ (.A1(_03382_),
    .A2(_03383_),
    .Y(_03386_),
    .B1(_03347_));
 sg13g2_or3_1 _09336_ (.A(_03346_),
    .B(_03384_),
    .C(_03386_),
    .X(_03387_));
 sg13g2_o21ai_1 _09337_ (.B1(_03346_),
    .Y(_03388_),
    .A1(_03384_),
    .A2(_03386_));
 sg13g2_and3_1 _09338_ (.X(_03389_),
    .A(_03324_),
    .B(_03387_),
    .C(_03388_));
 sg13g2_nand3_1 _09339_ (.B(_03387_),
    .C(_03388_),
    .A(_03324_),
    .Y(_03390_));
 sg13g2_a21oi_1 _09340_ (.A1(_03387_),
    .A2(_03388_),
    .Y(_03391_),
    .B1(_03324_));
 sg13g2_or3_1 _09341_ (.A(_03323_),
    .B(_03389_),
    .C(_03391_),
    .X(_03392_));
 sg13g2_o21ai_1 _09342_ (.B1(_03323_),
    .Y(_03393_),
    .A1(_03389_),
    .A2(_03391_));
 sg13g2_nand3_1 _09343_ (.B(_03392_),
    .C(_03393_),
    .A(_03290_),
    .Y(_03394_));
 sg13g2_a21oi_1 _09344_ (.A1(_03392_),
    .A2(_03393_),
    .Y(_03395_),
    .B1(_03290_));
 sg13g2_a21o_1 _09345_ (.A2(_03393_),
    .A1(_03392_),
    .B1(_03290_),
    .X(_03396_));
 sg13g2_nand2_1 _09346_ (.Y(_03397_),
    .A(_03394_),
    .B(_03396_));
 sg13g2_xor2_1 _09347_ (.B(_03397_),
    .A(_03289_),
    .X(_03398_));
 sg13g2_o21ai_1 _09348_ (.B1(_03264_),
    .Y(_03399_),
    .A1(_03157_),
    .A2(_03265_));
 sg13g2_nand2_1 _09349_ (.Y(_03400_),
    .A(_03398_),
    .B(_03399_));
 sg13g2_xor2_1 _09350_ (.B(_03399_),
    .A(_03398_),
    .X(_03401_));
 sg13g2_nor2b_1 _09351_ (.A(_03268_),
    .B_N(_03401_),
    .Y(_03402_));
 sg13g2_xnor2_1 _09352_ (.Y(_03403_),
    .A(_03268_),
    .B(_03401_));
 sg13g2_inv_1 _09353_ (.Y(_03404_),
    .A(_03403_));
 sg13g2_nand2_1 _09354_ (.Y(_03405_),
    .A(_03270_),
    .B(_03403_));
 sg13g2_xnor2_1 _09355_ (.Y(_03406_),
    .A(_03270_),
    .B(_03403_));
 sg13g2_inv_1 _09356_ (.Y(_03407_),
    .A(_03406_));
 sg13g2_xnor2_1 _09357_ (.Y(_03408_),
    .A(_03285_),
    .B(_03406_));
 sg13g2_o21ai_1 _09358_ (.B1(net1753),
    .Y(_03409_),
    .A1(net1469),
    .A2(net614));
 sg13g2_a21oi_1 _09359_ (.A1(net1469),
    .A2(_03408_),
    .Y(_00321_),
    .B1(_03409_));
 sg13g2_o21ai_1 _09360_ (.B1(_03394_),
    .Y(_03410_),
    .A1(_03289_),
    .A2(_03395_));
 sg13g2_o21ai_1 _09361_ (.B1(_03321_),
    .Y(_03411_),
    .A1(_03292_),
    .A2(_03322_));
 sg13g2_o21ai_1 _09362_ (.B1(_03301_),
    .Y(_03412_),
    .A1(_03294_),
    .A2(_03302_));
 sg13g2_nand2_1 _09363_ (.Y(_03413_),
    .A(_03411_),
    .B(_03412_));
 sg13g2_xor2_1 _09364_ (.B(_03412_),
    .A(_03411_),
    .X(_03414_));
 sg13g2_o21ai_1 _09365_ (.B1(_03390_),
    .Y(_03415_),
    .A1(_03323_),
    .A2(_03391_));
 sg13g2_o21ai_1 _09366_ (.B1(_03318_),
    .Y(_03416_),
    .A1(_03304_),
    .A2(_03319_));
 sg13g2_o21ai_1 _09367_ (.B1(_03344_),
    .Y(_03417_),
    .A1(_03326_),
    .A2(_03345_));
 sg13g2_a22oi_1 _09368_ (.Y(_03418_),
    .B1(net1558),
    .B2(net1491),
    .A2(net1549),
    .A1(net1495));
 sg13g2_nand4_1 _09369_ (.B(net1495),
    .C(net1550),
    .A(net1491),
    .Y(_03419_),
    .D(net1558));
 sg13g2_nor2b_1 _09370_ (.A(_03418_),
    .B_N(_03419_),
    .Y(_03420_));
 sg13g2_and2_1 _09371_ (.A(net1499),
    .B(net1544),
    .X(_03421_));
 sg13g2_nand2_2 _09372_ (.Y(_03422_),
    .A(net1501),
    .B(net1532));
 sg13g2_nor2_1 _09373_ (.A(_03297_),
    .B(_03422_),
    .Y(_03423_));
 sg13g2_a22oi_1 _09374_ (.Y(_03424_),
    .B1(net1537),
    .B2(net1501),
    .A2(net1532),
    .A1(net1505));
 sg13g2_nor2_1 _09375_ (.A(_03423_),
    .B(_03424_),
    .Y(_03425_));
 sg13g2_xor2_1 _09376_ (.B(_03425_),
    .A(_03421_),
    .X(_03426_));
 sg13g2_o21ai_1 _09377_ (.B1(_03298_),
    .Y(_03427_),
    .A1(_03296_),
    .A2(_03299_));
 sg13g2_nand2_1 _09378_ (.Y(_03428_),
    .A(_03426_),
    .B(_03427_));
 sg13g2_xor2_1 _09379_ (.B(_03427_),
    .A(_03426_),
    .X(_03429_));
 sg13g2_xnor2_1 _09380_ (.Y(_03430_),
    .A(_03420_),
    .B(_03429_));
 sg13g2_o21ai_1 _09381_ (.B1(_03315_),
    .Y(_03431_),
    .A1(_03307_),
    .A2(_03316_));
 sg13g2_o21ai_1 _09382_ (.B1(_03312_),
    .Y(_03432_),
    .A1(_03309_),
    .A2(_03313_));
 sg13g2_inv_1 _09383_ (.Y(_03433_),
    .A(_03432_));
 sg13g2_o21ai_1 _09384_ (.B1(_03330_),
    .Y(_03434_),
    .A1(_03328_),
    .A2(_03331_));
 sg13g2_nand2_1 _09385_ (.Y(_03435_),
    .A(net1508),
    .B(net1530));
 sg13g2_nand2_2 _09386_ (.Y(_03436_),
    .A(net1510),
    .B(\cordic_inst.MUX_cordic_state$write_1__VAL_1[63] ));
 sg13g2_nand2_1 _09387_ (.Y(_03437_),
    .A(net1562),
    .B(net1515));
 sg13g2_or2_1 _09388_ (.X(_03438_),
    .B(_03436_),
    .A(_03311_));
 sg13g2_xnor2_1 _09389_ (.Y(_03439_),
    .A(_03310_),
    .B(_03437_));
 sg13g2_xor2_1 _09390_ (.B(_03439_),
    .A(_03435_),
    .X(_03440_));
 sg13g2_nand2_1 _09391_ (.Y(_03441_),
    .A(_03434_),
    .B(_03440_));
 sg13g2_xnor2_1 _09392_ (.Y(_03442_),
    .A(_03434_),
    .B(_03440_));
 sg13g2_xnor2_1 _09393_ (.Y(_03443_),
    .A(_03433_),
    .B(_03442_));
 sg13g2_nand2b_1 _09394_ (.Y(_03444_),
    .B(_03431_),
    .A_N(_03443_));
 sg13g2_xor2_1 _09395_ (.B(_03443_),
    .A(_03431_),
    .X(_03445_));
 sg13g2_xor2_1 _09396_ (.B(_03445_),
    .A(_03430_),
    .X(_03446_));
 sg13g2_nand2_1 _09397_ (.Y(_03447_),
    .A(_03417_),
    .B(_03446_));
 sg13g2_xnor2_1 _09398_ (.Y(_03448_),
    .A(_03417_),
    .B(_03446_));
 sg13g2_nand2b_1 _09399_ (.Y(_03449_),
    .B(_03416_),
    .A_N(_03448_));
 sg13g2_xor2_1 _09400_ (.B(_03448_),
    .A(_03416_),
    .X(_03450_));
 sg13g2_o21ai_1 _09401_ (.B1(_03385_),
    .Y(_03451_),
    .A1(_03346_),
    .A2(_03386_));
 sg13g2_o21ai_1 _09402_ (.B1(_03341_),
    .Y(_03452_),
    .A1(_03333_),
    .A2(_03342_));
 sg13g2_inv_1 _09403_ (.Y(_03453_),
    .A(_03452_));
 sg13g2_o21ai_1 _09404_ (.B1(_03357_),
    .Y(_03454_),
    .A1(_03349_),
    .A2(_03358_));
 sg13g2_nand2_1 _09405_ (.Y(_03455_),
    .A(net1566),
    .B(net1728));
 sg13g2_nand2_1 _09406_ (.Y(_03456_),
    .A(net1570),
    .B(net1715));
 sg13g2_and4_1 _09407_ (.A(net1571),
    .B(net1574),
    .C(net1719),
    .D(net1721),
    .X(_03457_));
 sg13g2_a22oi_1 _09408_ (.Y(_03458_),
    .B1(net1721),
    .B2(net1570),
    .A2(net1719),
    .A1(net1574));
 sg13g2_nor3_1 _09409_ (.A(_03455_),
    .B(_03457_),
    .C(_03458_),
    .Y(_03459_));
 sg13g2_o21ai_1 _09410_ (.B1(_03455_),
    .Y(_03460_),
    .A1(_03457_),
    .A2(_03458_));
 sg13g2_nor2b_1 _09411_ (.A(_03459_),
    .B_N(_03460_),
    .Y(_03461_));
 sg13g2_inv_1 _09412_ (.Y(_03462_),
    .A(_03461_));
 sg13g2_o21ai_1 _09413_ (.B1(_03337_),
    .Y(_03463_),
    .A1(_03335_),
    .A2(_03338_));
 sg13g2_nand2_1 _09414_ (.Y(_03464_),
    .A(net1580),
    .B(net1710));
 sg13g2_nand2_1 _09415_ (.Y(_03465_),
    .A(net1585),
    .B(net1701));
 sg13g2_and4_1 _09416_ (.A(net1585),
    .B(net1592),
    .C(net1701),
    .D(net1704),
    .X(_03466_));
 sg13g2_a22oi_1 _09417_ (.Y(_03467_),
    .B1(net1704),
    .B2(net1585),
    .A2(net1701),
    .A1(net1592));
 sg13g2_nor3_1 _09418_ (.A(_03464_),
    .B(_03466_),
    .C(_03467_),
    .Y(_03468_));
 sg13g2_o21ai_1 _09419_ (.B1(_03464_),
    .Y(_03469_),
    .A1(_03466_),
    .A2(_03467_));
 sg13g2_nor2b_1 _09420_ (.A(_03468_),
    .B_N(_03469_),
    .Y(_03470_));
 sg13g2_nand2_1 _09421_ (.Y(_03471_),
    .A(_03463_),
    .B(_03470_));
 sg13g2_xnor2_1 _09422_ (.Y(_03472_),
    .A(_03463_),
    .B(_03470_));
 sg13g2_xnor2_1 _09423_ (.Y(_03473_),
    .A(_03462_),
    .B(_03472_));
 sg13g2_nand2b_1 _09424_ (.Y(_03474_),
    .B(_03454_),
    .A_N(_03473_));
 sg13g2_xor2_1 _09425_ (.B(_03473_),
    .A(_03454_),
    .X(_03475_));
 sg13g2_xnor2_1 _09426_ (.Y(_03476_),
    .A(_03453_),
    .B(_03475_));
 sg13g2_o21ai_1 _09427_ (.B1(_03380_),
    .Y(_03477_),
    .A1(_03359_),
    .A2(_03381_));
 sg13g2_o21ai_1 _09428_ (.B1(_03354_),
    .Y(_03478_),
    .A1(_03351_),
    .A2(_03355_));
 sg13g2_inv_1 _09429_ (.Y(_03479_),
    .A(_03478_));
 sg13g2_o21ai_1 _09430_ (.B1(_03363_),
    .Y(_03480_),
    .A1(_03361_),
    .A2(_03364_));
 sg13g2_nand2_1 _09431_ (.Y(_03481_),
    .A(net1598),
    .B(net1696));
 sg13g2_nand2_1 _09432_ (.Y(_03482_),
    .A(net1603),
    .B(net1687));
 sg13g2_nand2_1 _09433_ (.Y(_03483_),
    .A(net1607),
    .B(net1687));
 sg13g2_or2_1 _09434_ (.X(_03484_),
    .B(_03482_),
    .A(_03353_));
 sg13g2_xnor2_1 _09435_ (.Y(_03485_),
    .A(_03352_),
    .B(_03483_));
 sg13g2_xor2_1 _09436_ (.B(_03485_),
    .A(_03481_),
    .X(_03486_));
 sg13g2_nand2_1 _09437_ (.Y(_03487_),
    .A(_03480_),
    .B(_03486_));
 sg13g2_xnor2_1 _09438_ (.Y(_03488_),
    .A(_03480_),
    .B(_03486_));
 sg13g2_xnor2_1 _09439_ (.Y(_03489_),
    .A(_03479_),
    .B(_03488_));
 sg13g2_o21ai_1 _09440_ (.B1(_03375_),
    .Y(_03490_),
    .A1(_03366_),
    .A2(_03376_));
 sg13g2_o21ai_1 _09441_ (.B1(_03370_),
    .Y(_03491_),
    .A1(_03368_),
    .A2(_03371_));
 sg13g2_nand2_1 _09442_ (.Y(_03492_),
    .A(net1631),
    .B(net1668));
 sg13g2_and4_1 _09443_ (.A(net1636),
    .B(net1646),
    .C(net1660),
    .D(net1663),
    .X(_03493_));
 sg13g2_nand4_1 _09444_ (.B(net1646),
    .C(net1660),
    .A(net1636),
    .Y(_03494_),
    .D(net1663));
 sg13g2_a22oi_1 _09445_ (.Y(_03495_),
    .B1(net1663),
    .B2(net1636),
    .A2(net1660),
    .A1(net1646));
 sg13g2_or3_1 _09446_ (.A(_03492_),
    .B(_03493_),
    .C(_03495_),
    .X(_03496_));
 sg13g2_o21ai_1 _09447_ (.B1(_03492_),
    .Y(_03497_),
    .A1(_03493_),
    .A2(_03495_));
 sg13g2_and3_1 _09448_ (.X(_03498_),
    .A(_03491_),
    .B(_03496_),
    .C(_03497_));
 sg13g2_nand3_1 _09449_ (.B(_03496_),
    .C(_03497_),
    .A(_03491_),
    .Y(_03499_));
 sg13g2_a21oi_1 _09450_ (.A1(_03496_),
    .A2(_03497_),
    .Y(_03500_),
    .B1(_03491_));
 sg13g2_nand2_1 _09451_ (.Y(_03501_),
    .A(net1612),
    .B(net1681));
 sg13g2_nand2_1 _09452_ (.Y(_03502_),
    .A(net1618),
    .B(net1671));
 sg13g2_and4_1 _09453_ (.A(net1618),
    .B(net1623),
    .C(net1671),
    .D(net1675),
    .X(_03503_));
 sg13g2_a22oi_1 _09454_ (.Y(_03504_),
    .B1(net1675),
    .B2(net1618),
    .A2(net1671),
    .A1(net1623));
 sg13g2_nor3_1 _09455_ (.A(_03501_),
    .B(_03503_),
    .C(_03504_),
    .Y(_03505_));
 sg13g2_o21ai_1 _09456_ (.B1(_03501_),
    .Y(_03506_),
    .A1(_03503_),
    .A2(_03504_));
 sg13g2_nand2b_1 _09457_ (.Y(_03507_),
    .B(_03506_),
    .A_N(_03505_));
 sg13g2_or3_1 _09458_ (.A(_03498_),
    .B(_03500_),
    .C(_03507_),
    .X(_03508_));
 sg13g2_o21ai_1 _09459_ (.B1(_03507_),
    .Y(_03509_),
    .A1(_03498_),
    .A2(_03500_));
 sg13g2_and3_1 _09460_ (.X(_03510_),
    .A(_03490_),
    .B(_03508_),
    .C(_03509_));
 sg13g2_nand3_1 _09461_ (.B(_03508_),
    .C(_03509_),
    .A(_03490_),
    .Y(_03511_));
 sg13g2_a21oi_1 _09462_ (.A1(_03508_),
    .A2(_03509_),
    .Y(_03512_),
    .B1(_03490_));
 sg13g2_or3_1 _09463_ (.A(_03489_),
    .B(_03510_),
    .C(_03512_),
    .X(_03513_));
 sg13g2_o21ai_1 _09464_ (.B1(_03489_),
    .Y(_03514_),
    .A1(_03510_),
    .A2(_03512_));
 sg13g2_and3_1 _09465_ (.X(_03515_),
    .A(_03477_),
    .B(_03513_),
    .C(_03514_));
 sg13g2_nand3_1 _09466_ (.B(_03513_),
    .C(_03514_),
    .A(_03477_),
    .Y(_03516_));
 sg13g2_a21oi_1 _09467_ (.A1(_03513_),
    .A2(_03514_),
    .Y(_03517_),
    .B1(_03477_));
 sg13g2_or3_1 _09468_ (.A(_03476_),
    .B(_03515_),
    .C(_03517_),
    .X(_03518_));
 sg13g2_o21ai_1 _09469_ (.B1(_03476_),
    .Y(_03519_),
    .A1(_03515_),
    .A2(_03517_));
 sg13g2_and3_1 _09470_ (.X(_03520_),
    .A(_03451_),
    .B(_03518_),
    .C(_03519_));
 sg13g2_nand3_1 _09471_ (.B(_03518_),
    .C(_03519_),
    .A(_03451_),
    .Y(_03521_));
 sg13g2_a21oi_1 _09472_ (.A1(_03518_),
    .A2(_03519_),
    .Y(_03522_),
    .B1(_03451_));
 sg13g2_or3_1 _09473_ (.A(_03450_),
    .B(_03520_),
    .C(_03522_),
    .X(_03523_));
 sg13g2_o21ai_1 _09474_ (.B1(_03450_),
    .Y(_03524_),
    .A1(_03520_),
    .A2(_03522_));
 sg13g2_and3_1 _09475_ (.X(_03525_),
    .A(_03415_),
    .B(_03523_),
    .C(_03524_));
 sg13g2_nand3_1 _09476_ (.B(_03523_),
    .C(_03524_),
    .A(_03415_),
    .Y(_03526_));
 sg13g2_a21o_1 _09477_ (.A2(_03524_),
    .A1(_03523_),
    .B1(_03415_),
    .X(_03527_));
 sg13g2_nand3_1 _09478_ (.B(_03526_),
    .C(_03527_),
    .A(_03414_),
    .Y(_03528_));
 sg13g2_a21o_1 _09479_ (.A2(_03527_),
    .A1(_03526_),
    .B1(_03414_),
    .X(_03529_));
 sg13g2_nand3_1 _09480_ (.B(_03528_),
    .C(_03529_),
    .A(_03410_),
    .Y(_03530_));
 sg13g2_a21oi_1 _09481_ (.A1(_03528_),
    .A2(_03529_),
    .Y(_03531_),
    .B1(_03410_));
 sg13g2_a21o_1 _09482_ (.A2(_03529_),
    .A1(_03528_),
    .B1(_03410_),
    .X(_03532_));
 sg13g2_a21oi_1 _09483_ (.A1(_03530_),
    .A2(_03532_),
    .Y(_03533_),
    .B1(_03287_));
 sg13g2_and3_2 _09484_ (.X(_03534_),
    .A(_03287_),
    .B(_03530_),
    .C(_03532_));
 sg13g2_nor3_1 _09485_ (.A(_03400_),
    .B(_03533_),
    .C(_03534_),
    .Y(_03535_));
 sg13g2_or3_1 _09486_ (.A(_03400_),
    .B(_03533_),
    .C(_03534_),
    .X(_03536_));
 sg13g2_o21ai_1 _09487_ (.B1(_03400_),
    .Y(_03537_),
    .A1(_03533_),
    .A2(_03534_));
 sg13g2_and3_1 _09488_ (.X(_03538_),
    .A(_03402_),
    .B(_03536_),
    .C(_03537_));
 sg13g2_nand3_1 _09489_ (.B(_03536_),
    .C(_03537_),
    .A(_03402_),
    .Y(_03539_));
 sg13g2_a21oi_1 _09490_ (.A1(_03536_),
    .A2(_03537_),
    .Y(_03540_),
    .B1(_03402_));
 sg13g2_or2_1 _09491_ (.X(_03541_),
    .B(_03540_),
    .A(_03538_));
 sg13g2_o21ai_1 _09492_ (.B1(_03405_),
    .Y(_03542_),
    .A1(_03273_),
    .A2(_03404_));
 sg13g2_a21oi_1 _09493_ (.A1(_03281_),
    .A2(_03407_),
    .Y(_03543_),
    .B1(_03542_));
 sg13g2_xor2_1 _09494_ (.B(_03543_),
    .A(_03541_),
    .X(_03544_));
 sg13g2_o21ai_1 _09495_ (.B1(net1751),
    .Y(_03545_),
    .A1(net1398),
    .A2(_03544_));
 sg13g2_a21oi_1 _09496_ (.A1(net1398),
    .A2(_05548_),
    .Y(_00322_),
    .B1(_03545_));
 sg13g2_a21o_1 _09497_ (.A2(_03527_),
    .A1(_03414_),
    .B1(_03525_),
    .X(_03546_));
 sg13g2_nand2_1 _09498_ (.Y(_03547_),
    .A(_03447_),
    .B(_03449_));
 sg13g2_or2_1 _09499_ (.X(_03548_),
    .B(_03428_),
    .A(_03419_));
 sg13g2_nand2_1 _09500_ (.Y(_03549_),
    .A(_03419_),
    .B(_03428_));
 sg13g2_a22oi_1 _09501_ (.Y(_03550_),
    .B1(_03548_),
    .B2(_03549_),
    .A2(_03429_),
    .A1(_03420_));
 sg13g2_a21oi_2 _09502_ (.B1(_03550_),
    .Y(_03551_),
    .A2(_03449_),
    .A1(_03447_));
 sg13g2_inv_1 _09503_ (.Y(_03552_),
    .A(_03551_));
 sg13g2_xnor2_1 _09504_ (.Y(_03553_),
    .A(_03547_),
    .B(_03550_));
 sg13g2_o21ai_1 _09505_ (.B1(_03521_),
    .Y(_03554_),
    .A1(_03450_),
    .A2(_03522_));
 sg13g2_o21ai_1 _09506_ (.B1(_03444_),
    .Y(_03555_),
    .A1(_03430_),
    .A2(_03445_));
 sg13g2_o21ai_1 _09507_ (.B1(_03474_),
    .Y(_03556_),
    .A1(_03453_),
    .A2(_03475_));
 sg13g2_a21oi_2 _09508_ (.B1(_03423_),
    .Y(_03557_),
    .A2(_03425_),
    .A1(_03421_));
 sg13g2_nand2_1 _09509_ (.Y(_03558_),
    .A(net1498),
    .B(net1537));
 sg13g2_nand2_1 _09510_ (.Y(_03559_),
    .A(net1500),
    .B(net1527));
 sg13g2_nand2_1 _09511_ (.Y(_03560_),
    .A(net1503),
    .B(net1527));
 sg13g2_or2_1 _09512_ (.X(_03561_),
    .B(_03560_),
    .A(_03422_));
 sg13g2_xnor2_1 _09513_ (.Y(_03562_),
    .A(_03422_),
    .B(_03560_));
 sg13g2_xor2_1 _09514_ (.B(_03562_),
    .A(_03558_),
    .X(_03563_));
 sg13g2_nand2b_1 _09515_ (.Y(_03564_),
    .B(_03563_),
    .A_N(_03557_));
 sg13g2_xnor2_1 _09516_ (.Y(_03565_),
    .A(_03557_),
    .B(_03563_));
 sg13g2_and2_1 _09517_ (.A(net1487),
    .B(net1558),
    .X(_03566_));
 sg13g2_nand2_2 _09518_ (.Y(_03567_),
    .A(net1487),
    .B(net1558));
 sg13g2_a22oi_1 _09519_ (.Y(_03568_),
    .B1(net1549),
    .B2(net1490),
    .A2(net1543),
    .A1(net1493));
 sg13g2_nand4_1 _09520_ (.B(net1493),
    .C(net1543),
    .A(net1491),
    .Y(_03569_),
    .D(net1549));
 sg13g2_nor2b_1 _09521_ (.A(_03568_),
    .B_N(_03569_),
    .Y(_03570_));
 sg13g2_xnor2_1 _09522_ (.Y(_03571_),
    .A(_03567_),
    .B(_03570_));
 sg13g2_nand2_1 _09523_ (.Y(_03572_),
    .A(_03565_),
    .B(_03571_));
 sg13g2_xnor2_1 _09524_ (.Y(_03573_),
    .A(_03565_),
    .B(_03571_));
 sg13g2_o21ai_1 _09525_ (.B1(_03441_),
    .Y(_03574_),
    .A1(_03433_),
    .A2(_03442_));
 sg13g2_o21ai_1 _09526_ (.B1(_03438_),
    .Y(_03575_),
    .A1(_03435_),
    .A2(_03439_));
 sg13g2_or2_1 _09527_ (.X(_03576_),
    .B(_03459_),
    .A(_03457_));
 sg13g2_nand2_1 _09528_ (.Y(_03577_),
    .A(net1508),
    .B(net1520));
 sg13g2_nand2_1 _09529_ (.Y(_03578_),
    .A(net1510),
    .B(net1728));
 sg13g2_nand2_1 _09530_ (.Y(_03579_),
    .A(net1562),
    .B(net1728));
 sg13g2_or2_1 _09531_ (.X(_03580_),
    .B(_03578_),
    .A(_03437_));
 sg13g2_xnor2_1 _09532_ (.Y(_03581_),
    .A(_03436_),
    .B(_03579_));
 sg13g2_xor2_1 _09533_ (.B(_03581_),
    .A(_03577_),
    .X(_03582_));
 sg13g2_xnor2_1 _09534_ (.Y(_03583_),
    .A(_03576_),
    .B(_03582_));
 sg13g2_nor2b_1 _09535_ (.A(_03583_),
    .B_N(_03575_),
    .Y(_03584_));
 sg13g2_xor2_1 _09536_ (.B(_03583_),
    .A(_03575_),
    .X(_03585_));
 sg13g2_nand2b_1 _09537_ (.Y(_03586_),
    .B(_03574_),
    .A_N(_03585_));
 sg13g2_xor2_1 _09538_ (.B(_03585_),
    .A(_03574_),
    .X(_03587_));
 sg13g2_xor2_1 _09539_ (.B(_03587_),
    .A(_03573_),
    .X(_03588_));
 sg13g2_xnor2_1 _09540_ (.Y(_03589_),
    .A(_03556_),
    .B(_03588_));
 sg13g2_nor2b_1 _09541_ (.A(_03589_),
    .B_N(_03555_),
    .Y(_03590_));
 sg13g2_xnor2_1 _09542_ (.Y(_03591_),
    .A(_03555_),
    .B(_03589_));
 sg13g2_o21ai_1 _09543_ (.B1(_03516_),
    .Y(_03592_),
    .A1(_03476_),
    .A2(_03517_));
 sg13g2_o21ai_1 _09544_ (.B1(_03471_),
    .Y(_03593_),
    .A1(_03462_),
    .A2(_03472_));
 sg13g2_o21ai_1 _09545_ (.B1(_03487_),
    .Y(_03594_),
    .A1(_03479_),
    .A2(_03488_));
 sg13g2_inv_1 _09546_ (.Y(_03595_),
    .A(_03594_));
 sg13g2_nand2_1 _09547_ (.Y(_03596_),
    .A(net1566),
    .B(net1721));
 sg13g2_nand2_1 _09548_ (.Y(_03597_),
    .A(net1570),
    .B(net1710));
 sg13g2_nand2_1 _09549_ (.Y(_03598_),
    .A(net1575),
    .B(net1710));
 sg13g2_xor2_1 _09550_ (.B(_03598_),
    .A(_03456_),
    .X(_03599_));
 sg13g2_nand2b_1 _09551_ (.Y(_03600_),
    .B(_03599_),
    .A_N(_03596_));
 sg13g2_xnor2_1 _09552_ (.Y(_03601_),
    .A(_03596_),
    .B(_03599_));
 sg13g2_or2_1 _09553_ (.X(_03602_),
    .B(_03468_),
    .A(_03466_));
 sg13g2_nand2_1 _09554_ (.Y(_03603_),
    .A(net1580),
    .B(net1704));
 sg13g2_nand2_1 _09555_ (.Y(_03604_),
    .A(net1585),
    .B(net1696));
 sg13g2_nand2_1 _09556_ (.Y(_03605_),
    .A(net1592),
    .B(net1696));
 sg13g2_xor2_1 _09557_ (.B(_03605_),
    .A(_03465_),
    .X(_03606_));
 sg13g2_nand2b_1 _09558_ (.Y(_03607_),
    .B(_03606_),
    .A_N(_03603_));
 sg13g2_xnor2_1 _09559_ (.Y(_03608_),
    .A(_03603_),
    .B(_03606_));
 sg13g2_and2_1 _09560_ (.A(_03602_),
    .B(_03608_),
    .X(_03609_));
 sg13g2_xnor2_1 _09561_ (.Y(_03610_),
    .A(_03602_),
    .B(_03608_));
 sg13g2_inv_1 _09562_ (.Y(_03611_),
    .A(_03610_));
 sg13g2_xor2_1 _09563_ (.B(_03610_),
    .A(_03601_),
    .X(_03612_));
 sg13g2_xor2_1 _09564_ (.B(_03612_),
    .A(_03594_),
    .X(_03613_));
 sg13g2_nand2b_1 _09565_ (.Y(_03614_),
    .B(_03593_),
    .A_N(_03613_));
 sg13g2_xnor2_1 _09566_ (.Y(_03615_),
    .A(_03593_),
    .B(_03613_));
 sg13g2_o21ai_1 _09567_ (.B1(_03511_),
    .Y(_03616_),
    .A1(_03489_),
    .A2(_03512_));
 sg13g2_o21ai_1 _09568_ (.B1(_03499_),
    .Y(_03617_),
    .A1(_03500_),
    .A2(_03507_));
 sg13g2_o21ai_1 _09569_ (.B1(_03494_),
    .Y(_03618_),
    .A1(_03492_),
    .A2(_03495_));
 sg13g2_nand2_1 _09570_ (.Y(_03619_),
    .A(net1631),
    .B(net1663));
 sg13g2_and4_1 _09571_ (.A(net1636),
    .B(net1646),
    .C(net1657),
    .D(net1661),
    .X(_03620_));
 sg13g2_a22oi_1 _09572_ (.Y(_03621_),
    .B1(net1661),
    .B2(net1636),
    .A2(net1657),
    .A1(net1646));
 sg13g2_or3_1 _09573_ (.A(_03619_),
    .B(_03620_),
    .C(_03621_),
    .X(_03622_));
 sg13g2_o21ai_1 _09574_ (.B1(_03619_),
    .Y(_03623_),
    .A1(_03620_),
    .A2(_03621_));
 sg13g2_nand3_1 _09575_ (.B(_03622_),
    .C(_03623_),
    .A(_03618_),
    .Y(_03624_));
 sg13g2_a21o_1 _09576_ (.A2(_03623_),
    .A1(_03622_),
    .B1(_03618_),
    .X(_03625_));
 sg13g2_nand2_1 _09577_ (.Y(_03626_),
    .A(net1614),
    .B(net1675));
 sg13g2_nand2_1 _09578_ (.Y(_03627_),
    .A(net1618),
    .B(net1668));
 sg13g2_nand2_1 _09579_ (.Y(_03628_),
    .A(net1623),
    .B(net1668));
 sg13g2_xor2_1 _09580_ (.B(_03628_),
    .A(_03502_),
    .X(_03629_));
 sg13g2_nand2b_1 _09581_ (.Y(_03630_),
    .B(_03629_),
    .A_N(_03626_));
 sg13g2_xnor2_1 _09582_ (.Y(_03631_),
    .A(_03626_),
    .B(_03629_));
 sg13g2_nand3_1 _09583_ (.B(_03625_),
    .C(_03631_),
    .A(_03624_),
    .Y(_03632_));
 sg13g2_a21o_1 _09584_ (.A2(_03625_),
    .A1(_03624_),
    .B1(_03631_),
    .X(_03633_));
 sg13g2_nand3_1 _09585_ (.B(_03632_),
    .C(_03633_),
    .A(_03617_),
    .Y(_03634_));
 sg13g2_a21o_1 _09586_ (.A2(_03633_),
    .A1(_03632_),
    .B1(_03617_),
    .X(_03635_));
 sg13g2_o21ai_1 _09587_ (.B1(_03484_),
    .Y(_03636_),
    .A1(_03481_),
    .A2(_03485_));
 sg13g2_or2_1 _09588_ (.X(_03637_),
    .B(_03505_),
    .A(_03503_));
 sg13g2_nand2_1 _09589_ (.Y(_03638_),
    .A(net1600),
    .B(net1691));
 sg13g2_nand2_2 _09590_ (.Y(_03639_),
    .A(net1605),
    .B(net1681));
 sg13g2_nand2_1 _09591_ (.Y(_03640_),
    .A(net1607),
    .B(net1681));
 sg13g2_or2_1 _09592_ (.X(_03641_),
    .B(_03639_),
    .A(_03483_));
 sg13g2_xnor2_1 _09593_ (.Y(_03642_),
    .A(_03482_),
    .B(_03640_));
 sg13g2_xor2_1 _09594_ (.B(_03642_),
    .A(_03638_),
    .X(_03643_));
 sg13g2_xnor2_1 _09595_ (.Y(_03644_),
    .A(_03637_),
    .B(_03643_));
 sg13g2_nor2b_1 _09596_ (.A(_03644_),
    .B_N(_03636_),
    .Y(_03645_));
 sg13g2_xnor2_1 _09597_ (.Y(_03646_),
    .A(_03636_),
    .B(_03644_));
 sg13g2_nand3_1 _09598_ (.B(_03635_),
    .C(_03646_),
    .A(_03634_),
    .Y(_03647_));
 sg13g2_a21o_1 _09599_ (.A2(_03635_),
    .A1(_03634_),
    .B1(_03646_),
    .X(_03648_));
 sg13g2_nand3_1 _09600_ (.B(_03647_),
    .C(_03648_),
    .A(_03616_),
    .Y(_03649_));
 sg13g2_a21o_1 _09601_ (.A2(_03648_),
    .A1(_03647_),
    .B1(_03616_),
    .X(_03650_));
 sg13g2_nand3_1 _09602_ (.B(_03649_),
    .C(_03650_),
    .A(_03615_),
    .Y(_03651_));
 sg13g2_a21o_1 _09603_ (.A2(_03650_),
    .A1(_03649_),
    .B1(_03615_),
    .X(_03652_));
 sg13g2_nand3_1 _09604_ (.B(_03651_),
    .C(_03652_),
    .A(_03592_),
    .Y(_03653_));
 sg13g2_a21o_1 _09605_ (.A2(_03652_),
    .A1(_03651_),
    .B1(_03592_),
    .X(_03654_));
 sg13g2_nand3_1 _09606_ (.B(_03653_),
    .C(_03654_),
    .A(_03591_),
    .Y(_03655_));
 sg13g2_a21o_1 _09607_ (.A2(_03654_),
    .A1(_03653_),
    .B1(_03591_),
    .X(_03656_));
 sg13g2_nand3_1 _09608_ (.B(_03655_),
    .C(_03656_),
    .A(_03554_),
    .Y(_03657_));
 sg13g2_a21o_1 _09609_ (.A2(_03656_),
    .A1(_03655_),
    .B1(_03554_),
    .X(_03658_));
 sg13g2_nand3_1 _09610_ (.B(_03657_),
    .C(_03658_),
    .A(_03553_),
    .Y(_03659_));
 sg13g2_a21o_1 _09611_ (.A2(_03658_),
    .A1(_03657_),
    .B1(_03553_),
    .X(_03660_));
 sg13g2_and3_1 _09612_ (.X(_03661_),
    .A(_03546_),
    .B(_03659_),
    .C(_03660_));
 sg13g2_a21oi_1 _09613_ (.A1(_03659_),
    .A2(_03660_),
    .Y(_03662_),
    .B1(_03546_));
 sg13g2_o21ai_1 _09614_ (.B1(_03413_),
    .Y(_03663_),
    .A1(_03661_),
    .A2(_03662_));
 sg13g2_or3_1 _09615_ (.A(_03413_),
    .B(_03661_),
    .C(_03662_),
    .X(_03664_));
 sg13g2_o21ai_1 _09616_ (.B1(_03530_),
    .Y(_03665_),
    .A1(_03288_),
    .A2(_03531_));
 sg13g2_nand3_1 _09617_ (.B(_03664_),
    .C(_03665_),
    .A(_03663_),
    .Y(_03666_));
 sg13g2_a21o_1 _09618_ (.A2(_03664_),
    .A1(_03663_),
    .B1(_03665_),
    .X(_03667_));
 sg13g2_and2_1 _09619_ (.A(_03666_),
    .B(_03667_),
    .X(_03668_));
 sg13g2_a21oi_1 _09620_ (.A1(_03666_),
    .A2(_03667_),
    .Y(_03669_),
    .B1(_03535_));
 sg13g2_and3_1 _09621_ (.X(_03670_),
    .A(_03535_),
    .B(_03666_),
    .C(_03667_));
 sg13g2_or2_1 _09622_ (.X(_03671_),
    .B(_03670_),
    .A(_03669_));
 sg13g2_o21ai_1 _09623_ (.B1(_03539_),
    .Y(_03672_),
    .A1(_03541_),
    .A2(_03543_));
 sg13g2_xor2_1 _09624_ (.B(_03672_),
    .A(_03671_),
    .X(_03673_));
 sg13g2_o21ai_1 _09625_ (.B1(net1751),
    .Y(_03674_),
    .A1(net1470),
    .A2(net618));
 sg13g2_a21oi_1 _09626_ (.A1(net1470),
    .A2(_03673_),
    .Y(_00323_),
    .B1(_03674_));
 sg13g2_nor4_1 _09627_ (.A(_03538_),
    .B(_03540_),
    .C(_03669_),
    .D(_03670_),
    .Y(_03675_));
 sg13g2_a221oi_1 _09628_ (.B2(_03542_),
    .C1(_03670_),
    .B1(_03675_),
    .A1(_03538_),
    .Y(_03676_),
    .A2(_03668_));
 sg13g2_nand3b_1 _09629_ (.B(_03407_),
    .C(_03675_),
    .Y(_03677_),
    .A_N(_03274_));
 sg13g2_o21ai_1 _09630_ (.B1(_03676_),
    .Y(_03678_),
    .A1(_03280_),
    .A2(_03677_));
 sg13g2_nand2b_2 _09631_ (.Y(_03679_),
    .B(_03664_),
    .A_N(_03661_));
 sg13g2_nand2_2 _09632_ (.Y(_03680_),
    .A(_03657_),
    .B(_03659_));
 sg13g2_a21oi_2 _09633_ (.B1(_03590_),
    .Y(_03681_),
    .A2(_03588_),
    .A1(_03556_));
 sg13g2_nor2_1 _09634_ (.A(_03567_),
    .B(_03568_),
    .Y(_03682_));
 sg13g2_a21o_1 _09635_ (.A2(_03569_),
    .A1(_03567_),
    .B1(_03682_),
    .X(_03683_));
 sg13g2_a21oi_1 _09636_ (.A1(_03564_),
    .A2(_03572_),
    .Y(_03684_),
    .B1(_03683_));
 sg13g2_nand3_1 _09637_ (.B(_03572_),
    .C(_03683_),
    .A(_03564_),
    .Y(_03685_));
 sg13g2_nand2b_1 _09638_ (.Y(_03686_),
    .B(_03685_),
    .A_N(_03684_));
 sg13g2_nor2_1 _09639_ (.A(_03548_),
    .B(_03686_),
    .Y(_03687_));
 sg13g2_xor2_1 _09640_ (.B(_03686_),
    .A(_03548_),
    .X(_03688_));
 sg13g2_nand2b_1 _09641_ (.Y(_03689_),
    .B(_03688_),
    .A_N(_03681_));
 sg13g2_xor2_1 _09642_ (.B(_03688_),
    .A(_03681_),
    .X(_03690_));
 sg13g2_nand2_2 _09643_ (.Y(_03691_),
    .A(_03653_),
    .B(_03655_));
 sg13g2_o21ai_1 _09644_ (.B1(_03586_),
    .Y(_03692_),
    .A1(_03573_),
    .A2(_03587_));
 sg13g2_o21ai_1 _09645_ (.B1(_03614_),
    .Y(_03693_),
    .A1(_03595_),
    .A2(_03612_));
 sg13g2_a21o_2 _09646_ (.A2(_03582_),
    .A1(_03576_),
    .B1(_03584_),
    .X(_03694_));
 sg13g2_o21ai_1 _09647_ (.B1(_03580_),
    .Y(_03695_),
    .A1(_03577_),
    .A2(_03581_));
 sg13g2_o21ai_1 _09648_ (.B1(_03600_),
    .Y(_03696_),
    .A1(_03456_),
    .A2(_03598_));
 sg13g2_nand2_1 _09649_ (.Y(_03697_),
    .A(net1508),
    .B(net1514));
 sg13g2_nand2_1 _09650_ (.Y(_03698_),
    .A(net1510),
    .B(net1721));
 sg13g2_nand2_1 _09651_ (.Y(_03699_),
    .A(net1562),
    .B(net1721));
 sg13g2_or2_1 _09652_ (.X(_03700_),
    .B(_03698_),
    .A(_03579_));
 sg13g2_xnor2_1 _09653_ (.Y(_03701_),
    .A(_03578_),
    .B(_03699_));
 sg13g2_xor2_1 _09654_ (.B(_03701_),
    .A(_03697_),
    .X(_03702_));
 sg13g2_xnor2_1 _09655_ (.Y(_03703_),
    .A(_03696_),
    .B(_03702_));
 sg13g2_nor2b_1 _09656_ (.A(_03703_),
    .B_N(_03695_),
    .Y(_03704_));
 sg13g2_xor2_1 _09657_ (.B(_03703_),
    .A(_03695_),
    .X(_03705_));
 sg13g2_nand2b_1 _09658_ (.Y(_03706_),
    .B(_03694_),
    .A_N(_03705_));
 sg13g2_xor2_1 _09659_ (.B(_03705_),
    .A(_03694_),
    .X(_03707_));
 sg13g2_and2_1 _09660_ (.A(net1487),
    .B(net1549),
    .X(_03708_));
 sg13g2_nand2_2 _09661_ (.Y(_03709_),
    .A(net1488),
    .B(net1549));
 sg13g2_nand2_1 _09662_ (.Y(_03710_),
    .A(net1494),
    .B(net1537));
 sg13g2_nor3_1 _09663_ (.A(_05552_),
    .B(_05573_),
    .C(_03710_),
    .Y(_03711_));
 sg13g2_a22oi_1 _09664_ (.Y(_03712_),
    .B1(net1543),
    .B2(net1490),
    .A2(net1537),
    .A1(net1494));
 sg13g2_nor2_1 _09665_ (.A(_03711_),
    .B(_03712_),
    .Y(_03713_));
 sg13g2_xnor2_1 _09666_ (.Y(_03714_),
    .A(_03709_),
    .B(_03713_));
 sg13g2_o21ai_1 _09667_ (.B1(_03561_),
    .Y(_03715_),
    .A1(_03558_),
    .A2(_03562_));
 sg13g2_nand2_1 _09668_ (.Y(_03716_),
    .A(net1498),
    .B(net1532));
 sg13g2_nand2_1 _09669_ (.Y(_03717_),
    .A(net1500),
    .B(net1519));
 sg13g2_nand2_1 _09670_ (.Y(_03718_),
    .A(net1503),
    .B(net1520));
 sg13g2_xor2_1 _09671_ (.B(_03718_),
    .A(_03559_),
    .X(_03719_));
 sg13g2_nand2b_1 _09672_ (.Y(_03720_),
    .B(_03719_),
    .A_N(_03716_));
 sg13g2_xnor2_1 _09673_ (.Y(_03721_),
    .A(_03716_),
    .B(_03719_));
 sg13g2_nand2_1 _09674_ (.Y(_03722_),
    .A(_03715_),
    .B(_03721_));
 sg13g2_xor2_1 _09675_ (.B(_03721_),
    .A(_03715_),
    .X(_03723_));
 sg13g2_nand2_1 _09676_ (.Y(_03724_),
    .A(_03714_),
    .B(_03723_));
 sg13g2_xnor2_1 _09677_ (.Y(_03725_),
    .A(_03714_),
    .B(_03723_));
 sg13g2_xor2_1 _09678_ (.B(_03725_),
    .A(_03707_),
    .X(_03726_));
 sg13g2_nand2_1 _09679_ (.Y(_03727_),
    .A(_03693_),
    .B(_03726_));
 sg13g2_xnor2_1 _09680_ (.Y(_03728_),
    .A(_03693_),
    .B(_03726_));
 sg13g2_nand2b_1 _09681_ (.Y(_03729_),
    .B(_03692_),
    .A_N(_03728_));
 sg13g2_xor2_1 _09682_ (.B(_03728_),
    .A(_03692_),
    .X(_03730_));
 sg13g2_nand2_1 _09683_ (.Y(_03731_),
    .A(_03649_),
    .B(_03651_));
 sg13g2_nand2_1 _09684_ (.Y(_03732_),
    .A(_03634_),
    .B(_03647_));
 sg13g2_nand2_1 _09685_ (.Y(_03733_),
    .A(_03624_),
    .B(_03632_));
 sg13g2_nand2b_1 _09686_ (.Y(_03734_),
    .B(_03622_),
    .A_N(_03620_));
 sg13g2_o21ai_1 _09687_ (.B1(net1657),
    .Y(_03735_),
    .A1(net1639),
    .A2(net1649));
 sg13g2_nand3_1 _09688_ (.B(net1649),
    .C(net1657),
    .A(net1639),
    .Y(_03736_));
 sg13g2_nor2b_1 _09689_ (.A(_03735_),
    .B_N(_03736_),
    .Y(_03737_));
 sg13g2_nand2_1 _09690_ (.Y(_03738_),
    .A(net1631),
    .B(net1660));
 sg13g2_xnor2_1 _09691_ (.Y(_03739_),
    .A(_03737_),
    .B(_03738_));
 sg13g2_nand2_1 _09692_ (.Y(_03740_),
    .A(_03734_),
    .B(_03739_));
 sg13g2_xnor2_1 _09693_ (.Y(_03741_),
    .A(_03734_),
    .B(_03739_));
 sg13g2_nand2_1 _09694_ (.Y(_03742_),
    .A(net1614),
    .B(net1671));
 sg13g2_nand2_1 _09695_ (.Y(_03743_),
    .A(net1619),
    .B(net1663));
 sg13g2_nand2_2 _09696_ (.Y(_03744_),
    .A(net1623),
    .B(net1664));
 sg13g2_xor2_1 _09697_ (.B(_03744_),
    .A(_03627_),
    .X(_03745_));
 sg13g2_nand2b_1 _09698_ (.Y(_03746_),
    .B(_03745_),
    .A_N(_03742_));
 sg13g2_xor2_1 _09699_ (.B(_03745_),
    .A(_03742_),
    .X(_03747_));
 sg13g2_xor2_1 _09700_ (.B(_03747_),
    .A(_03741_),
    .X(_03748_));
 sg13g2_nand2_1 _09701_ (.Y(_03749_),
    .A(_03733_),
    .B(_03748_));
 sg13g2_xnor2_1 _09702_ (.Y(_03750_),
    .A(_03733_),
    .B(_03748_));
 sg13g2_o21ai_1 _09703_ (.B1(_03641_),
    .Y(_03751_),
    .A1(_03638_),
    .A2(_03642_));
 sg13g2_inv_1 _09704_ (.Y(_03752_),
    .A(_03751_));
 sg13g2_o21ai_1 _09705_ (.B1(_03630_),
    .Y(_03753_),
    .A1(_03502_),
    .A2(_03628_));
 sg13g2_nand2_1 _09706_ (.Y(_03754_),
    .A(net1598),
    .B(net1687));
 sg13g2_nand2_1 _09707_ (.Y(_03755_),
    .A(net1603),
    .B(net1675));
 sg13g2_nand2_2 _09708_ (.Y(_03756_),
    .A(net1607),
    .B(net1675));
 sg13g2_xnor2_1 _09709_ (.Y(_03757_),
    .A(_03639_),
    .B(_03756_));
 sg13g2_or2_1 _09710_ (.X(_03758_),
    .B(_03757_),
    .A(_03754_));
 sg13g2_xor2_1 _09711_ (.B(_03757_),
    .A(_03754_),
    .X(_03759_));
 sg13g2_nand2_1 _09712_ (.Y(_03760_),
    .A(_03753_),
    .B(_03759_));
 sg13g2_xnor2_1 _09713_ (.Y(_03761_),
    .A(_03753_),
    .B(_03759_));
 sg13g2_xnor2_1 _09714_ (.Y(_03762_),
    .A(_03752_),
    .B(_03761_));
 sg13g2_xor2_1 _09715_ (.B(_03762_),
    .A(_03750_),
    .X(_03763_));
 sg13g2_nand2_1 _09716_ (.Y(_03764_),
    .A(_03732_),
    .B(_03763_));
 sg13g2_xnor2_1 _09717_ (.Y(_03765_),
    .A(_03732_),
    .B(_03763_));
 sg13g2_a21o_1 _09718_ (.A2(_03611_),
    .A1(_03601_),
    .B1(_03609_),
    .X(_03766_));
 sg13g2_a21o_2 _09719_ (.A2(_03643_),
    .A1(_03637_),
    .B1(_03645_),
    .X(_03767_));
 sg13g2_nand2_1 _09720_ (.Y(_03768_),
    .A(net1566),
    .B(net1715));
 sg13g2_nand2_1 _09721_ (.Y(_03769_),
    .A(net1570),
    .B(net1704));
 sg13g2_nand2_1 _09722_ (.Y(_03770_),
    .A(net1575),
    .B(net1704));
 sg13g2_xor2_1 _09723_ (.B(_03770_),
    .A(_03597_),
    .X(_03771_));
 sg13g2_nand2b_1 _09724_ (.Y(_03772_),
    .B(_03771_),
    .A_N(_03768_));
 sg13g2_xor2_1 _09725_ (.B(_03771_),
    .A(_03768_),
    .X(_03773_));
 sg13g2_o21ai_1 _09726_ (.B1(_03607_),
    .Y(_03774_),
    .A1(_03465_),
    .A2(_03605_));
 sg13g2_nand2_1 _09727_ (.Y(_03775_),
    .A(net1581),
    .B(net1701));
 sg13g2_nand2_1 _09728_ (.Y(_03776_),
    .A(net1585),
    .B(net1691));
 sg13g2_nand2_1 _09729_ (.Y(_03777_),
    .A(net1592),
    .B(net1691));
 sg13g2_xor2_1 _09730_ (.B(_03777_),
    .A(_03604_),
    .X(_03778_));
 sg13g2_nand2b_1 _09731_ (.Y(_03779_),
    .B(_03778_),
    .A_N(_03775_));
 sg13g2_xnor2_1 _09732_ (.Y(_03780_),
    .A(_03775_),
    .B(_03778_));
 sg13g2_xnor2_1 _09733_ (.Y(_03781_),
    .A(_03774_),
    .B(_03780_));
 sg13g2_nor2_1 _09734_ (.A(_03773_),
    .B(_03781_),
    .Y(_03782_));
 sg13g2_xnor2_1 _09735_ (.Y(_03783_),
    .A(_03773_),
    .B(_03781_));
 sg13g2_nand2b_1 _09736_ (.Y(_03784_),
    .B(_03767_),
    .A_N(_03783_));
 sg13g2_xor2_1 _09737_ (.B(_03783_),
    .A(_03767_),
    .X(_03785_));
 sg13g2_nand2b_1 _09738_ (.Y(_03786_),
    .B(_03766_),
    .A_N(_03785_));
 sg13g2_xor2_1 _09739_ (.B(_03785_),
    .A(_03766_),
    .X(_03787_));
 sg13g2_xor2_1 _09740_ (.B(_03787_),
    .A(_03765_),
    .X(_03788_));
 sg13g2_nand2_1 _09741_ (.Y(_03789_),
    .A(_03731_),
    .B(_03788_));
 sg13g2_xnor2_1 _09742_ (.Y(_03790_),
    .A(_03731_),
    .B(_03788_));
 sg13g2_xor2_1 _09743_ (.B(_03790_),
    .A(_03730_),
    .X(_03791_));
 sg13g2_nand2_1 _09744_ (.Y(_03792_),
    .A(_03691_),
    .B(_03791_));
 sg13g2_xnor2_1 _09745_ (.Y(_03793_),
    .A(_03691_),
    .B(_03791_));
 sg13g2_xor2_1 _09746_ (.B(_03793_),
    .A(_03690_),
    .X(_03794_));
 sg13g2_nand2_1 _09747_ (.Y(_03795_),
    .A(_03680_),
    .B(_03794_));
 sg13g2_xnor2_1 _09748_ (.Y(_03796_),
    .A(_03680_),
    .B(_03794_));
 sg13g2_xnor2_1 _09749_ (.Y(_03797_),
    .A(_03551_),
    .B(_03796_));
 sg13g2_nand2_1 _09750_ (.Y(_03798_),
    .A(_03679_),
    .B(_03797_));
 sg13g2_xor2_1 _09751_ (.B(_03797_),
    .A(_03679_),
    .X(_03799_));
 sg13g2_nor2b_1 _09752_ (.A(_03666_),
    .B_N(_03799_),
    .Y(_03800_));
 sg13g2_xor2_1 _09753_ (.B(_03799_),
    .A(_03666_),
    .X(_03801_));
 sg13g2_inv_1 _09754_ (.Y(_03802_),
    .A(_03801_));
 sg13g2_xnor2_1 _09755_ (.Y(_03803_),
    .A(_03678_),
    .B(_03802_));
 sg13g2_o21ai_1 _09756_ (.B1(net1751),
    .Y(_03804_),
    .A1(net1470),
    .A2(net624));
 sg13g2_a21oi_1 _09757_ (.A1(net1470),
    .A2(_03803_),
    .Y(_00324_),
    .B1(_03804_));
 sg13g2_a21oi_1 _09758_ (.A1(_03678_),
    .A2(_03802_),
    .Y(_03805_),
    .B1(_03800_));
 sg13g2_o21ai_1 _09759_ (.B1(_03792_),
    .Y(_03806_),
    .A1(_03690_),
    .A2(_03793_));
 sg13g2_nor2_2 _09760_ (.A(_05574_),
    .B(_03567_),
    .Y(_03807_));
 sg13g2_nand2_2 _09761_ (.Y(_03808_),
    .A(net1549),
    .B(_03566_));
 sg13g2_o21ai_1 _09762_ (.B1(_03808_),
    .Y(_03809_),
    .A1(_03566_),
    .A2(_03708_));
 sg13g2_a21o_1 _09763_ (.A2(_03713_),
    .A1(_03708_),
    .B1(_03711_),
    .X(_03810_));
 sg13g2_nand2b_1 _09764_ (.Y(_03811_),
    .B(_03810_),
    .A_N(_03809_));
 sg13g2_xor2_1 _09765_ (.B(_03810_),
    .A(_03809_),
    .X(_03812_));
 sg13g2_a21o_1 _09766_ (.A2(_03724_),
    .A1(_03722_),
    .B1(_03812_),
    .X(_03813_));
 sg13g2_nand3_1 _09767_ (.B(_03724_),
    .C(_03812_),
    .A(_03722_),
    .Y(_03814_));
 sg13g2_nand2_1 _09768_ (.Y(_03815_),
    .A(_03813_),
    .B(_03814_));
 sg13g2_nor2_1 _09769_ (.A(_03682_),
    .B(_03684_),
    .Y(_03816_));
 sg13g2_xnor2_1 _09770_ (.Y(_03817_),
    .A(_03815_),
    .B(_03816_));
 sg13g2_a21oi_1 _09771_ (.A1(_03727_),
    .A2(_03729_),
    .Y(_03818_),
    .B1(_03817_));
 sg13g2_nand3_1 _09772_ (.B(_03729_),
    .C(_03817_),
    .A(_03727_),
    .Y(_03819_));
 sg13g2_nor2b_1 _09773_ (.A(_03818_),
    .B_N(_03819_),
    .Y(_03820_));
 sg13g2_xnor2_1 _09774_ (.Y(_03821_),
    .A(_03687_),
    .B(_03820_));
 sg13g2_o21ai_1 _09775_ (.B1(_03789_),
    .Y(_03822_),
    .A1(_03730_),
    .A2(_03790_));
 sg13g2_o21ai_1 _09776_ (.B1(_03764_),
    .Y(_03823_),
    .A1(_03765_),
    .A2(_03787_));
 sg13g2_o21ai_1 _09777_ (.B1(_03749_),
    .Y(_03824_),
    .A1(_03750_),
    .A2(_03762_));
 sg13g2_o21ai_1 _09778_ (.B1(_03740_),
    .Y(_03825_),
    .A1(_03741_),
    .A2(_03747_));
 sg13g2_nand2_1 _09779_ (.Y(_03826_),
    .A(net1614),
    .B(net1669));
 sg13g2_nand2_1 _09780_ (.Y(_03827_),
    .A(net1619),
    .B(net1660));
 sg13g2_nand2_1 _09781_ (.Y(_03828_),
    .A(net1623),
    .B(net1660));
 sg13g2_or2_1 _09782_ (.X(_03829_),
    .B(_03827_),
    .A(_03744_));
 sg13g2_xor2_1 _09783_ (.B(_03828_),
    .A(_03743_),
    .X(_03830_));
 sg13g2_nand2b_1 _09784_ (.Y(_03831_),
    .B(_03830_),
    .A_N(_03826_));
 sg13g2_xor2_1 _09785_ (.B(_03830_),
    .A(_03826_),
    .X(_03832_));
 sg13g2_o21ai_1 _09786_ (.B1(_03736_),
    .Y(_03833_),
    .A1(_03735_),
    .A2(_03738_));
 sg13g2_nand2_1 _09787_ (.Y(_03834_),
    .A(net1631),
    .B(net1657));
 sg13g2_xnor2_1 _09788_ (.Y(_03835_),
    .A(_03737_),
    .B(_03834_));
 sg13g2_or2_1 _09789_ (.X(_03836_),
    .B(_03736_),
    .A(_05558_));
 sg13g2_inv_4 _09790_ (.A(_03836_),
    .Y(_03837_));
 sg13g2_xnor2_1 _09791_ (.Y(_03838_),
    .A(_03833_),
    .B(_03835_));
 sg13g2_xor2_1 _09792_ (.B(_03838_),
    .A(_03832_),
    .X(_03839_));
 sg13g2_nand2_1 _09793_ (.Y(_03840_),
    .A(_03825_),
    .B(_03839_));
 sg13g2_xnor2_1 _09794_ (.Y(_03841_),
    .A(_03825_),
    .B(_03839_));
 sg13g2_o21ai_1 _09795_ (.B1(_03758_),
    .Y(_03842_),
    .A1(_03639_),
    .A2(_03756_));
 sg13g2_inv_1 _09796_ (.Y(_03843_),
    .A(_03842_));
 sg13g2_o21ai_1 _09797_ (.B1(_03746_),
    .Y(_03844_),
    .A1(_03627_),
    .A2(_03744_));
 sg13g2_nand2_1 _09798_ (.Y(_03845_),
    .A(net1598),
    .B(net1681));
 sg13g2_nand2_1 _09799_ (.Y(_03846_),
    .A(net1603),
    .B(net1671));
 sg13g2_nand2_1 _09800_ (.Y(_03847_),
    .A(net1607),
    .B(net1671));
 sg13g2_or2_1 _09801_ (.X(_03848_),
    .B(_03846_),
    .A(_03756_));
 sg13g2_xnor2_1 _09802_ (.Y(_03849_),
    .A(_03755_),
    .B(_03847_));
 sg13g2_xor2_1 _09803_ (.B(_03849_),
    .A(_03845_),
    .X(_03850_));
 sg13g2_nand2_1 _09804_ (.Y(_03851_),
    .A(_03844_),
    .B(_03850_));
 sg13g2_xnor2_1 _09805_ (.Y(_03852_),
    .A(_03844_),
    .B(_03850_));
 sg13g2_xnor2_1 _09806_ (.Y(_03853_),
    .A(_03843_),
    .B(_03852_));
 sg13g2_xor2_1 _09807_ (.B(_03853_),
    .A(_03841_),
    .X(_03854_));
 sg13g2_nand2_1 _09808_ (.Y(_03855_),
    .A(_03824_),
    .B(_03854_));
 sg13g2_xnor2_1 _09809_ (.Y(_03856_),
    .A(_03824_),
    .B(_03854_));
 sg13g2_a21oi_1 _09810_ (.A1(_03774_),
    .A2(_03780_),
    .Y(_03857_),
    .B1(_03782_));
 sg13g2_o21ai_1 _09811_ (.B1(_03760_),
    .Y(_03858_),
    .A1(_03752_),
    .A2(_03761_));
 sg13g2_nand2_1 _09812_ (.Y(_03859_),
    .A(net1566),
    .B(net1710));
 sg13g2_nand2_1 _09813_ (.Y(_03860_),
    .A(net1571),
    .B(net1701));
 sg13g2_nand2_1 _09814_ (.Y(_03861_),
    .A(net1574),
    .B(net1701));
 sg13g2_xor2_1 _09815_ (.B(_03861_),
    .A(_03769_),
    .X(_03862_));
 sg13g2_nand2b_1 _09816_ (.Y(_03863_),
    .B(_03862_),
    .A_N(_03859_));
 sg13g2_xnor2_1 _09817_ (.Y(_03864_),
    .A(_03859_),
    .B(_03862_));
 sg13g2_inv_1 _09818_ (.Y(_03865_),
    .A(_03864_));
 sg13g2_o21ai_1 _09819_ (.B1(_03779_),
    .Y(_03866_),
    .A1(_03604_),
    .A2(_03777_));
 sg13g2_nand2_1 _09820_ (.Y(_03867_),
    .A(net1580),
    .B(net1696));
 sg13g2_nand2_1 _09821_ (.Y(_03868_),
    .A(net1586),
    .B(net1687));
 sg13g2_nand2_1 _09822_ (.Y(_03869_),
    .A(net1592),
    .B(net1687));
 sg13g2_xor2_1 _09823_ (.B(_03869_),
    .A(_03776_),
    .X(_03870_));
 sg13g2_nand2b_1 _09824_ (.Y(_03871_),
    .B(_03870_),
    .A_N(_03867_));
 sg13g2_xnor2_1 _09825_ (.Y(_03872_),
    .A(_03867_),
    .B(_03870_));
 sg13g2_nand2_1 _09826_ (.Y(_03873_),
    .A(_03866_),
    .B(_03872_));
 sg13g2_xnor2_1 _09827_ (.Y(_03874_),
    .A(_03866_),
    .B(_03872_));
 sg13g2_xnor2_1 _09828_ (.Y(_03875_),
    .A(_03865_),
    .B(_03874_));
 sg13g2_nand2b_1 _09829_ (.Y(_03876_),
    .B(_03858_),
    .A_N(_03875_));
 sg13g2_xor2_1 _09830_ (.B(_03875_),
    .A(_03858_),
    .X(_03877_));
 sg13g2_xnor2_1 _09831_ (.Y(_03878_),
    .A(_03857_),
    .B(_03877_));
 sg13g2_xor2_1 _09832_ (.B(_03878_),
    .A(_03856_),
    .X(_03879_));
 sg13g2_nand2_1 _09833_ (.Y(_03880_),
    .A(_03823_),
    .B(_03879_));
 sg13g2_xnor2_1 _09834_ (.Y(_03881_),
    .A(_03823_),
    .B(_03879_));
 sg13g2_o21ai_1 _09835_ (.B1(_03706_),
    .Y(_03882_),
    .A1(_03707_),
    .A2(_03725_));
 sg13g2_inv_1 _09836_ (.Y(_03883_),
    .A(_03882_));
 sg13g2_nand2_1 _09837_ (.Y(_03884_),
    .A(_03784_),
    .B(_03786_));
 sg13g2_a21o_1 _09838_ (.A2(_03702_),
    .A1(_03696_),
    .B1(_03704_),
    .X(_03885_));
 sg13g2_o21ai_1 _09839_ (.B1(_03700_),
    .Y(_03886_),
    .A1(_03697_),
    .A2(_03701_));
 sg13g2_inv_1 _09840_ (.Y(_03887_),
    .A(_03886_));
 sg13g2_o21ai_1 _09841_ (.B1(_03772_),
    .Y(_03888_),
    .A1(_03597_),
    .A2(_03770_));
 sg13g2_nand2_1 _09842_ (.Y(_03889_),
    .A(net1508),
    .B(net1728));
 sg13g2_nand2_1 _09843_ (.Y(_03890_),
    .A(net1510),
    .B(net1715));
 sg13g2_nand2_1 _09844_ (.Y(_03891_),
    .A(net1562),
    .B(net1715));
 sg13g2_or2_1 _09845_ (.X(_03892_),
    .B(_03890_),
    .A(_03699_));
 sg13g2_xnor2_1 _09846_ (.Y(_03893_),
    .A(_03698_),
    .B(_03891_));
 sg13g2_xor2_1 _09847_ (.B(_03893_),
    .A(_03889_),
    .X(_03894_));
 sg13g2_nand2_1 _09848_ (.Y(_03895_),
    .A(_03888_),
    .B(_03894_));
 sg13g2_xnor2_1 _09849_ (.Y(_03896_),
    .A(_03888_),
    .B(_03894_));
 sg13g2_xnor2_1 _09850_ (.Y(_03897_),
    .A(_03887_),
    .B(_03896_));
 sg13g2_nand2b_1 _09851_ (.Y(_03898_),
    .B(_03885_),
    .A_N(_03897_));
 sg13g2_xor2_1 _09852_ (.B(_03897_),
    .A(_03885_),
    .X(_03899_));
 sg13g2_nand2_2 _09853_ (.Y(_03900_),
    .A(net1487),
    .B(net1543));
 sg13g2_nand2_1 _09854_ (.Y(_03901_),
    .A(net1490),
    .B(net1532));
 sg13g2_nor2_1 _09855_ (.A(_03710_),
    .B(_03901_),
    .Y(_03902_));
 sg13g2_a22oi_1 _09856_ (.Y(_03903_),
    .B1(net1537),
    .B2(net1490),
    .A2(net1532),
    .A1(net1494));
 sg13g2_nor3_1 _09857_ (.A(_03900_),
    .B(_03902_),
    .C(_03903_),
    .Y(_03904_));
 sg13g2_o21ai_1 _09858_ (.B1(_03900_),
    .Y(_03905_),
    .A1(_03902_),
    .A2(_03903_));
 sg13g2_nand2b_1 _09859_ (.Y(_03906_),
    .B(_03905_),
    .A_N(_03904_));
 sg13g2_o21ai_1 _09860_ (.B1(_03720_),
    .Y(_03907_),
    .A1(_03559_),
    .A2(_03718_));
 sg13g2_nand2_1 _09861_ (.Y(_03908_),
    .A(net1498),
    .B(net1527));
 sg13g2_nand2_1 _09862_ (.Y(_03909_),
    .A(net1500),
    .B(net1514));
 sg13g2_nand2_1 _09863_ (.Y(_03910_),
    .A(net1504),
    .B(net1514));
 sg13g2_xor2_1 _09864_ (.B(_03910_),
    .A(_03717_),
    .X(_03911_));
 sg13g2_nand2b_1 _09865_ (.Y(_03912_),
    .B(_03911_),
    .A_N(_03908_));
 sg13g2_xnor2_1 _09866_ (.Y(_03913_),
    .A(_03908_),
    .B(_03911_));
 sg13g2_nand2_1 _09867_ (.Y(_03914_),
    .A(_03907_),
    .B(_03913_));
 sg13g2_xnor2_1 _09868_ (.Y(_03915_),
    .A(_03907_),
    .B(_03913_));
 sg13g2_xnor2_1 _09869_ (.Y(_03916_),
    .A(_03906_),
    .B(_03915_));
 sg13g2_xor2_1 _09870_ (.B(_03916_),
    .A(_03899_),
    .X(_03917_));
 sg13g2_nand2_1 _09871_ (.Y(_03918_),
    .A(_03884_),
    .B(_03917_));
 sg13g2_xnor2_1 _09872_ (.Y(_03919_),
    .A(_03884_),
    .B(_03917_));
 sg13g2_xnor2_1 _09873_ (.Y(_03920_),
    .A(_03883_),
    .B(_03919_));
 sg13g2_xor2_1 _09874_ (.B(_03920_),
    .A(_03881_),
    .X(_03921_));
 sg13g2_nand2_1 _09875_ (.Y(_03922_),
    .A(_03822_),
    .B(_03921_));
 sg13g2_xnor2_1 _09876_ (.Y(_03923_),
    .A(_03822_),
    .B(_03921_));
 sg13g2_xor2_1 _09877_ (.B(_03923_),
    .A(_03821_),
    .X(_03924_));
 sg13g2_and2_1 _09878_ (.A(_03806_),
    .B(_03924_),
    .X(_03925_));
 sg13g2_xnor2_1 _09879_ (.Y(_03926_),
    .A(_03806_),
    .B(_03924_));
 sg13g2_nor2_1 _09880_ (.A(_03689_),
    .B(_03926_),
    .Y(_03927_));
 sg13g2_xor2_1 _09881_ (.B(_03926_),
    .A(_03689_),
    .X(_03928_));
 sg13g2_o21ai_1 _09882_ (.B1(_03795_),
    .Y(_03929_),
    .A1(_03552_),
    .A2(_03796_));
 sg13g2_nand2_1 _09883_ (.Y(_03930_),
    .A(_03928_),
    .B(_03929_));
 sg13g2_xor2_1 _09884_ (.B(_03929_),
    .A(_03928_),
    .X(_03931_));
 sg13g2_nor2b_1 _09885_ (.A(_03798_),
    .B_N(_03931_),
    .Y(_03932_));
 sg13g2_xnor2_1 _09886_ (.Y(_03933_),
    .A(_03798_),
    .B(_03931_));
 sg13g2_xnor2_1 _09887_ (.Y(_03934_),
    .A(_03805_),
    .B(_03933_));
 sg13g2_o21ai_1 _09888_ (.B1(net1758),
    .Y(_03935_),
    .A1(net1398),
    .A2(_03934_));
 sg13g2_a21oi_1 _09889_ (.A1(net1399),
    .A2(_05547_),
    .Y(_00325_),
    .B1(_03935_));
 sg13g2_a21oi_1 _09890_ (.A1(_03687_),
    .A2(_03819_),
    .Y(_03936_),
    .B1(_03818_));
 sg13g2_o21ai_1 _09891_ (.B1(_03922_),
    .Y(_03937_),
    .A1(_03821_),
    .A2(_03923_));
 sg13g2_o21ai_1 _09892_ (.B1(_03880_),
    .Y(_03938_),
    .A1(_03881_),
    .A2(_03920_));
 sg13g2_o21ai_1 _09893_ (.B1(_03855_),
    .Y(_03939_),
    .A1(_03856_),
    .A2(_03878_));
 sg13g2_o21ai_1 _09894_ (.B1(_03840_),
    .Y(_03940_),
    .A1(_03841_),
    .A2(_03853_));
 sg13g2_o21ai_1 _09895_ (.B1(_03836_),
    .Y(_03941_),
    .A1(_03832_),
    .A2(_03838_));
 sg13g2_a21oi_2 _09896_ (.B1(_03837_),
    .Y(_03942_),
    .A2(_03834_),
    .A1(_03735_));
 sg13g2_nand2_1 _09897_ (.Y(_03943_),
    .A(net1612),
    .B(net1663));
 sg13g2_and2_1 _09898_ (.A(net1624),
    .B(net1657),
    .X(_03944_));
 sg13g2_nand2b_1 _09899_ (.Y(_03945_),
    .B(_03944_),
    .A_N(_03827_));
 sg13g2_xnor2_1 _09900_ (.Y(_03946_),
    .A(_03827_),
    .B(_03944_));
 sg13g2_nand2b_1 _09901_ (.Y(_03947_),
    .B(_03946_),
    .A_N(_03943_));
 sg13g2_xnor2_1 _09902_ (.Y(_03948_),
    .A(_03943_),
    .B(_03946_));
 sg13g2_xnor2_1 _09903_ (.Y(_03949_),
    .A(_03942_),
    .B(_03948_));
 sg13g2_nor2b_1 _09904_ (.A(_03949_),
    .B_N(_03941_),
    .Y(_03950_));
 sg13g2_nand2b_1 _09905_ (.Y(_03951_),
    .B(_03949_),
    .A_N(_03941_));
 sg13g2_nand2b_1 _09906_ (.Y(_03952_),
    .B(_03951_),
    .A_N(_03950_));
 sg13g2_o21ai_1 _09907_ (.B1(_03848_),
    .Y(_03953_),
    .A1(_03845_),
    .A2(_03849_));
 sg13g2_and2_1 _09908_ (.A(_03829_),
    .B(_03831_),
    .X(_03954_));
 sg13g2_nand2_1 _09909_ (.Y(_03955_),
    .A(net1598),
    .B(net1675));
 sg13g2_nand2_1 _09910_ (.Y(_03956_),
    .A(net1603),
    .B(net1669));
 sg13g2_nand2_1 _09911_ (.Y(_03957_),
    .A(net1607),
    .B(net1669));
 sg13g2_or2_1 _09912_ (.X(_03958_),
    .B(_03956_),
    .A(_03847_));
 sg13g2_xnor2_1 _09913_ (.Y(_03959_),
    .A(_03846_),
    .B(_03957_));
 sg13g2_xor2_1 _09914_ (.B(_03959_),
    .A(_03955_),
    .X(_03960_));
 sg13g2_nor2b_1 _09915_ (.A(_03954_),
    .B_N(_03960_),
    .Y(_03961_));
 sg13g2_xnor2_1 _09916_ (.Y(_03962_),
    .A(_03954_),
    .B(_03960_));
 sg13g2_xor2_1 _09917_ (.B(_03962_),
    .A(_03953_),
    .X(_03963_));
 sg13g2_xnor2_1 _09918_ (.Y(_03964_),
    .A(_03952_),
    .B(_03963_));
 sg13g2_nand2_1 _09919_ (.Y(_03965_),
    .A(_03940_),
    .B(_03964_));
 sg13g2_xnor2_1 _09920_ (.Y(_03966_),
    .A(_03940_),
    .B(_03964_));
 sg13g2_o21ai_1 _09921_ (.B1(_03873_),
    .Y(_03967_),
    .A1(_03865_),
    .A2(_03874_));
 sg13g2_o21ai_1 _09922_ (.B1(_03851_),
    .Y(_03968_),
    .A1(_03843_),
    .A2(_03852_));
 sg13g2_nand2_1 _09923_ (.Y(_03969_),
    .A(net1567),
    .B(net1704));
 sg13g2_nand2_1 _09924_ (.Y(_03970_),
    .A(net1570),
    .B(net1696));
 sg13g2_nand2_1 _09925_ (.Y(_03971_),
    .A(net1574),
    .B(net1696));
 sg13g2_xor2_1 _09926_ (.B(_03971_),
    .A(_03860_),
    .X(_03972_));
 sg13g2_nand2b_1 _09927_ (.Y(_03973_),
    .B(_03972_),
    .A_N(_03969_));
 sg13g2_xnor2_1 _09928_ (.Y(_03974_),
    .A(_03969_),
    .B(_03972_));
 sg13g2_inv_1 _09929_ (.Y(_03975_),
    .A(_03974_));
 sg13g2_o21ai_1 _09930_ (.B1(_03871_),
    .Y(_03976_),
    .A1(_03776_),
    .A2(_03869_));
 sg13g2_nand2_1 _09931_ (.Y(_03977_),
    .A(net1580),
    .B(net1691));
 sg13g2_nand2_1 _09932_ (.Y(_03978_),
    .A(net1586),
    .B(net1682));
 sg13g2_nand2_1 _09933_ (.Y(_03979_),
    .A(net1593),
    .B(net1682));
 sg13g2_xor2_1 _09934_ (.B(_03979_),
    .A(_03868_),
    .X(_03980_));
 sg13g2_nand2b_1 _09935_ (.Y(_03981_),
    .B(_03980_),
    .A_N(_03977_));
 sg13g2_xnor2_1 _09936_ (.Y(_03982_),
    .A(_03977_),
    .B(_03980_));
 sg13g2_nand2_1 _09937_ (.Y(_03983_),
    .A(_03976_),
    .B(_03982_));
 sg13g2_xnor2_1 _09938_ (.Y(_03984_),
    .A(_03976_),
    .B(_03982_));
 sg13g2_xnor2_1 _09939_ (.Y(_03985_),
    .A(_03975_),
    .B(_03984_));
 sg13g2_nand2b_1 _09940_ (.Y(_03986_),
    .B(_03968_),
    .A_N(_03985_));
 sg13g2_xor2_1 _09941_ (.B(_03985_),
    .A(_03968_),
    .X(_03987_));
 sg13g2_nand2b_1 _09942_ (.Y(_03988_),
    .B(_03967_),
    .A_N(_03987_));
 sg13g2_xor2_1 _09943_ (.B(_03987_),
    .A(_03967_),
    .X(_03989_));
 sg13g2_xor2_1 _09944_ (.B(_03989_),
    .A(_03966_),
    .X(_03990_));
 sg13g2_nand2_1 _09945_ (.Y(_03991_),
    .A(_03939_),
    .B(_03990_));
 sg13g2_xnor2_1 _09946_ (.Y(_03992_),
    .A(_03939_),
    .B(_03990_));
 sg13g2_o21ai_1 _09947_ (.B1(_03898_),
    .Y(_03993_),
    .A1(_03899_),
    .A2(_03916_));
 sg13g2_o21ai_1 _09948_ (.B1(_03876_),
    .Y(_03994_),
    .A1(_03857_),
    .A2(_03877_));
 sg13g2_o21ai_1 _09949_ (.B1(_03895_),
    .Y(_03995_),
    .A1(_03887_),
    .A2(_03896_));
 sg13g2_o21ai_1 _09950_ (.B1(_03892_),
    .Y(_03996_),
    .A1(_03889_),
    .A2(_03893_));
 sg13g2_o21ai_1 _09951_ (.B1(_03863_),
    .Y(_03997_),
    .A1(_03769_),
    .A2(_03861_));
 sg13g2_nand2_1 _09952_ (.Y(_03998_),
    .A(net1508),
    .B(net1721));
 sg13g2_nand2_1 _09953_ (.Y(_03999_),
    .A(net1510),
    .B(net1710));
 sg13g2_nand2_1 _09954_ (.Y(_04000_),
    .A(net1562),
    .B(net1710));
 sg13g2_or2_1 _09955_ (.X(_04001_),
    .B(_03999_),
    .A(_03891_));
 sg13g2_xnor2_1 _09956_ (.Y(_04002_),
    .A(_03890_),
    .B(_04000_));
 sg13g2_xor2_1 _09957_ (.B(_04002_),
    .A(_03998_),
    .X(_04003_));
 sg13g2_xnor2_1 _09958_ (.Y(_04004_),
    .A(_03997_),
    .B(_04003_));
 sg13g2_nor2b_1 _09959_ (.A(_04004_),
    .B_N(_03996_),
    .Y(_04005_));
 sg13g2_xor2_1 _09960_ (.B(_04004_),
    .A(_03996_),
    .X(_04006_));
 sg13g2_nand2b_1 _09961_ (.Y(_04007_),
    .B(_03995_),
    .A_N(_04006_));
 sg13g2_xor2_1 _09962_ (.B(_04006_),
    .A(_03995_),
    .X(_04008_));
 sg13g2_and2_1 _09963_ (.A(net1487),
    .B(net1537),
    .X(_04009_));
 sg13g2_nand2_1 _09964_ (.Y(_04010_),
    .A(net1487),
    .B(net1537));
 sg13g2_nand2_1 _09965_ (.Y(_04011_),
    .A(net1494),
    .B(net1530));
 sg13g2_xor2_1 _09966_ (.B(_04011_),
    .A(_03901_),
    .X(_04012_));
 sg13g2_nand2_1 _09967_ (.Y(_04013_),
    .A(_04009_),
    .B(_04012_));
 sg13g2_xnor2_1 _09968_ (.Y(_04014_),
    .A(_04009_),
    .B(_04012_));
 sg13g2_o21ai_1 _09969_ (.B1(_03912_),
    .Y(_04015_),
    .A1(_03717_),
    .A2(_03910_));
 sg13g2_nand2_1 _09970_ (.Y(_04016_),
    .A(net1498),
    .B(net1519));
 sg13g2_nand2_1 _09971_ (.Y(_04017_),
    .A(net1500),
    .B(net1728));
 sg13g2_nand2_1 _09972_ (.Y(_04018_),
    .A(net1504),
    .B(net1728));
 sg13g2_xor2_1 _09973_ (.B(_04018_),
    .A(_03909_),
    .X(_04019_));
 sg13g2_nand2b_1 _09974_ (.Y(_04020_),
    .B(_04019_),
    .A_N(_04016_));
 sg13g2_xnor2_1 _09975_ (.Y(_04021_),
    .A(_04016_),
    .B(_04019_));
 sg13g2_nand2_1 _09976_ (.Y(_04022_),
    .A(_04015_),
    .B(_04021_));
 sg13g2_xnor2_1 _09977_ (.Y(_04023_),
    .A(_04015_),
    .B(_04021_));
 sg13g2_xnor2_1 _09978_ (.Y(_04024_),
    .A(_04014_),
    .B(_04023_));
 sg13g2_xor2_1 _09979_ (.B(_04024_),
    .A(_04008_),
    .X(_04025_));
 sg13g2_xnor2_1 _09980_ (.Y(_04026_),
    .A(_03994_),
    .B(_04025_));
 sg13g2_nor2b_1 _09981_ (.A(_04026_),
    .B_N(_03993_),
    .Y(_04027_));
 sg13g2_xor2_1 _09982_ (.B(_04026_),
    .A(_03993_),
    .X(_04028_));
 sg13g2_xor2_1 _09983_ (.B(_04028_),
    .A(_03992_),
    .X(_04029_));
 sg13g2_nand2_1 _09984_ (.Y(_04030_),
    .A(_03938_),
    .B(_04029_));
 sg13g2_xnor2_1 _09985_ (.Y(_04031_),
    .A(_03938_),
    .B(_04029_));
 sg13g2_and3_1 _09986_ (.X(_04032_),
    .A(_03684_),
    .B(_03813_),
    .C(_03814_));
 sg13g2_inv_1 _09987_ (.Y(_04033_),
    .A(_04032_));
 sg13g2_o21ai_1 _09988_ (.B1(_03918_),
    .Y(_04034_),
    .A1(_03883_),
    .A2(_03919_));
 sg13g2_o21ai_1 _09989_ (.B1(_03914_),
    .Y(_04035_),
    .A1(_03906_),
    .A2(_03915_));
 sg13g2_or2_1 _09990_ (.X(_04036_),
    .B(_03904_),
    .A(_03902_));
 sg13g2_o21ai_1 _09991_ (.B1(net1488),
    .Y(_04037_),
    .A1(net1543),
    .A2(net1549));
 sg13g2_nor2_2 _09992_ (.A(_05573_),
    .B(_03709_),
    .Y(_04038_));
 sg13g2_nor2_1 _09993_ (.A(_03567_),
    .B(_04038_),
    .Y(_04039_));
 sg13g2_nor2_1 _09994_ (.A(_04037_),
    .B(_04038_),
    .Y(_04040_));
 sg13g2_xnor2_1 _09995_ (.Y(_04041_),
    .A(_03567_),
    .B(_04040_));
 sg13g2_inv_1 _09996_ (.Y(_04042_),
    .A(_04041_));
 sg13g2_nand2_1 _09997_ (.Y(_04043_),
    .A(_04036_),
    .B(_04041_));
 sg13g2_xnor2_1 _09998_ (.Y(_04044_),
    .A(_04036_),
    .B(_04041_));
 sg13g2_xnor2_1 _09999_ (.Y(_04045_),
    .A(_03807_),
    .B(_04044_));
 sg13g2_nand2_1 _10000_ (.Y(_04046_),
    .A(_04035_),
    .B(_04045_));
 sg13g2_xnor2_1 _10001_ (.Y(_04047_),
    .A(_04035_),
    .B(_04045_));
 sg13g2_xor2_1 _10002_ (.B(_04047_),
    .A(_03811_),
    .X(_04048_));
 sg13g2_nand2_1 _10003_ (.Y(_04049_),
    .A(_03682_),
    .B(_03814_));
 sg13g2_nand2_1 _10004_ (.Y(_04050_),
    .A(_03813_),
    .B(_04049_));
 sg13g2_nand2_1 _10005_ (.Y(_04051_),
    .A(_04048_),
    .B(_04050_));
 sg13g2_xor2_1 _10006_ (.B(_04050_),
    .A(_04048_),
    .X(_04052_));
 sg13g2_nand2_1 _10007_ (.Y(_04053_),
    .A(_04034_),
    .B(_04052_));
 sg13g2_xnor2_1 _10008_ (.Y(_04054_),
    .A(_04034_),
    .B(_04052_));
 sg13g2_xnor2_1 _10009_ (.Y(_04055_),
    .A(_04033_),
    .B(_04054_));
 sg13g2_xor2_1 _10010_ (.B(_04055_),
    .A(_04031_),
    .X(_04056_));
 sg13g2_nand2_1 _10011_ (.Y(_04057_),
    .A(_03937_),
    .B(_04056_));
 sg13g2_xnor2_1 _10012_ (.Y(_04058_),
    .A(_03937_),
    .B(_04056_));
 sg13g2_xor2_1 _10013_ (.B(_04058_),
    .A(_03936_),
    .X(_04059_));
 sg13g2_o21ai_1 _10014_ (.B1(_04059_),
    .Y(_04060_),
    .A1(_03925_),
    .A2(_03927_));
 sg13g2_or3_1 _10015_ (.A(_03925_),
    .B(_03927_),
    .C(_04059_),
    .X(_04061_));
 sg13g2_and2_1 _10016_ (.A(_04060_),
    .B(_04061_),
    .X(_04062_));
 sg13g2_nor2b_1 _10017_ (.A(_03930_),
    .B_N(_04062_),
    .Y(_04063_));
 sg13g2_xnor2_1 _10018_ (.Y(_04064_),
    .A(_03930_),
    .B(_04062_));
 sg13g2_and2_1 _10019_ (.A(_03802_),
    .B(_03933_),
    .X(_04065_));
 sg13g2_a21o_1 _10020_ (.A2(_03933_),
    .A1(_03800_),
    .B1(_03932_),
    .X(_04066_));
 sg13g2_a21o_2 _10021_ (.A2(_04065_),
    .A1(_03678_),
    .B1(_04066_),
    .X(_04067_));
 sg13g2_xor2_1 _10022_ (.B(_04067_),
    .A(_04064_),
    .X(_04068_));
 sg13g2_o21ai_1 _10023_ (.B1(net1757),
    .Y(_04069_),
    .A1(net1398),
    .A2(_04068_));
 sg13g2_a21oi_1 _10024_ (.A1(net1398),
    .A2(_05546_),
    .Y(_00326_),
    .B1(_04069_));
 sg13g2_o21ai_1 _10025_ (.B1(_04053_),
    .Y(_04070_),
    .A1(_04033_),
    .A2(_04054_));
 sg13g2_o21ai_1 _10026_ (.B1(_04030_),
    .Y(_04071_),
    .A1(_04031_),
    .A2(_04055_));
 sg13g2_o21ai_1 _10027_ (.B1(_03991_),
    .Y(_04072_),
    .A1(_03992_),
    .A2(_04028_));
 sg13g2_o21ai_1 _10028_ (.B1(_03965_),
    .Y(_04073_),
    .A1(_03966_),
    .A2(_03989_));
 sg13g2_a21o_1 _10029_ (.A2(_03963_),
    .A1(_03951_),
    .B1(_03950_),
    .X(_04074_));
 sg13g2_a21o_1 _10030_ (.A2(_03948_),
    .A1(_03942_),
    .B1(_03837_),
    .X(_04075_));
 sg13g2_o21ai_1 _10031_ (.B1(net1657),
    .Y(_04076_),
    .A1(net1616),
    .A2(net1624));
 sg13g2_a21o_2 _10032_ (.A2(_03944_),
    .A1(net1616),
    .B1(_04076_),
    .X(_04077_));
 sg13g2_nand2_1 _10033_ (.Y(_04078_),
    .A(net1612),
    .B(net1660));
 sg13g2_nor2_1 _10034_ (.A(_04077_),
    .B(_04078_),
    .Y(_04079_));
 sg13g2_xor2_1 _10035_ (.B(_04078_),
    .A(_04077_),
    .X(_04080_));
 sg13g2_xor2_1 _10036_ (.B(_04080_),
    .A(_03942_),
    .X(_04081_));
 sg13g2_nand2_1 _10037_ (.Y(_04082_),
    .A(_04075_),
    .B(_04081_));
 sg13g2_xnor2_1 _10038_ (.Y(_04083_),
    .A(_04075_),
    .B(_04081_));
 sg13g2_o21ai_1 _10039_ (.B1(_03958_),
    .Y(_04084_),
    .A1(_03955_),
    .A2(_03959_));
 sg13g2_and2_1 _10040_ (.A(_03945_),
    .B(_03947_),
    .X(_04085_));
 sg13g2_nand2_1 _10041_ (.Y(_04086_),
    .A(net1598),
    .B(net1673));
 sg13g2_nand2_2 _10042_ (.Y(_04087_),
    .A(net1603),
    .B(net1663));
 sg13g2_nand2_1 _10043_ (.Y(_04088_),
    .A(net1607),
    .B(net1663));
 sg13g2_or2_1 _10044_ (.X(_04089_),
    .B(_04087_),
    .A(_03957_));
 sg13g2_xnor2_1 _10045_ (.Y(_04090_),
    .A(_03956_),
    .B(_04088_));
 sg13g2_xor2_1 _10046_ (.B(_04090_),
    .A(_04086_),
    .X(_04091_));
 sg13g2_nor2b_1 _10047_ (.A(_04085_),
    .B_N(_04091_),
    .Y(_04092_));
 sg13g2_xnor2_1 _10048_ (.Y(_04093_),
    .A(_04085_),
    .B(_04091_));
 sg13g2_xnor2_1 _10049_ (.Y(_04094_),
    .A(_04084_),
    .B(_04093_));
 sg13g2_xor2_1 _10050_ (.B(_04094_),
    .A(_04083_),
    .X(_04095_));
 sg13g2_and2_1 _10051_ (.A(_04074_),
    .B(_04095_),
    .X(_04096_));
 sg13g2_or2_1 _10052_ (.X(_04097_),
    .B(_04095_),
    .A(_04074_));
 sg13g2_nand2b_1 _10053_ (.Y(_04098_),
    .B(_04097_),
    .A_N(_04096_));
 sg13g2_o21ai_1 _10054_ (.B1(_03983_),
    .Y(_04099_),
    .A1(_03975_),
    .A2(_03984_));
 sg13g2_a21o_1 _10055_ (.A2(_03962_),
    .A1(_03953_),
    .B1(_03961_),
    .X(_04100_));
 sg13g2_nand2_1 _10056_ (.Y(_04101_),
    .A(net1566),
    .B(net1701));
 sg13g2_nand2_1 _10057_ (.Y(_04102_),
    .A(net1570),
    .B(net1692));
 sg13g2_nand2_1 _10058_ (.Y(_04103_),
    .A(net1574),
    .B(net1692));
 sg13g2_xor2_1 _10059_ (.B(_04103_),
    .A(_03970_),
    .X(_04104_));
 sg13g2_nand2b_1 _10060_ (.Y(_04105_),
    .B(_04104_),
    .A_N(_04101_));
 sg13g2_xnor2_1 _10061_ (.Y(_04106_),
    .A(_04101_),
    .B(_04104_));
 sg13g2_inv_1 _10062_ (.Y(_04107_),
    .A(_04106_));
 sg13g2_o21ai_1 _10063_ (.B1(_03981_),
    .Y(_04108_),
    .A1(_03868_),
    .A2(_03979_));
 sg13g2_nand2_1 _10064_ (.Y(_04109_),
    .A(net1580),
    .B(net1687));
 sg13g2_nand2_1 _10065_ (.Y(_04110_),
    .A(net1584),
    .B(net1677));
 sg13g2_nand2_1 _10066_ (.Y(_04111_),
    .A(net1593),
    .B(net1677));
 sg13g2_xor2_1 _10067_ (.B(_04111_),
    .A(_03978_),
    .X(_04112_));
 sg13g2_nand2b_1 _10068_ (.Y(_04113_),
    .B(_04112_),
    .A_N(_04109_));
 sg13g2_xnor2_1 _10069_ (.Y(_04114_),
    .A(_04109_),
    .B(_04112_));
 sg13g2_nand2_1 _10070_ (.Y(_04115_),
    .A(_04108_),
    .B(_04114_));
 sg13g2_xnor2_1 _10071_ (.Y(_04116_),
    .A(_04108_),
    .B(_04114_));
 sg13g2_xnor2_1 _10072_ (.Y(_04117_),
    .A(_04106_),
    .B(_04116_));
 sg13g2_xnor2_1 _10073_ (.Y(_04118_),
    .A(_04100_),
    .B(_04117_));
 sg13g2_nor2b_1 _10074_ (.A(_04118_),
    .B_N(_04099_),
    .Y(_04119_));
 sg13g2_xnor2_1 _10075_ (.Y(_04120_),
    .A(_04099_),
    .B(_04118_));
 sg13g2_xnor2_1 _10076_ (.Y(_04121_),
    .A(_04098_),
    .B(_04120_));
 sg13g2_nand2_1 _10077_ (.Y(_04122_),
    .A(_04073_),
    .B(_04121_));
 sg13g2_xnor2_1 _10078_ (.Y(_04123_),
    .A(_04073_),
    .B(_04121_));
 sg13g2_o21ai_1 _10079_ (.B1(_04007_),
    .Y(_04124_),
    .A1(_04008_),
    .A2(_04024_));
 sg13g2_nand2_2 _10080_ (.Y(_04125_),
    .A(_03986_),
    .B(_03988_));
 sg13g2_a21o_1 _10081_ (.A2(_04003_),
    .A1(_03997_),
    .B1(_04005_),
    .X(_04126_));
 sg13g2_o21ai_1 _10082_ (.B1(_04001_),
    .Y(_04127_),
    .A1(_03998_),
    .A2(_04002_));
 sg13g2_o21ai_1 _10083_ (.B1(_03973_),
    .Y(_04128_),
    .A1(_03860_),
    .A2(_03971_));
 sg13g2_nand2_1 _10084_ (.Y(_04129_),
    .A(net1508),
    .B(net1715));
 sg13g2_nand2_1 _10085_ (.Y(_04130_),
    .A(net1510),
    .B(net1704));
 sg13g2_nand2_1 _10086_ (.Y(_04131_),
    .A(net1562),
    .B(net1704));
 sg13g2_or2_1 _10087_ (.X(_04132_),
    .B(_04130_),
    .A(_04000_));
 sg13g2_xnor2_1 _10088_ (.Y(_04133_),
    .A(_03999_),
    .B(_04131_));
 sg13g2_xor2_1 _10089_ (.B(_04133_),
    .A(_04129_),
    .X(_04134_));
 sg13g2_xnor2_1 _10090_ (.Y(_04135_),
    .A(_04128_),
    .B(_04134_));
 sg13g2_nor2b_1 _10091_ (.A(_04135_),
    .B_N(_04127_),
    .Y(_04136_));
 sg13g2_xor2_1 _10092_ (.B(_04135_),
    .A(_04127_),
    .X(_04137_));
 sg13g2_nand2b_1 _10093_ (.Y(_04138_),
    .B(_04126_),
    .A_N(_04137_));
 sg13g2_xor2_1 _10094_ (.B(_04137_),
    .A(_04126_),
    .X(_04139_));
 sg13g2_and2_1 _10095_ (.A(net1487),
    .B(net1532),
    .X(_04140_));
 sg13g2_nand2_1 _10096_ (.Y(_04141_),
    .A(net1487),
    .B(net1532));
 sg13g2_nand2_1 _10097_ (.Y(_04142_),
    .A(net1493),
    .B(net1519));
 sg13g2_nor3_1 _10098_ (.A(_05552_),
    .B(_05571_),
    .C(_04142_),
    .Y(_04143_));
 sg13g2_a22oi_1 _10099_ (.Y(_04144_),
    .B1(net1527),
    .B2(net1490),
    .A2(net1519),
    .A1(net1493));
 sg13g2_nor2_1 _10100_ (.A(_04143_),
    .B(_04144_),
    .Y(_04145_));
 sg13g2_xnor2_1 _10101_ (.Y(_04146_),
    .A(_04141_),
    .B(_04145_));
 sg13g2_inv_1 _10102_ (.Y(_04147_),
    .A(_04146_));
 sg13g2_o21ai_1 _10103_ (.B1(_04020_),
    .Y(_04148_),
    .A1(_03909_),
    .A2(_04018_));
 sg13g2_nand2_1 _10104_ (.Y(_04149_),
    .A(net1498),
    .B(net1514));
 sg13g2_nand2_1 _10105_ (.Y(_04150_),
    .A(net1501),
    .B(net1721));
 sg13g2_nand2_1 _10106_ (.Y(_04151_),
    .A(net1504),
    .B(net1721));
 sg13g2_xor2_1 _10107_ (.B(_04151_),
    .A(_04017_),
    .X(_04152_));
 sg13g2_nand2b_1 _10108_ (.Y(_04153_),
    .B(_04152_),
    .A_N(_04149_));
 sg13g2_xnor2_1 _10109_ (.Y(_04154_),
    .A(_04149_),
    .B(_04152_));
 sg13g2_nand2_1 _10110_ (.Y(_04155_),
    .A(_04148_),
    .B(_04154_));
 sg13g2_xnor2_1 _10111_ (.Y(_04156_),
    .A(_04148_),
    .B(_04154_));
 sg13g2_xnor2_1 _10112_ (.Y(_04157_),
    .A(_04147_),
    .B(_04156_));
 sg13g2_xor2_1 _10113_ (.B(_04157_),
    .A(_04139_),
    .X(_04158_));
 sg13g2_xnor2_1 _10114_ (.Y(_04159_),
    .A(_04125_),
    .B(_04158_));
 sg13g2_nor2b_1 _10115_ (.A(_04159_),
    .B_N(_04124_),
    .Y(_04160_));
 sg13g2_xor2_1 _10116_ (.B(_04159_),
    .A(_04124_),
    .X(_04161_));
 sg13g2_xor2_1 _10117_ (.B(_04161_),
    .A(_04123_),
    .X(_04162_));
 sg13g2_xnor2_1 _10118_ (.Y(_04163_),
    .A(_04072_),
    .B(_04162_));
 sg13g2_a21o_1 _10119_ (.A2(_04025_),
    .A1(_03994_),
    .B1(_04027_),
    .X(_04164_));
 sg13g2_o21ai_1 _10120_ (.B1(_04046_),
    .Y(_04165_),
    .A1(_03811_),
    .A2(_04047_));
 sg13g2_o21ai_1 _10121_ (.B1(_04043_),
    .Y(_04166_),
    .A1(_03808_),
    .A2(_04044_));
 sg13g2_o21ai_1 _10122_ (.B1(_04022_),
    .Y(_04167_),
    .A1(_04014_),
    .A2(_04023_));
 sg13g2_inv_1 _10123_ (.Y(_04168_),
    .A(_04167_));
 sg13g2_a21o_2 _10124_ (.A2(_04040_),
    .A1(_03566_),
    .B1(_04038_),
    .X(_04169_));
 sg13g2_o21ai_1 _10125_ (.B1(_04013_),
    .Y(_04170_),
    .A1(_03901_),
    .A2(_04011_));
 sg13g2_nand2_1 _10126_ (.Y(_04171_),
    .A(net1543),
    .B(_04009_));
 sg13g2_nand2_1 _10127_ (.Y(_04172_),
    .A(_03900_),
    .B(_04010_));
 sg13g2_nand2_1 _10128_ (.Y(_04173_),
    .A(_04171_),
    .B(_04172_));
 sg13g2_xnor2_1 _10129_ (.Y(_04174_),
    .A(_03708_),
    .B(_04173_));
 sg13g2_inv_1 _10130_ (.Y(_04175_),
    .A(_04174_));
 sg13g2_xnor2_1 _10131_ (.Y(_04176_),
    .A(_04170_),
    .B(_04174_));
 sg13g2_nor2b_1 _10132_ (.A(_04176_),
    .B_N(_04169_),
    .Y(_04177_));
 sg13g2_xor2_1 _10133_ (.B(_04176_),
    .A(_04169_),
    .X(_04178_));
 sg13g2_xor2_1 _10134_ (.B(_04178_),
    .A(_04167_),
    .X(_04179_));
 sg13g2_nand2b_1 _10135_ (.Y(_04180_),
    .B(_04166_),
    .A_N(_04179_));
 sg13g2_xnor2_1 _10136_ (.Y(_04181_),
    .A(_04166_),
    .B(_04179_));
 sg13g2_nand2_1 _10137_ (.Y(_04182_),
    .A(_04165_),
    .B(_04181_));
 sg13g2_xnor2_1 _10138_ (.Y(_04183_),
    .A(_04165_),
    .B(_04181_));
 sg13g2_xnor2_1 _10139_ (.Y(_04184_),
    .A(_03566_),
    .B(_04183_));
 sg13g2_nand2_1 _10140_ (.Y(_04185_),
    .A(_04164_),
    .B(_04184_));
 sg13g2_xnor2_1 _10141_ (.Y(_04186_),
    .A(_04164_),
    .B(_04184_));
 sg13g2_xor2_1 _10142_ (.B(_04186_),
    .A(_04051_),
    .X(_04187_));
 sg13g2_nor2b_1 _10143_ (.A(_04163_),
    .B_N(_04187_),
    .Y(_04188_));
 sg13g2_xnor2_1 _10144_ (.Y(_04189_),
    .A(_04163_),
    .B(_04187_));
 sg13g2_xnor2_1 _10145_ (.Y(_04190_),
    .A(_04071_),
    .B(_04189_));
 sg13g2_nor2b_1 _10146_ (.A(_04190_),
    .B_N(_04070_),
    .Y(_04191_));
 sg13g2_xnor2_1 _10147_ (.Y(_04192_),
    .A(_04070_),
    .B(_04190_));
 sg13g2_o21ai_1 _10148_ (.B1(_04057_),
    .Y(_04193_),
    .A1(_03936_),
    .A2(_04058_));
 sg13g2_nand2_1 _10149_ (.Y(_04194_),
    .A(_04192_),
    .B(_04193_));
 sg13g2_xnor2_1 _10150_ (.Y(_04195_),
    .A(_04192_),
    .B(_04193_));
 sg13g2_nand2_1 _10151_ (.Y(_04196_),
    .A(_04060_),
    .B(_04195_));
 sg13g2_nor2_1 _10152_ (.A(_04060_),
    .B(_04195_),
    .Y(_04197_));
 sg13g2_xor2_1 _10153_ (.B(_04195_),
    .A(_04060_),
    .X(_04198_));
 sg13g2_a21oi_1 _10154_ (.A1(_04064_),
    .A2(_04067_),
    .Y(_04199_),
    .B1(_04063_));
 sg13g2_xnor2_1 _10155_ (.Y(_04200_),
    .A(_04198_),
    .B(_04199_));
 sg13g2_o21ai_1 _10156_ (.B1(net1757),
    .Y(_04201_),
    .A1(net1398),
    .A2(_04200_));
 sg13g2_a21oi_1 _10157_ (.A1(net1399),
    .A2(_05545_),
    .Y(_00327_),
    .B1(_04201_));
 sg13g2_and2_1 _10158_ (.A(_04064_),
    .B(_04198_),
    .X(_04202_));
 sg13g2_a21o_1 _10159_ (.A2(_04196_),
    .A1(_04063_),
    .B1(_04197_),
    .X(_04203_));
 sg13g2_a21o_1 _10160_ (.A2(_04202_),
    .A1(_04067_),
    .B1(_04203_),
    .X(_04204_));
 sg13g2_o21ai_1 _10161_ (.B1(_04185_),
    .Y(_04205_),
    .A1(_04051_),
    .A2(_04186_));
 sg13g2_a21o_1 _10162_ (.A2(_04162_),
    .A1(_04072_),
    .B1(_04188_),
    .X(_04206_));
 sg13g2_o21ai_1 _10163_ (.B1(_04122_),
    .Y(_04207_),
    .A1(_04123_),
    .A2(_04161_));
 sg13g2_a21o_2 _10164_ (.A2(_04120_),
    .A1(_04097_),
    .B1(_04096_),
    .X(_04208_));
 sg13g2_o21ai_1 _10165_ (.B1(_04082_),
    .Y(_04209_),
    .A1(_04083_),
    .A2(_04094_));
 sg13g2_a21o_1 _10166_ (.A2(_04080_),
    .A1(_03942_),
    .B1(_03837_),
    .X(_04210_));
 sg13g2_nand2_1 _10167_ (.Y(_04211_),
    .A(net1612),
    .B(\cordic_inst.MUX_cordic_state$write_1__VAL_1[79] ));
 sg13g2_nor2_1 _10168_ (.A(_04077_),
    .B(_04211_),
    .Y(_04212_));
 sg13g2_xor2_1 _10169_ (.B(_04211_),
    .A(_04077_),
    .X(_04213_));
 sg13g2_xor2_1 _10170_ (.B(_04213_),
    .A(_03942_),
    .X(_04214_));
 sg13g2_nand2_1 _10171_ (.Y(_04215_),
    .A(_04210_),
    .B(_04214_));
 sg13g2_xnor2_1 _10172_ (.Y(_04216_),
    .A(_04210_),
    .B(_04214_));
 sg13g2_o21ai_1 _10173_ (.B1(_04089_),
    .Y(_04217_),
    .A1(_04086_),
    .A2(_04090_));
 sg13g2_a21oi_1 _10174_ (.A1(net1616),
    .A2(_03944_),
    .Y(_04218_),
    .B1(_04079_));
 sg13g2_nand2_1 _10175_ (.Y(_04219_),
    .A(net1601),
    .B(net1669));
 sg13g2_nand2_1 _10176_ (.Y(_04220_),
    .A(net1606),
    .B(net1658));
 sg13g2_nand2_1 _10177_ (.Y(_04221_),
    .A(net1608),
    .B(net1660));
 sg13g2_xnor2_1 _10178_ (.Y(_04222_),
    .A(_04087_),
    .B(_04221_));
 sg13g2_or2_1 _10179_ (.X(_04223_),
    .B(_04222_),
    .A(_04219_));
 sg13g2_xor2_1 _10180_ (.B(_04222_),
    .A(_04219_),
    .X(_04224_));
 sg13g2_nor2b_1 _10181_ (.A(_04218_),
    .B_N(_04224_),
    .Y(_04225_));
 sg13g2_xnor2_1 _10182_ (.Y(_04226_),
    .A(_04218_),
    .B(_04224_));
 sg13g2_xnor2_1 _10183_ (.Y(_04227_),
    .A(_04217_),
    .B(_04226_));
 sg13g2_xor2_1 _10184_ (.B(_04227_),
    .A(_04216_),
    .X(_04228_));
 sg13g2_nand2_1 _10185_ (.Y(_04229_),
    .A(_04209_),
    .B(_04228_));
 sg13g2_xnor2_1 _10186_ (.Y(_04230_),
    .A(_04209_),
    .B(_04228_));
 sg13g2_o21ai_1 _10187_ (.B1(_04115_),
    .Y(_04231_),
    .A1(_04107_),
    .A2(_04116_));
 sg13g2_inv_1 _10188_ (.Y(_04232_),
    .A(_04231_));
 sg13g2_a21o_1 _10189_ (.A2(_04093_),
    .A1(_04084_),
    .B1(_04092_),
    .X(_04233_));
 sg13g2_nand2_1 _10190_ (.Y(_04234_),
    .A(net1566),
    .B(net1697));
 sg13g2_nand2_1 _10191_ (.Y(_04235_),
    .A(net1572),
    .B(net1684));
 sg13g2_nand2_1 _10192_ (.Y(_04236_),
    .A(net1574),
    .B(net1687));
 sg13g2_xor2_1 _10193_ (.B(_04236_),
    .A(_04102_),
    .X(_04237_));
 sg13g2_nand2b_1 _10194_ (.Y(_04238_),
    .B(_04237_),
    .A_N(_04234_));
 sg13g2_xnor2_1 _10195_ (.Y(_04239_),
    .A(_04234_),
    .B(_04237_));
 sg13g2_inv_1 _10196_ (.Y(_04240_),
    .A(_04239_));
 sg13g2_o21ai_1 _10197_ (.B1(_04113_),
    .Y(_04241_),
    .A1(_03978_),
    .A2(_04111_));
 sg13g2_nand2_1 _10198_ (.Y(_04242_),
    .A(net1579),
    .B(net1682));
 sg13g2_nand2_1 _10199_ (.Y(_04243_),
    .A(net1584),
    .B(net1673));
 sg13g2_nand2_1 _10200_ (.Y(_04244_),
    .A(net1591),
    .B(net1673));
 sg13g2_xor2_1 _10201_ (.B(_04244_),
    .A(_04110_),
    .X(_04245_));
 sg13g2_nand2b_1 _10202_ (.Y(_04246_),
    .B(_04245_),
    .A_N(_04242_));
 sg13g2_xnor2_1 _10203_ (.Y(_04247_),
    .A(_04242_),
    .B(_04245_));
 sg13g2_nand2_1 _10204_ (.Y(_04248_),
    .A(_04241_),
    .B(_04247_));
 sg13g2_xnor2_1 _10205_ (.Y(_04249_),
    .A(_04241_),
    .B(_04247_));
 sg13g2_xnor2_1 _10206_ (.Y(_04250_),
    .A(_04240_),
    .B(_04249_));
 sg13g2_nand2b_1 _10207_ (.Y(_04251_),
    .B(_04233_),
    .A_N(_04250_));
 sg13g2_xor2_1 _10208_ (.B(_04250_),
    .A(_04233_),
    .X(_04252_));
 sg13g2_xnor2_1 _10209_ (.Y(_04253_),
    .A(_04232_),
    .B(_04252_));
 sg13g2_xor2_1 _10210_ (.B(_04253_),
    .A(_04230_),
    .X(_04254_));
 sg13g2_and2_1 _10211_ (.A(_04208_),
    .B(_04254_),
    .X(_04255_));
 sg13g2_or2_1 _10212_ (.X(_04256_),
    .B(_04254_),
    .A(_04208_));
 sg13g2_nand2b_1 _10213_ (.Y(_04257_),
    .B(_04256_),
    .A_N(_04255_));
 sg13g2_o21ai_1 _10214_ (.B1(_04138_),
    .Y(_04258_),
    .A1(_04139_),
    .A2(_04157_));
 sg13g2_a21o_2 _10215_ (.A2(_04117_),
    .A1(_04100_),
    .B1(_04119_),
    .X(_04259_));
 sg13g2_a21o_1 _10216_ (.A2(_04134_),
    .A1(_04128_),
    .B1(_04136_),
    .X(_04260_));
 sg13g2_o21ai_1 _10217_ (.B1(_04132_),
    .Y(_04261_),
    .A1(_04129_),
    .A2(_04133_));
 sg13g2_o21ai_1 _10218_ (.B1(_04105_),
    .Y(_04262_),
    .A1(_03970_),
    .A2(_04103_));
 sg13g2_nand2_1 _10219_ (.Y(_04263_),
    .A(net1509),
    .B(net1711));
 sg13g2_nand2_1 _10220_ (.Y(_04264_),
    .A(net1510),
    .B(net1702));
 sg13g2_nand2_1 _10221_ (.Y(_04265_),
    .A(net1562),
    .B(net1702));
 sg13g2_or2_1 _10222_ (.X(_04266_),
    .B(_04264_),
    .A(_04131_));
 sg13g2_xnor2_1 _10223_ (.Y(_04267_),
    .A(_04130_),
    .B(_04265_));
 sg13g2_xor2_1 _10224_ (.B(_04267_),
    .A(_04263_),
    .X(_04268_));
 sg13g2_xnor2_1 _10225_ (.Y(_04269_),
    .A(_04262_),
    .B(_04268_));
 sg13g2_nor2b_1 _10226_ (.A(_04269_),
    .B_N(_04261_),
    .Y(_04270_));
 sg13g2_xor2_1 _10227_ (.B(_04269_),
    .A(_04261_),
    .X(_04271_));
 sg13g2_nand2b_1 _10228_ (.Y(_04272_),
    .B(_04260_),
    .A_N(_04271_));
 sg13g2_xor2_1 _10229_ (.B(_04271_),
    .A(_04260_),
    .X(_04273_));
 sg13g2_and2_1 _10230_ (.A(net1488),
    .B(net1527),
    .X(_04274_));
 sg13g2_nand2_1 _10231_ (.Y(_04275_),
    .A(net1488),
    .B(net1527));
 sg13g2_nor3_1 _10232_ (.A(_05552_),
    .B(_05570_),
    .C(_04142_),
    .Y(_04276_));
 sg13g2_a22oi_1 _10233_ (.Y(_04277_),
    .B1(net1519),
    .B2(net1490),
    .A2(net1514),
    .A1(net1493));
 sg13g2_nor2_1 _10234_ (.A(_04276_),
    .B(_04277_),
    .Y(_04278_));
 sg13g2_xnor2_1 _10235_ (.Y(_04279_),
    .A(_04275_),
    .B(_04278_));
 sg13g2_inv_1 _10236_ (.Y(_04280_),
    .A(_04279_));
 sg13g2_o21ai_1 _10237_ (.B1(_04153_),
    .Y(_04281_),
    .A1(_04017_),
    .A2(_04151_));
 sg13g2_nand2_1 _10238_ (.Y(_04282_),
    .A(net1498),
    .B(net1728));
 sg13g2_nand2_1 _10239_ (.Y(_04283_),
    .A(net1500),
    .B(net1716));
 sg13g2_nand2_1 _10240_ (.Y(_04284_),
    .A(net1504),
    .B(net1715));
 sg13g2_xor2_1 _10241_ (.B(_04284_),
    .A(_04150_),
    .X(_04285_));
 sg13g2_nand2b_1 _10242_ (.Y(_04286_),
    .B(_04285_),
    .A_N(_04282_));
 sg13g2_xnor2_1 _10243_ (.Y(_04287_),
    .A(_04282_),
    .B(_04285_));
 sg13g2_nand2_1 _10244_ (.Y(_04288_),
    .A(_04281_),
    .B(_04287_));
 sg13g2_xnor2_1 _10245_ (.Y(_04289_),
    .A(_04281_),
    .B(_04287_));
 sg13g2_xnor2_1 _10246_ (.Y(_04290_),
    .A(_04280_),
    .B(_04289_));
 sg13g2_xor2_1 _10247_ (.B(_04290_),
    .A(_04273_),
    .X(_04291_));
 sg13g2_xnor2_1 _10248_ (.Y(_04292_),
    .A(_04259_),
    .B(_04291_));
 sg13g2_nor2b_1 _10249_ (.A(_04292_),
    .B_N(_04258_),
    .Y(_04293_));
 sg13g2_xnor2_1 _10250_ (.Y(_04294_),
    .A(_04258_),
    .B(_04292_));
 sg13g2_xnor2_1 _10251_ (.Y(_04295_),
    .A(_04257_),
    .B(_04294_));
 sg13g2_nand2_1 _10252_ (.Y(_04296_),
    .A(_04207_),
    .B(_04295_));
 sg13g2_xnor2_1 _10253_ (.Y(_04297_),
    .A(_04207_),
    .B(_04295_));
 sg13g2_o21ai_1 _10254_ (.B1(_04182_),
    .Y(_04298_),
    .A1(_03567_),
    .A2(_04183_));
 sg13g2_a21o_1 _10255_ (.A2(_04158_),
    .A1(_04125_),
    .B1(_04160_),
    .X(_04299_));
 sg13g2_o21ai_1 _10256_ (.B1(_04180_),
    .Y(_04300_),
    .A1(_04168_),
    .A2(_04178_));
 sg13g2_a21o_1 _10257_ (.A2(_04174_),
    .A1(_04170_),
    .B1(_04177_),
    .X(_04301_));
 sg13g2_o21ai_1 _10258_ (.B1(_04155_),
    .Y(_04302_),
    .A1(_04147_),
    .A2(_04156_));
 sg13g2_o21ai_1 _10259_ (.B1(_04171_),
    .Y(_04303_),
    .A1(_03709_),
    .A2(_04173_));
 sg13g2_a21o_1 _10260_ (.A2(_04145_),
    .A1(_04140_),
    .B1(_04143_),
    .X(_04304_));
 sg13g2_nand2_1 _10261_ (.Y(_04305_),
    .A(net1536),
    .B(_04009_));
 sg13g2_o21ai_1 _10262_ (.B1(_04305_),
    .Y(_04306_),
    .A1(_04009_),
    .A2(_04140_));
 sg13g2_xor2_1 _10263_ (.B(_04306_),
    .A(_03900_),
    .X(_04307_));
 sg13g2_inv_1 _10264_ (.Y(_04308_),
    .A(_04307_));
 sg13g2_xnor2_1 _10265_ (.Y(_04309_),
    .A(_04304_),
    .B(_04307_));
 sg13g2_nor2b_1 _10266_ (.A(_04309_),
    .B_N(_04303_),
    .Y(_04310_));
 sg13g2_xnor2_1 _10267_ (.Y(_04311_),
    .A(_04303_),
    .B(_04309_));
 sg13g2_xnor2_1 _10268_ (.Y(_04312_),
    .A(_04302_),
    .B(_04311_));
 sg13g2_nor2b_1 _10269_ (.A(_04312_),
    .B_N(_04301_),
    .Y(_04313_));
 sg13g2_xor2_1 _10270_ (.B(_04312_),
    .A(_04301_),
    .X(_04314_));
 sg13g2_nand2b_1 _10271_ (.Y(_04315_),
    .B(_04300_),
    .A_N(_04314_));
 sg13g2_xor2_1 _10272_ (.B(_04314_),
    .A(_04300_),
    .X(_04316_));
 sg13g2_xor2_1 _10273_ (.B(_04316_),
    .A(_03809_),
    .X(_04317_));
 sg13g2_and2_1 _10274_ (.A(_04299_),
    .B(_04317_),
    .X(_04318_));
 sg13g2_xor2_1 _10275_ (.B(_04317_),
    .A(_04299_),
    .X(_04319_));
 sg13g2_xnor2_1 _10276_ (.Y(_04320_),
    .A(_04298_),
    .B(_04319_));
 sg13g2_xor2_1 _10277_ (.B(_04320_),
    .A(_04297_),
    .X(_04321_));
 sg13g2_xnor2_1 _10278_ (.Y(_04322_),
    .A(_04206_),
    .B(_04321_));
 sg13g2_nor2b_1 _10279_ (.A(_04322_),
    .B_N(_04205_),
    .Y(_04323_));
 sg13g2_xnor2_1 _10280_ (.Y(_04324_),
    .A(_04205_),
    .B(_04322_));
 sg13g2_a21oi_1 _10281_ (.A1(_04071_),
    .A2(_04189_),
    .Y(_04325_),
    .B1(_04191_));
 sg13g2_nand2b_1 _10282_ (.Y(_04326_),
    .B(_04324_),
    .A_N(_04325_));
 sg13g2_xor2_1 _10283_ (.B(_04325_),
    .A(_04324_),
    .X(_04327_));
 sg13g2_nor2_1 _10284_ (.A(_04194_),
    .B(_04327_),
    .Y(_04328_));
 sg13g2_xor2_1 _10285_ (.B(_04327_),
    .A(_04194_),
    .X(_04329_));
 sg13g2_xnor2_1 _10286_ (.Y(_04330_),
    .A(_04204_),
    .B(_04329_));
 sg13g2_inv_1 _10287_ (.Y(_04331_),
    .A(_04330_));
 sg13g2_o21ai_1 _10288_ (.B1(net1757),
    .Y(_04332_),
    .A1(net1472),
    .A2(net621));
 sg13g2_a21oi_1 _10289_ (.A1(net1472),
    .A2(_04330_),
    .Y(_00328_),
    .B1(net622));
 sg13g2_a21oi_1 _10290_ (.A1(_04204_),
    .A2(_04329_),
    .Y(_04333_),
    .B1(_04328_));
 sg13g2_a21oi_1 _10291_ (.A1(_04298_),
    .A2(_04319_),
    .Y(_04334_),
    .B1(_04318_));
 sg13g2_o21ai_1 _10292_ (.B1(_04296_),
    .Y(_04335_),
    .A1(_04297_),
    .A2(_04320_));
 sg13g2_a21o_1 _10293_ (.A2(_04294_),
    .A1(_04256_),
    .B1(_04255_),
    .X(_04336_));
 sg13g2_o21ai_1 _10294_ (.B1(_04229_),
    .Y(_04337_),
    .A1(_04230_),
    .A2(_04253_));
 sg13g2_o21ai_1 _10295_ (.B1(_04215_),
    .Y(_04338_),
    .A1(_04216_),
    .A2(_04227_));
 sg13g2_nand2_2 _10296_ (.Y(_04339_),
    .A(_03837_),
    .B(_04213_));
 sg13g2_or3_1 _10297_ (.A(_03837_),
    .B(_03942_),
    .C(_04213_),
    .X(_04340_));
 sg13g2_nand2_2 _10298_ (.Y(_04341_),
    .A(_04339_),
    .B(_04340_));
 sg13g2_o21ai_1 _10299_ (.B1(_04223_),
    .Y(_04342_),
    .A1(_04087_),
    .A2(_04221_));
 sg13g2_a21oi_2 _10300_ (.B1(_04212_),
    .Y(_04343_),
    .A2(_03944_),
    .A1(net1616));
 sg13g2_nand2_1 _10301_ (.Y(_04344_),
    .A(net1601),
    .B(net1665));
 sg13g2_nand2_1 _10302_ (.Y(_04345_),
    .A(net1608),
    .B(net1655));
 sg13g2_nor2_1 _10303_ (.A(_05556_),
    .B(_04345_),
    .Y(_04346_));
 sg13g2_xor2_1 _10304_ (.B(_04345_),
    .A(_04220_),
    .X(_04347_));
 sg13g2_nand2b_1 _10305_ (.Y(_04348_),
    .B(_04347_),
    .A_N(_04344_));
 sg13g2_xnor2_1 _10306_ (.Y(_04349_),
    .A(_04344_),
    .B(_04347_));
 sg13g2_nor2b_1 _10307_ (.A(_04343_),
    .B_N(_04349_),
    .Y(_04350_));
 sg13g2_xnor2_1 _10308_ (.Y(_04351_),
    .A(_04343_),
    .B(_04349_));
 sg13g2_xnor2_1 _10309_ (.Y(_04352_),
    .A(_04342_),
    .B(_04351_));
 sg13g2_xor2_1 _10310_ (.B(_04352_),
    .A(_04341_),
    .X(_04353_));
 sg13g2_nand2_1 _10311_ (.Y(_04354_),
    .A(_04338_),
    .B(_04353_));
 sg13g2_xnor2_1 _10312_ (.Y(_04355_),
    .A(_04338_),
    .B(_04353_));
 sg13g2_o21ai_1 _10313_ (.B1(_04248_),
    .Y(_04356_),
    .A1(_04240_),
    .A2(_04249_));
 sg13g2_inv_1 _10314_ (.Y(_04357_),
    .A(_04356_));
 sg13g2_a21o_1 _10315_ (.A2(_04226_),
    .A1(_04217_),
    .B1(_04225_),
    .X(_04358_));
 sg13g2_nand2_1 _10316_ (.Y(_04359_),
    .A(net1568),
    .B(net1692));
 sg13g2_nand2_1 _10317_ (.Y(_04360_),
    .A(net1572),
    .B(net1679));
 sg13g2_nand2_1 _10318_ (.Y(_04361_),
    .A(net1576),
    .B(net1679));
 sg13g2_xor2_1 _10319_ (.B(_04361_),
    .A(_04235_),
    .X(_04362_));
 sg13g2_nand2b_1 _10320_ (.Y(_04363_),
    .B(_04362_),
    .A_N(_04359_));
 sg13g2_xnor2_1 _10321_ (.Y(_04364_),
    .A(_04359_),
    .B(_04362_));
 sg13g2_inv_1 _10322_ (.Y(_04365_),
    .A(_04364_));
 sg13g2_o21ai_1 _10323_ (.B1(_04246_),
    .Y(_04366_),
    .A1(_04110_),
    .A2(_04244_));
 sg13g2_nand2_1 _10324_ (.Y(_04367_),
    .A(net1579),
    .B(net1677));
 sg13g2_nand2_1 _10325_ (.Y(_04368_),
    .A(net1584),
    .B(net1666));
 sg13g2_nand2_1 _10326_ (.Y(_04369_),
    .A(net1591),
    .B(net1666));
 sg13g2_xor2_1 _10327_ (.B(_04369_),
    .A(_04243_),
    .X(_04370_));
 sg13g2_nand2b_1 _10328_ (.Y(_04371_),
    .B(_04370_),
    .A_N(_04367_));
 sg13g2_xnor2_1 _10329_ (.Y(_04372_),
    .A(_04367_),
    .B(_04370_));
 sg13g2_nand2_1 _10330_ (.Y(_04373_),
    .A(_04366_),
    .B(_04372_));
 sg13g2_xnor2_1 _10331_ (.Y(_04374_),
    .A(_04366_),
    .B(_04372_));
 sg13g2_xnor2_1 _10332_ (.Y(_04375_),
    .A(_04365_),
    .B(_04374_));
 sg13g2_nand2b_1 _10333_ (.Y(_04376_),
    .B(_04358_),
    .A_N(_04375_));
 sg13g2_xor2_1 _10334_ (.B(_04375_),
    .A(_04358_),
    .X(_04377_));
 sg13g2_xnor2_1 _10335_ (.Y(_04378_),
    .A(_04357_),
    .B(_04377_));
 sg13g2_xor2_1 _10336_ (.B(_04378_),
    .A(_04355_),
    .X(_04379_));
 sg13g2_nand2_1 _10337_ (.Y(_04380_),
    .A(_04337_),
    .B(_04379_));
 sg13g2_xnor2_1 _10338_ (.Y(_04381_),
    .A(_04337_),
    .B(_04379_));
 sg13g2_o21ai_1 _10339_ (.B1(_04272_),
    .Y(_04382_),
    .A1(_04273_),
    .A2(_04290_));
 sg13g2_o21ai_1 _10340_ (.B1(_04251_),
    .Y(_04383_),
    .A1(_04232_),
    .A2(_04252_));
 sg13g2_a21o_1 _10341_ (.A2(_04268_),
    .A1(_04262_),
    .B1(_04270_),
    .X(_04384_));
 sg13g2_o21ai_1 _10342_ (.B1(_04266_),
    .Y(_04385_),
    .A1(_04263_),
    .A2(_04267_));
 sg13g2_o21ai_1 _10343_ (.B1(_04238_),
    .Y(_04386_),
    .A1(_04102_),
    .A2(_04236_));
 sg13g2_nand2_1 _10344_ (.Y(_04387_),
    .A(net1508),
    .B(net1705));
 sg13g2_nand2_1 _10345_ (.Y(_04388_),
    .A(net1512),
    .B(net1697));
 sg13g2_nand2_1 _10346_ (.Y(_04389_),
    .A(net1564),
    .B(net1697));
 sg13g2_or2_1 _10347_ (.X(_04390_),
    .B(_04388_),
    .A(_04265_));
 sg13g2_xnor2_1 _10348_ (.Y(_04391_),
    .A(_04264_),
    .B(_04389_));
 sg13g2_xor2_1 _10349_ (.B(_04391_),
    .A(_04387_),
    .X(_04392_));
 sg13g2_xnor2_1 _10350_ (.Y(_04393_),
    .A(_04386_),
    .B(_04392_));
 sg13g2_nor2b_1 _10351_ (.A(_04393_),
    .B_N(_04385_),
    .Y(_04394_));
 sg13g2_xor2_1 _10352_ (.B(_04393_),
    .A(_04385_),
    .X(_04395_));
 sg13g2_nand2b_1 _10353_ (.Y(_04396_),
    .B(_04384_),
    .A_N(_04395_));
 sg13g2_xor2_1 _10354_ (.B(_04395_),
    .A(_04384_),
    .X(_04397_));
 sg13g2_and2_1 _10355_ (.A(net1488),
    .B(net1519),
    .X(_04398_));
 sg13g2_nand2_1 _10356_ (.Y(_04399_),
    .A(net1488),
    .B(net1519));
 sg13g2_nand2_1 _10357_ (.Y(_04400_),
    .A(net1493),
    .B(net1729));
 sg13g2_nor3_1 _10358_ (.A(_05552_),
    .B(_05570_),
    .C(_04400_),
    .Y(_04401_));
 sg13g2_a22oi_1 _10359_ (.Y(_04402_),
    .B1(net1515),
    .B2(net1490),
    .A2(net1729),
    .A1(net1493));
 sg13g2_nor2_1 _10360_ (.A(_04401_),
    .B(_04402_),
    .Y(_04403_));
 sg13g2_xnor2_1 _10361_ (.Y(_04404_),
    .A(_04399_),
    .B(_04403_));
 sg13g2_inv_1 _10362_ (.Y(_04405_),
    .A(_04404_));
 sg13g2_o21ai_1 _10363_ (.B1(_04286_),
    .Y(_04406_),
    .A1(_04150_),
    .A2(_04284_));
 sg13g2_nand2_1 _10364_ (.Y(_04407_),
    .A(net1498),
    .B(net1722));
 sg13g2_nand2_1 _10365_ (.Y(_04408_),
    .A(net1500),
    .B(net1711));
 sg13g2_nand2_1 _10366_ (.Y(_04409_),
    .A(net1504),
    .B(net1711));
 sg13g2_xor2_1 _10367_ (.B(_04409_),
    .A(_04283_),
    .X(_04410_));
 sg13g2_nand2b_1 _10368_ (.Y(_04411_),
    .B(_04410_),
    .A_N(_04407_));
 sg13g2_xnor2_1 _10369_ (.Y(_04412_),
    .A(_04407_),
    .B(_04410_));
 sg13g2_nand2_1 _10370_ (.Y(_04413_),
    .A(_04406_),
    .B(_04412_));
 sg13g2_xnor2_1 _10371_ (.Y(_04414_),
    .A(_04406_),
    .B(_04412_));
 sg13g2_xnor2_1 _10372_ (.Y(_04415_),
    .A(_04405_),
    .B(_04414_));
 sg13g2_xor2_1 _10373_ (.B(_04415_),
    .A(_04397_),
    .X(_04416_));
 sg13g2_xnor2_1 _10374_ (.Y(_04417_),
    .A(_04383_),
    .B(_04416_));
 sg13g2_nor2b_1 _10375_ (.A(_04417_),
    .B_N(_04382_),
    .Y(_04418_));
 sg13g2_xor2_1 _10376_ (.B(_04417_),
    .A(_04382_),
    .X(_04419_));
 sg13g2_xor2_1 _10377_ (.B(_04419_),
    .A(_04381_),
    .X(_04420_));
 sg13g2_nand2_1 _10378_ (.Y(_04421_),
    .A(_04336_),
    .B(_04420_));
 sg13g2_xnor2_1 _10379_ (.Y(_04422_),
    .A(_04336_),
    .B(_04420_));
 sg13g2_o21ai_1 _10380_ (.B1(_04315_),
    .Y(_04423_),
    .A1(_03809_),
    .A2(_04316_));
 sg13g2_a21o_2 _10381_ (.A2(_04291_),
    .A1(_04259_),
    .B1(_04293_),
    .X(_04424_));
 sg13g2_nand2_1 _10382_ (.Y(_04425_),
    .A(net1543),
    .B(_03807_));
 sg13g2_o21ai_1 _10383_ (.B1(_04425_),
    .Y(_04426_),
    .A1(_03807_),
    .A2(_04041_));
 sg13g2_a21o_1 _10384_ (.A2(_04311_),
    .A1(_04302_),
    .B1(_04313_),
    .X(_04427_));
 sg13g2_a21o_1 _10385_ (.A2(_04307_),
    .A1(_04304_),
    .B1(_04310_),
    .X(_04428_));
 sg13g2_o21ai_1 _10386_ (.B1(_04288_),
    .Y(_04429_),
    .A1(_04280_),
    .A2(_04289_));
 sg13g2_inv_1 _10387_ (.Y(_04430_),
    .A(_04429_));
 sg13g2_o21ai_1 _10388_ (.B1(_04305_),
    .Y(_04431_),
    .A1(_03900_),
    .A2(_04306_));
 sg13g2_a21o_1 _10389_ (.A2(_04278_),
    .A1(_04274_),
    .B1(_04276_),
    .X(_04432_));
 sg13g2_nand2_1 _10390_ (.Y(_04433_),
    .A(net1527),
    .B(_04140_));
 sg13g2_o21ai_1 _10391_ (.B1(_04433_),
    .Y(_04434_),
    .A1(_04140_),
    .A2(_04274_));
 sg13g2_xnor2_1 _10392_ (.Y(_04435_),
    .A(_04009_),
    .B(_04434_));
 sg13g2_xnor2_1 _10393_ (.Y(_04436_),
    .A(_04432_),
    .B(_04435_));
 sg13g2_nor2b_1 _10394_ (.A(_04436_),
    .B_N(_04431_),
    .Y(_04437_));
 sg13g2_xor2_1 _10395_ (.B(_04436_),
    .A(_04431_),
    .X(_04438_));
 sg13g2_xor2_1 _10396_ (.B(_04438_),
    .A(_04429_),
    .X(_04439_));
 sg13g2_nand2b_1 _10397_ (.Y(_04440_),
    .B(_04428_),
    .A_N(_04439_));
 sg13g2_xnor2_1 _10398_ (.Y(_04441_),
    .A(_04428_),
    .B(_04439_));
 sg13g2_nand2_1 _10399_ (.Y(_04442_),
    .A(_04427_),
    .B(_04441_));
 sg13g2_xnor2_1 _10400_ (.Y(_04443_),
    .A(_04427_),
    .B(_04441_));
 sg13g2_xor2_1 _10401_ (.B(_04443_),
    .A(_04426_),
    .X(_04444_));
 sg13g2_xnor2_1 _10402_ (.Y(_04445_),
    .A(_04424_),
    .B(_04444_));
 sg13g2_nor2b_1 _10403_ (.A(_04445_),
    .B_N(_04423_),
    .Y(_04446_));
 sg13g2_xor2_1 _10404_ (.B(_04445_),
    .A(_04423_),
    .X(_04447_));
 sg13g2_xor2_1 _10405_ (.B(_04447_),
    .A(_04422_),
    .X(_04448_));
 sg13g2_nand2_1 _10406_ (.Y(_04449_),
    .A(_04335_),
    .B(_04448_));
 sg13g2_xnor2_1 _10407_ (.Y(_04450_),
    .A(_04335_),
    .B(_04448_));
 sg13g2_xor2_1 _10408_ (.B(_04450_),
    .A(_04334_),
    .X(_04451_));
 sg13g2_a21o_1 _10409_ (.A2(_04321_),
    .A1(_04206_),
    .B1(_04323_),
    .X(_04452_));
 sg13g2_nand2_1 _10410_ (.Y(_04453_),
    .A(_04451_),
    .B(_04452_));
 sg13g2_xor2_1 _10411_ (.B(_04452_),
    .A(_04451_),
    .X(_04454_));
 sg13g2_nor2b_1 _10412_ (.A(_04326_),
    .B_N(_04454_),
    .Y(_04455_));
 sg13g2_xnor2_1 _10413_ (.Y(_04456_),
    .A(_04326_),
    .B(_04454_));
 sg13g2_xnor2_1 _10414_ (.Y(_04457_),
    .A(_04333_),
    .B(_04456_));
 sg13g2_o21ai_1 _10415_ (.B1(net1757),
    .Y(_04458_),
    .A1(net1400),
    .A2(_04457_));
 sg13g2_a21oi_1 _10416_ (.A1(net1400),
    .A2(_05544_),
    .Y(_00329_),
    .B1(_04458_));
 sg13g2_and2_1 _10417_ (.A(_04329_),
    .B(_04456_),
    .X(_04459_));
 sg13g2_a21o_1 _10418_ (.A2(_04456_),
    .A1(_04328_),
    .B1(_04455_),
    .X(_04460_));
 sg13g2_a21o_1 _10419_ (.A2(_04459_),
    .A1(_04204_),
    .B1(_04460_),
    .X(_04461_));
 sg13g2_a21o_1 _10420_ (.A2(_04444_),
    .A1(_04424_),
    .B1(_04446_),
    .X(_04462_));
 sg13g2_o21ai_1 _10421_ (.B1(_04421_),
    .Y(_04463_),
    .A1(_04422_),
    .A2(_04447_));
 sg13g2_o21ai_1 _10422_ (.B1(_04380_),
    .Y(_04464_),
    .A1(_04381_),
    .A2(_04419_));
 sg13g2_o21ai_1 _10423_ (.B1(_04354_),
    .Y(_04465_),
    .A1(_04355_),
    .A2(_04378_));
 sg13g2_o21ai_1 _10424_ (.B1(_04339_),
    .Y(_04466_),
    .A1(_04341_),
    .A2(_04352_));
 sg13g2_o21ai_1 _10425_ (.B1(_04348_),
    .Y(_04467_),
    .A1(_04220_),
    .A2(_04345_));
 sg13g2_o21ai_1 _10426_ (.B1(net1655),
    .Y(_04468_),
    .A1(net1606),
    .A2(net1608));
 sg13g2_or2_1 _10427_ (.X(_04469_),
    .B(_04468_),
    .A(_04346_));
 sg13g2_nand2_1 _10428_ (.Y(_04470_),
    .A(net1601),
    .B(net1659));
 sg13g2_nor2_1 _10429_ (.A(_04469_),
    .B(_04470_),
    .Y(_04471_));
 sg13g2_xor2_1 _10430_ (.B(_04470_),
    .A(_04469_),
    .X(_04472_));
 sg13g2_nor2b_1 _10431_ (.A(_04343_),
    .B_N(_04472_),
    .Y(_04473_));
 sg13g2_xnor2_1 _10432_ (.Y(_04474_),
    .A(_04343_),
    .B(_04472_));
 sg13g2_xnor2_1 _10433_ (.Y(_04475_),
    .A(_04467_),
    .B(_04474_));
 sg13g2_xor2_1 _10434_ (.B(_04475_),
    .A(_04341_),
    .X(_04476_));
 sg13g2_nand2_1 _10435_ (.Y(_04477_),
    .A(_04466_),
    .B(_04476_));
 sg13g2_xnor2_1 _10436_ (.Y(_04478_),
    .A(_04466_),
    .B(_04476_));
 sg13g2_o21ai_1 _10437_ (.B1(_04373_),
    .Y(_04479_),
    .A1(_04365_),
    .A2(_04374_));
 sg13g2_inv_1 _10438_ (.Y(_04480_),
    .A(_04479_));
 sg13g2_a21o_1 _10439_ (.A2(_04351_),
    .A1(_04342_),
    .B1(_04350_),
    .X(_04481_));
 sg13g2_nand2_1 _10440_ (.Y(_04482_),
    .A(net1568),
    .B(net1684));
 sg13g2_nand2_1 _10441_ (.Y(_04483_),
    .A(net1572),
    .B(net1674));
 sg13g2_nand2_1 _10442_ (.Y(_04484_),
    .A(net1576),
    .B(net1677));
 sg13g2_xor2_1 _10443_ (.B(_04484_),
    .A(_04360_),
    .X(_04485_));
 sg13g2_nand2b_1 _10444_ (.Y(_04486_),
    .B(_04485_),
    .A_N(_04482_));
 sg13g2_xnor2_1 _10445_ (.Y(_04487_),
    .A(_04482_),
    .B(_04485_));
 sg13g2_inv_1 _10446_ (.Y(_04488_),
    .A(_04487_));
 sg13g2_o21ai_1 _10447_ (.B1(_04371_),
    .Y(_04489_),
    .A1(_04243_),
    .A2(_04369_));
 sg13g2_nand2_1 _10448_ (.Y(_04490_),
    .A(net1579),
    .B(net1673));
 sg13g2_nand2_1 _10449_ (.Y(_04491_),
    .A(net1584),
    .B(net1662));
 sg13g2_nand2_1 _10450_ (.Y(_04492_),
    .A(net1591),
    .B(net1665));
 sg13g2_xor2_1 _10451_ (.B(_04492_),
    .A(_04368_),
    .X(_04493_));
 sg13g2_nand2b_1 _10452_ (.Y(_04494_),
    .B(_04493_),
    .A_N(_04490_));
 sg13g2_xnor2_1 _10453_ (.Y(_04495_),
    .A(_04490_),
    .B(_04493_));
 sg13g2_nand2_1 _10454_ (.Y(_04496_),
    .A(_04489_),
    .B(_04495_));
 sg13g2_xnor2_1 _10455_ (.Y(_04497_),
    .A(_04489_),
    .B(_04495_));
 sg13g2_xnor2_1 _10456_ (.Y(_04498_),
    .A(_04488_),
    .B(_04497_));
 sg13g2_nand2b_1 _10457_ (.Y(_04499_),
    .B(_04481_),
    .A_N(_04498_));
 sg13g2_xor2_1 _10458_ (.B(_04498_),
    .A(_04481_),
    .X(_04500_));
 sg13g2_xnor2_1 _10459_ (.Y(_04501_),
    .A(_04480_),
    .B(_04500_));
 sg13g2_xor2_1 _10460_ (.B(_04501_),
    .A(_04478_),
    .X(_04502_));
 sg13g2_nand2_1 _10461_ (.Y(_04503_),
    .A(_04465_),
    .B(_04502_));
 sg13g2_xnor2_1 _10462_ (.Y(_04504_),
    .A(_04465_),
    .B(_04502_));
 sg13g2_o21ai_1 _10463_ (.B1(_04396_),
    .Y(_04505_),
    .A1(_04397_),
    .A2(_04415_));
 sg13g2_o21ai_1 _10464_ (.B1(_04376_),
    .Y(_04506_),
    .A1(_04357_),
    .A2(_04377_));
 sg13g2_a21o_1 _10465_ (.A2(_04392_),
    .A1(_04386_),
    .B1(_04394_),
    .X(_04507_));
 sg13g2_o21ai_1 _10466_ (.B1(_04390_),
    .Y(_04508_),
    .A1(_04387_),
    .A2(_04391_));
 sg13g2_o21ai_1 _10467_ (.B1(_04363_),
    .Y(_04509_),
    .A1(_04235_),
    .A2(_04361_));
 sg13g2_nand2_1 _10468_ (.Y(_04510_),
    .A(net1508),
    .B(net1702));
 sg13g2_nand2_1 _10469_ (.Y(_04511_),
    .A(net1512),
    .B(net1692));
 sg13g2_nand2_1 _10470_ (.Y(_04512_),
    .A(net1564),
    .B(net1692));
 sg13g2_or2_1 _10471_ (.X(_04513_),
    .B(_04511_),
    .A(_04389_));
 sg13g2_xnor2_1 _10472_ (.Y(_04514_),
    .A(_04388_),
    .B(_04512_));
 sg13g2_xor2_1 _10473_ (.B(_04514_),
    .A(_04510_),
    .X(_04515_));
 sg13g2_xnor2_1 _10474_ (.Y(_04516_),
    .A(_04509_),
    .B(_04515_));
 sg13g2_nor2b_1 _10475_ (.A(_04516_),
    .B_N(_04508_),
    .Y(_04517_));
 sg13g2_xor2_1 _10476_ (.B(_04516_),
    .A(_04508_),
    .X(_04518_));
 sg13g2_nand2b_1 _10477_ (.Y(_04519_),
    .B(_04507_),
    .A_N(_04518_));
 sg13g2_xor2_1 _10478_ (.B(_04518_),
    .A(_04507_),
    .X(_04520_));
 sg13g2_and2_1 _10479_ (.A(net1485),
    .B(net1515),
    .X(_04521_));
 sg13g2_nand2_1 _10480_ (.Y(_04522_),
    .A(net1485),
    .B(net1515));
 sg13g2_nor3_1 _10481_ (.A(_05552_),
    .B(_05569_),
    .C(_04400_),
    .Y(_04523_));
 sg13g2_a22oi_1 _10482_ (.Y(_04524_),
    .B1(net1729),
    .B2(net1490),
    .A2(net1722),
    .A1(net1493));
 sg13g2_nor2_1 _10483_ (.A(_04523_),
    .B(_04524_),
    .Y(_04525_));
 sg13g2_xnor2_1 _10484_ (.Y(_04526_),
    .A(_04522_),
    .B(_04525_));
 sg13g2_inv_1 _10485_ (.Y(_04527_),
    .A(_04526_));
 sg13g2_o21ai_1 _10486_ (.B1(_04411_),
    .Y(_04528_),
    .A1(_04283_),
    .A2(_04409_));
 sg13g2_nand2_1 _10487_ (.Y(_04529_),
    .A(net1498),
    .B(net1716));
 sg13g2_nand2_1 _10488_ (.Y(_04530_),
    .A(net1500),
    .B(net1705));
 sg13g2_nand2_1 _10489_ (.Y(_04531_),
    .A(net1503),
    .B(net1705));
 sg13g2_xor2_1 _10490_ (.B(_04531_),
    .A(_04408_),
    .X(_04532_));
 sg13g2_nand2b_1 _10491_ (.Y(_04533_),
    .B(_04532_),
    .A_N(_04529_));
 sg13g2_xnor2_1 _10492_ (.Y(_04534_),
    .A(_04529_),
    .B(_04532_));
 sg13g2_nand2_1 _10493_ (.Y(_04535_),
    .A(_04528_),
    .B(_04534_));
 sg13g2_xnor2_1 _10494_ (.Y(_04536_),
    .A(_04528_),
    .B(_04534_));
 sg13g2_xnor2_1 _10495_ (.Y(_04537_),
    .A(_04527_),
    .B(_04536_));
 sg13g2_xor2_1 _10496_ (.B(_04537_),
    .A(_04520_),
    .X(_04538_));
 sg13g2_xnor2_1 _10497_ (.Y(_04539_),
    .A(_04506_),
    .B(_04538_));
 sg13g2_nor2b_1 _10498_ (.A(_04539_),
    .B_N(_04505_),
    .Y(_04540_));
 sg13g2_xor2_1 _10499_ (.B(_04539_),
    .A(_04505_),
    .X(_04541_));
 sg13g2_xor2_1 _10500_ (.B(_04541_),
    .A(_04504_),
    .X(_04542_));
 sg13g2_nand2_1 _10501_ (.Y(_04543_),
    .A(_04464_),
    .B(_04542_));
 sg13g2_xnor2_1 _10502_ (.Y(_04544_),
    .A(_04464_),
    .B(_04542_));
 sg13g2_o21ai_1 _10503_ (.B1(_04442_),
    .Y(_04545_),
    .A1(_04426_),
    .A2(_04443_));
 sg13g2_a21o_2 _10504_ (.A2(_04416_),
    .A1(_04383_),
    .B1(_04418_),
    .X(_04546_));
 sg13g2_o21ai_1 _10505_ (.B1(_04440_),
    .Y(_04547_),
    .A1(_04430_),
    .A2(_04438_));
 sg13g2_a21o_1 _10506_ (.A2(_04435_),
    .A1(_04432_),
    .B1(_04437_),
    .X(_04548_));
 sg13g2_o21ai_1 _10507_ (.B1(_04413_),
    .Y(_04549_),
    .A1(_04405_),
    .A2(_04414_));
 sg13g2_inv_1 _10508_ (.Y(_04550_),
    .A(_04549_));
 sg13g2_o21ai_1 _10509_ (.B1(_04433_),
    .Y(_04551_),
    .A1(_04010_),
    .A2(_04434_));
 sg13g2_a21o_1 _10510_ (.A2(_04403_),
    .A1(_04398_),
    .B1(_04401_),
    .X(_04552_));
 sg13g2_nand2_1 _10511_ (.Y(_04553_),
    .A(net1519),
    .B(_04274_));
 sg13g2_o21ai_1 _10512_ (.B1(_04553_),
    .Y(_04554_),
    .A1(_04274_),
    .A2(_04398_));
 sg13g2_xnor2_1 _10513_ (.Y(_04555_),
    .A(_04140_),
    .B(_04554_));
 sg13g2_xnor2_1 _10514_ (.Y(_04556_),
    .A(_04552_),
    .B(_04555_));
 sg13g2_nor2b_1 _10515_ (.A(_04556_),
    .B_N(_04551_),
    .Y(_04557_));
 sg13g2_xor2_1 _10516_ (.B(_04556_),
    .A(_04551_),
    .X(_04558_));
 sg13g2_xor2_1 _10517_ (.B(_04558_),
    .A(_04549_),
    .X(_04559_));
 sg13g2_nand2b_1 _10518_ (.Y(_04560_),
    .B(_04548_),
    .A_N(_04559_));
 sg13g2_xor2_1 _10519_ (.B(_04559_),
    .A(_04548_),
    .X(_04561_));
 sg13g2_nor2b_1 _10520_ (.A(_04561_),
    .B_N(_04547_),
    .Y(_04562_));
 sg13g2_xor2_1 _10521_ (.B(_04561_),
    .A(_04547_),
    .X(_04563_));
 sg13g2_inv_1 _10522_ (.Y(_04564_),
    .A(_04563_));
 sg13g2_nor2_1 _10523_ (.A(_04169_),
    .B(_04174_),
    .Y(_04565_));
 sg13g2_xnor2_1 _10524_ (.Y(_04566_),
    .A(_04169_),
    .B(_04174_));
 sg13g2_xnor2_1 _10525_ (.Y(_04567_),
    .A(_04039_),
    .B(_04566_));
 sg13g2_xnor2_1 _10526_ (.Y(_04568_),
    .A(_04563_),
    .B(_04567_));
 sg13g2_and2_1 _10527_ (.A(_04546_),
    .B(_04568_),
    .X(_04569_));
 sg13g2_xor2_1 _10528_ (.B(_04568_),
    .A(_04546_),
    .X(_04570_));
 sg13g2_xnor2_1 _10529_ (.Y(_04571_),
    .A(_04545_),
    .B(_04570_));
 sg13g2_xor2_1 _10530_ (.B(_04571_),
    .A(_04544_),
    .X(_04572_));
 sg13g2_xnor2_1 _10531_ (.Y(_04573_),
    .A(_04463_),
    .B(_04572_));
 sg13g2_nor2b_1 _10532_ (.A(_04573_),
    .B_N(_04462_),
    .Y(_04574_));
 sg13g2_xor2_1 _10533_ (.B(_04573_),
    .A(_04462_),
    .X(_04575_));
 sg13g2_o21ai_1 _10534_ (.B1(_04449_),
    .Y(_04576_),
    .A1(_04334_),
    .A2(_04450_));
 sg13g2_nand2b_1 _10535_ (.Y(_04577_),
    .B(_04576_),
    .A_N(_04575_));
 sg13g2_xor2_1 _10536_ (.B(_04576_),
    .A(_04575_),
    .X(_04578_));
 sg13g2_nor2_1 _10537_ (.A(_04453_),
    .B(_04578_),
    .Y(_04579_));
 sg13g2_xor2_1 _10538_ (.B(_04578_),
    .A(_04453_),
    .X(_04580_));
 sg13g2_xnor2_1 _10539_ (.Y(_04581_),
    .A(_04461_),
    .B(_04580_));
 sg13g2_o21ai_1 _10540_ (.B1(net1759),
    .Y(_04582_),
    .A1(net1472),
    .A2(net628));
 sg13g2_a21oi_1 _10541_ (.A1(net1472),
    .A2(_04581_),
    .Y(_00330_),
    .B1(net629));
 sg13g2_a21oi_1 _10542_ (.A1(_04461_),
    .A2(_04580_),
    .Y(_04583_),
    .B1(_04579_));
 sg13g2_nand3_1 _10543_ (.B(_03807_),
    .C(_04174_),
    .A(net1543),
    .Y(_04584_));
 sg13g2_a21oi_1 _10544_ (.A1(_04545_),
    .A2(_04570_),
    .Y(_04585_),
    .B1(_04569_));
 sg13g2_nor2_1 _10545_ (.A(_04584_),
    .B(_04585_),
    .Y(_04586_));
 sg13g2_xnor2_1 _10546_ (.Y(_04587_),
    .A(_04584_),
    .B(_04585_));
 sg13g2_o21ai_1 _10547_ (.B1(_04543_),
    .Y(_04588_),
    .A1(_04544_),
    .A2(_04571_));
 sg13g2_o21ai_1 _10548_ (.B1(_04503_),
    .Y(_04589_),
    .A1(_04504_),
    .A2(_04541_));
 sg13g2_o21ai_1 _10549_ (.B1(_04477_),
    .Y(_04590_),
    .A1(_04478_),
    .A2(_04501_));
 sg13g2_o21ai_1 _10550_ (.B1(_04339_),
    .Y(_04591_),
    .A1(_04341_),
    .A2(_04475_));
 sg13g2_nor2_1 _10551_ (.A(_04346_),
    .B(_04471_),
    .Y(_04592_));
 sg13g2_nand2_1 _10552_ (.Y(_04593_),
    .A(net1601),
    .B(net1655));
 sg13g2_nor2_1 _10553_ (.A(_04469_),
    .B(_04593_),
    .Y(_04594_));
 sg13g2_xor2_1 _10554_ (.B(_04593_),
    .A(_04469_),
    .X(_04595_));
 sg13g2_nand2b_1 _10555_ (.Y(_04596_),
    .B(_04595_),
    .A_N(_04343_));
 sg13g2_xnor2_1 _10556_ (.Y(_04597_),
    .A(_04343_),
    .B(_04595_));
 sg13g2_inv_1 _10557_ (.Y(_04598_),
    .A(_04597_));
 sg13g2_xnor2_1 _10558_ (.Y(_04599_),
    .A(_04592_),
    .B(_04597_));
 sg13g2_inv_1 _10559_ (.Y(_04600_),
    .A(_04599_));
 sg13g2_xnor2_1 _10560_ (.Y(_04601_),
    .A(_04341_),
    .B(_04599_));
 sg13g2_nand2_1 _10561_ (.Y(_04602_),
    .A(_04591_),
    .B(_04601_));
 sg13g2_xnor2_1 _10562_ (.Y(_04603_),
    .A(_04591_),
    .B(_04601_));
 sg13g2_o21ai_1 _10563_ (.B1(_04496_),
    .Y(_04604_),
    .A1(_04488_),
    .A2(_04497_));
 sg13g2_a21o_1 _10564_ (.A2(_04474_),
    .A1(_04467_),
    .B1(_04473_),
    .X(_04605_));
 sg13g2_inv_1 _10565_ (.Y(_04606_),
    .A(_04605_));
 sg13g2_nand2_1 _10566_ (.Y(_04607_),
    .A(net1568),
    .B(net1683));
 sg13g2_nand2_1 _10567_ (.Y(_04608_),
    .A(net1572),
    .B(net1670));
 sg13g2_nand2_1 _10568_ (.Y(_04609_),
    .A(net1576),
    .B(net1670));
 sg13g2_xor2_1 _10569_ (.B(_04609_),
    .A(_04483_),
    .X(_04610_));
 sg13g2_nand2b_1 _10570_ (.Y(_04611_),
    .B(_04610_),
    .A_N(_04607_));
 sg13g2_xnor2_1 _10571_ (.Y(_04612_),
    .A(_04607_),
    .B(_04610_));
 sg13g2_inv_1 _10572_ (.Y(_04613_),
    .A(_04612_));
 sg13g2_o21ai_1 _10573_ (.B1(_04494_),
    .Y(_04614_),
    .A1(_04368_),
    .A2(_04492_));
 sg13g2_nand2_1 _10574_ (.Y(_04615_),
    .A(net1579),
    .B(net1667));
 sg13g2_nand2_1 _10575_ (.Y(_04616_),
    .A(net1584),
    .B(net1659));
 sg13g2_nand2_1 _10576_ (.Y(_04617_),
    .A(net1591),
    .B(net1659));
 sg13g2_xor2_1 _10577_ (.B(_04617_),
    .A(_04491_),
    .X(_04618_));
 sg13g2_nand2b_1 _10578_ (.Y(_04619_),
    .B(_04618_),
    .A_N(_04615_));
 sg13g2_xnor2_1 _10579_ (.Y(_04620_),
    .A(_04615_),
    .B(_04618_));
 sg13g2_nand2_1 _10580_ (.Y(_04621_),
    .A(_04614_),
    .B(_04620_));
 sg13g2_xnor2_1 _10581_ (.Y(_04622_),
    .A(_04614_),
    .B(_04620_));
 sg13g2_xnor2_1 _10582_ (.Y(_04623_),
    .A(_04613_),
    .B(_04622_));
 sg13g2_xor2_1 _10583_ (.B(_04623_),
    .A(_04605_),
    .X(_04624_));
 sg13g2_nand2b_1 _10584_ (.Y(_04625_),
    .B(_04604_),
    .A_N(_04624_));
 sg13g2_xor2_1 _10585_ (.B(_04624_),
    .A(_04604_),
    .X(_04626_));
 sg13g2_xor2_1 _10586_ (.B(_04626_),
    .A(_04603_),
    .X(_04627_));
 sg13g2_nand2_1 _10587_ (.Y(_04628_),
    .A(_04590_),
    .B(_04627_));
 sg13g2_xnor2_1 _10588_ (.Y(_04629_),
    .A(_04590_),
    .B(_04627_));
 sg13g2_o21ai_1 _10589_ (.B1(_04519_),
    .Y(_04630_),
    .A1(_04520_),
    .A2(_04537_));
 sg13g2_o21ai_1 _10590_ (.B1(_04499_),
    .Y(_04631_),
    .A1(_04480_),
    .A2(_04500_));
 sg13g2_a21o_1 _10591_ (.A2(_04515_),
    .A1(_04509_),
    .B1(_04517_),
    .X(_04632_));
 sg13g2_o21ai_1 _10592_ (.B1(_04513_),
    .Y(_04633_),
    .A1(_04510_),
    .A2(_04514_));
 sg13g2_o21ai_1 _10593_ (.B1(_04486_),
    .Y(_04634_),
    .A1(_04360_),
    .A2(_04484_));
 sg13g2_nand2_1 _10594_ (.Y(_04635_),
    .A(net1507),
    .B(net1697));
 sg13g2_nand2_1 _10595_ (.Y(_04636_),
    .A(net1512),
    .B(net1685));
 sg13g2_nand2_1 _10596_ (.Y(_04637_),
    .A(net1564),
    .B(net1684));
 sg13g2_or2_1 _10597_ (.X(_04638_),
    .B(_04636_),
    .A(_04512_));
 sg13g2_xnor2_1 _10598_ (.Y(_04639_),
    .A(_04511_),
    .B(_04637_));
 sg13g2_xor2_1 _10599_ (.B(_04639_),
    .A(_04635_),
    .X(_04640_));
 sg13g2_xnor2_1 _10600_ (.Y(_04641_),
    .A(_04634_),
    .B(_04640_));
 sg13g2_nor2b_1 _10601_ (.A(_04641_),
    .B_N(_04633_),
    .Y(_04642_));
 sg13g2_xor2_1 _10602_ (.B(_04641_),
    .A(_04633_),
    .X(_04643_));
 sg13g2_nand2b_1 _10603_ (.Y(_04644_),
    .B(_04632_),
    .A_N(_04643_));
 sg13g2_xor2_1 _10604_ (.B(_04643_),
    .A(_04632_),
    .X(_04645_));
 sg13g2_and2_1 _10605_ (.A(net1485),
    .B(net1729),
    .X(_04646_));
 sg13g2_nand2_1 _10606_ (.Y(_04647_),
    .A(net1485),
    .B(net1729));
 sg13g2_nand2_1 _10607_ (.Y(_04648_),
    .A(net1492),
    .B(net1716));
 sg13g2_nor3_1 _10608_ (.A(_05553_),
    .B(_05569_),
    .C(_04648_),
    .Y(_04649_));
 sg13g2_a22oi_1 _10609_ (.Y(_04650_),
    .B1(net1722),
    .B2(net1492),
    .A2(net1716),
    .A1(net1496));
 sg13g2_nor2_1 _10610_ (.A(_04649_),
    .B(_04650_),
    .Y(_04651_));
 sg13g2_xnor2_1 _10611_ (.Y(_04652_),
    .A(_04647_),
    .B(_04651_));
 sg13g2_inv_1 _10612_ (.Y(_04653_),
    .A(_04652_));
 sg13g2_o21ai_1 _10613_ (.B1(_04533_),
    .Y(_04654_),
    .A1(_04408_),
    .A2(_04531_));
 sg13g2_nand2_1 _10614_ (.Y(_04655_),
    .A(net1497),
    .B(net1711));
 sg13g2_nand2_1 _10615_ (.Y(_04656_),
    .A(net1500),
    .B(net1702));
 sg13g2_nand2_1 _10616_ (.Y(_04657_),
    .A(net1503),
    .B(net1702));
 sg13g2_xor2_1 _10617_ (.B(_04657_),
    .A(_04530_),
    .X(_04658_));
 sg13g2_nand2b_1 _10618_ (.Y(_04659_),
    .B(_04658_),
    .A_N(_04655_));
 sg13g2_xnor2_1 _10619_ (.Y(_04660_),
    .A(_04655_),
    .B(_04658_));
 sg13g2_nand2_1 _10620_ (.Y(_04661_),
    .A(_04654_),
    .B(_04660_));
 sg13g2_xnor2_1 _10621_ (.Y(_04662_),
    .A(_04654_),
    .B(_04660_));
 sg13g2_xnor2_1 _10622_ (.Y(_04663_),
    .A(_04653_),
    .B(_04662_));
 sg13g2_xor2_1 _10623_ (.B(_04663_),
    .A(_04645_),
    .X(_04664_));
 sg13g2_xnor2_1 _10624_ (.Y(_04665_),
    .A(_04631_),
    .B(_04664_));
 sg13g2_nor2b_1 _10625_ (.A(_04665_),
    .B_N(_04630_),
    .Y(_04666_));
 sg13g2_xor2_1 _10626_ (.B(_04665_),
    .A(_04630_),
    .X(_04667_));
 sg13g2_xor2_1 _10627_ (.B(_04667_),
    .A(_04629_),
    .X(_04668_));
 sg13g2_nand2_1 _10628_ (.Y(_04669_),
    .A(_04589_),
    .B(_04668_));
 sg13g2_xnor2_1 _10629_ (.Y(_04670_),
    .A(_04589_),
    .B(_04668_));
 sg13g2_a21oi_1 _10630_ (.A1(_04564_),
    .A2(_04567_),
    .Y(_04671_),
    .B1(_04562_));
 sg13g2_a21o_2 _10631_ (.A2(_04538_),
    .A1(_04506_),
    .B1(_04540_),
    .X(_04672_));
 sg13g2_o21ai_1 _10632_ (.B1(_04560_),
    .Y(_04673_),
    .A1(_04550_),
    .A2(_04558_));
 sg13g2_a21o_1 _10633_ (.A2(_04555_),
    .A1(_04552_),
    .B1(_04557_),
    .X(_04674_));
 sg13g2_o21ai_1 _10634_ (.B1(_04535_),
    .Y(_04675_),
    .A1(_04527_),
    .A2(_04536_));
 sg13g2_inv_1 _10635_ (.Y(_04676_),
    .A(_04675_));
 sg13g2_o21ai_1 _10636_ (.B1(_04553_),
    .Y(_04677_),
    .A1(_04141_),
    .A2(_04554_));
 sg13g2_a21o_1 _10637_ (.A2(_04525_),
    .A1(_04521_),
    .B1(_04523_),
    .X(_04678_));
 sg13g2_nand2_1 _10638_ (.Y(_04679_),
    .A(net1515),
    .B(_04398_));
 sg13g2_o21ai_1 _10639_ (.B1(_04679_),
    .Y(_04680_),
    .A1(_04398_),
    .A2(_04521_));
 sg13g2_xnor2_1 _10640_ (.Y(_04681_),
    .A(_04274_),
    .B(_04680_));
 sg13g2_xnor2_1 _10641_ (.Y(_04682_),
    .A(_04678_),
    .B(_04681_));
 sg13g2_nor2b_1 _10642_ (.A(_04682_),
    .B_N(_04677_),
    .Y(_04683_));
 sg13g2_xor2_1 _10643_ (.B(_04682_),
    .A(_04677_),
    .X(_04684_));
 sg13g2_xor2_1 _10644_ (.B(_04684_),
    .A(_04675_),
    .X(_04685_));
 sg13g2_nand2b_1 _10645_ (.Y(_04686_),
    .B(_04674_),
    .A_N(_04685_));
 sg13g2_xor2_1 _10646_ (.B(_04685_),
    .A(_04674_),
    .X(_04687_));
 sg13g2_nand2b_1 _10647_ (.Y(_04688_),
    .B(_04673_),
    .A_N(_04687_));
 sg13g2_xor2_1 _10648_ (.B(_04687_),
    .A(_04673_),
    .X(_04689_));
 sg13g2_nand2_1 _10649_ (.Y(_04690_),
    .A(_04303_),
    .B(_04307_));
 sg13g2_xnor2_1 _10650_ (.Y(_04691_),
    .A(_04303_),
    .B(_04307_));
 sg13g2_xor2_1 _10651_ (.B(_04691_),
    .A(_03809_),
    .X(_04692_));
 sg13g2_a21oi_1 _10652_ (.A1(_04038_),
    .A2(_04174_),
    .Y(_04693_),
    .B1(_03566_));
 sg13g2_nor2_1 _10653_ (.A(_04565_),
    .B(_04693_),
    .Y(_04694_));
 sg13g2_nand2_1 _10654_ (.Y(_04695_),
    .A(_04692_),
    .B(_04694_));
 sg13g2_xnor2_1 _10655_ (.Y(_04696_),
    .A(_04692_),
    .B(_04694_));
 sg13g2_xor2_1 _10656_ (.B(_04696_),
    .A(_04689_),
    .X(_04697_));
 sg13g2_nand2_1 _10657_ (.Y(_04698_),
    .A(_04672_),
    .B(_04697_));
 sg13g2_xnor2_1 _10658_ (.Y(_04699_),
    .A(_04672_),
    .B(_04697_));
 sg13g2_xnor2_1 _10659_ (.Y(_04700_),
    .A(_04671_),
    .B(_04699_));
 sg13g2_xor2_1 _10660_ (.B(_04700_),
    .A(_04670_),
    .X(_04701_));
 sg13g2_xnor2_1 _10661_ (.Y(_04702_),
    .A(_04588_),
    .B(_04701_));
 sg13g2_nor2_1 _10662_ (.A(_04587_),
    .B(_04702_),
    .Y(_04703_));
 sg13g2_xor2_1 _10663_ (.B(_04702_),
    .A(_04587_),
    .X(_04704_));
 sg13g2_a21oi_1 _10664_ (.A1(_04463_),
    .A2(_04572_),
    .Y(_04705_),
    .B1(_04574_));
 sg13g2_nor2b_1 _10665_ (.A(_04705_),
    .B_N(_04704_),
    .Y(_04706_));
 sg13g2_xnor2_1 _10666_ (.Y(_04707_),
    .A(_04704_),
    .B(_04705_));
 sg13g2_nand2b_1 _10667_ (.Y(_04708_),
    .B(_04707_),
    .A_N(_04577_));
 sg13g2_xnor2_1 _10668_ (.Y(_04709_),
    .A(_04577_),
    .B(_04707_));
 sg13g2_inv_1 _10669_ (.Y(_04710_),
    .A(_04709_));
 sg13g2_xnor2_1 _10670_ (.Y(_04711_),
    .A(_04583_),
    .B(_04709_));
 sg13g2_o21ai_1 _10671_ (.B1(net1757),
    .Y(_04712_),
    .A1(net1400),
    .A2(_04711_));
 sg13g2_a21oi_1 _10672_ (.A1(net1400),
    .A2(_05543_),
    .Y(_00331_),
    .B1(_04712_));
 sg13g2_a21oi_1 _10673_ (.A1(_04588_),
    .A2(_04701_),
    .Y(_04713_),
    .B1(_04703_));
 sg13g2_o21ai_1 _10674_ (.B1(_04698_),
    .Y(_04714_),
    .A1(_04671_),
    .A2(_04699_));
 sg13g2_nor2b_1 _10675_ (.A(_04695_),
    .B_N(_04714_),
    .Y(_04715_));
 sg13g2_xor2_1 _10676_ (.B(_04714_),
    .A(_04695_),
    .X(_04716_));
 sg13g2_o21ai_1 _10677_ (.B1(_04669_),
    .Y(_04717_),
    .A1(_04670_),
    .A2(_04700_));
 sg13g2_o21ai_1 _10678_ (.B1(_04628_),
    .Y(_04718_),
    .A1(_04629_),
    .A2(_04667_));
 sg13g2_o21ai_1 _10679_ (.B1(_04602_),
    .Y(_04719_),
    .A1(_04603_),
    .A2(_04626_));
 sg13g2_o21ai_1 _10680_ (.B1(_04339_),
    .Y(_04720_),
    .A1(_04341_),
    .A2(_04600_));
 sg13g2_nor2_1 _10681_ (.A(_04346_),
    .B(_04594_),
    .Y(_04721_));
 sg13g2_xnor2_1 _10682_ (.Y(_04722_),
    .A(_04597_),
    .B(_04721_));
 sg13g2_xnor2_1 _10683_ (.Y(_04723_),
    .A(_04341_),
    .B(_04722_));
 sg13g2_nand2_1 _10684_ (.Y(_04724_),
    .A(_04720_),
    .B(_04723_));
 sg13g2_xnor2_1 _10685_ (.Y(_04725_),
    .A(_04720_),
    .B(_04723_));
 sg13g2_o21ai_1 _10686_ (.B1(_04621_),
    .Y(_04726_),
    .A1(_04613_),
    .A2(_04622_));
 sg13g2_o21ai_1 _10687_ (.B1(_04596_),
    .Y(_04727_),
    .A1(_04592_),
    .A2(_04598_));
 sg13g2_nand2_1 _10688_ (.Y(_04728_),
    .A(net1568),
    .B(net1674));
 sg13g2_nand2_1 _10689_ (.Y(_04729_),
    .A(net1572),
    .B(net1667));
 sg13g2_nand2_1 _10690_ (.Y(_04730_),
    .A(net1576),
    .B(net1667));
 sg13g2_xor2_1 _10691_ (.B(_04730_),
    .A(_04608_),
    .X(_04731_));
 sg13g2_nand2b_1 _10692_ (.Y(_04732_),
    .B(_04731_),
    .A_N(_04728_));
 sg13g2_xnor2_1 _10693_ (.Y(_04733_),
    .A(_04728_),
    .B(_04731_));
 sg13g2_inv_1 _10694_ (.Y(_04734_),
    .A(_04733_));
 sg13g2_o21ai_1 _10695_ (.B1(_04619_),
    .Y(_04735_),
    .A1(_04491_),
    .A2(_04617_));
 sg13g2_nand2_1 _10696_ (.Y(_04736_),
    .A(net1579),
    .B(net1662));
 sg13g2_nand2_1 _10697_ (.Y(_04737_),
    .A(net1591),
    .B(net1655));
 sg13g2_xor2_1 _10698_ (.B(_04737_),
    .A(_04616_),
    .X(_04738_));
 sg13g2_nand2b_1 _10699_ (.Y(_04739_),
    .B(_04738_),
    .A_N(_04736_));
 sg13g2_xnor2_1 _10700_ (.Y(_04740_),
    .A(_04736_),
    .B(_04738_));
 sg13g2_nand2_1 _10701_ (.Y(_04741_),
    .A(_04735_),
    .B(_04740_));
 sg13g2_xnor2_1 _10702_ (.Y(_04742_),
    .A(_04735_),
    .B(_04740_));
 sg13g2_xnor2_1 _10703_ (.Y(_04743_),
    .A(_04733_),
    .B(_04742_));
 sg13g2_xnor2_1 _10704_ (.Y(_04744_),
    .A(_04727_),
    .B(_04743_));
 sg13g2_nor2b_1 _10705_ (.A(_04744_),
    .B_N(_04726_),
    .Y(_04745_));
 sg13g2_xor2_1 _10706_ (.B(_04744_),
    .A(_04726_),
    .X(_04746_));
 sg13g2_xor2_1 _10707_ (.B(_04746_),
    .A(_04725_),
    .X(_04747_));
 sg13g2_nand2_1 _10708_ (.Y(_04748_),
    .A(_04719_),
    .B(_04747_));
 sg13g2_xnor2_1 _10709_ (.Y(_04749_),
    .A(_04719_),
    .B(_04747_));
 sg13g2_o21ai_1 _10710_ (.B1(_04644_),
    .Y(_04750_),
    .A1(_04645_),
    .A2(_04663_));
 sg13g2_o21ai_1 _10711_ (.B1(_04625_),
    .Y(_04751_),
    .A1(_04606_),
    .A2(_04623_));
 sg13g2_a21o_1 _10712_ (.A2(_04640_),
    .A1(_04634_),
    .B1(_04642_),
    .X(_04752_));
 sg13g2_o21ai_1 _10713_ (.B1(_04638_),
    .Y(_04753_),
    .A1(_04635_),
    .A2(_04639_));
 sg13g2_o21ai_1 _10714_ (.B1(_04611_),
    .Y(_04754_),
    .A1(_04483_),
    .A2(_04609_));
 sg13g2_nand2_1 _10715_ (.Y(_04755_),
    .A(net1507),
    .B(net1693));
 sg13g2_nand2_1 _10716_ (.Y(_04756_),
    .A(net1512),
    .B(net1679));
 sg13g2_nand2_1 _10717_ (.Y(_04757_),
    .A(net1564),
    .B(net1683));
 sg13g2_or2_1 _10718_ (.X(_04758_),
    .B(_04756_),
    .A(_04637_));
 sg13g2_xnor2_1 _10719_ (.Y(_04759_),
    .A(_04636_),
    .B(_04757_));
 sg13g2_xor2_1 _10720_ (.B(_04759_),
    .A(_04755_),
    .X(_04760_));
 sg13g2_xnor2_1 _10721_ (.Y(_04761_),
    .A(_04754_),
    .B(_04760_));
 sg13g2_nor2b_1 _10722_ (.A(_04761_),
    .B_N(_04753_),
    .Y(_04762_));
 sg13g2_xor2_1 _10723_ (.B(_04761_),
    .A(_04753_),
    .X(_04763_));
 sg13g2_inv_1 _10724_ (.Y(_04764_),
    .A(_04763_));
 sg13g2_xnor2_1 _10725_ (.Y(_04765_),
    .A(_04752_),
    .B(_04764_));
 sg13g2_and2_1 _10726_ (.A(net1485),
    .B(net1722),
    .X(_04766_));
 sg13g2_nand2_1 _10727_ (.Y(_04767_),
    .A(net1492),
    .B(net1711));
 sg13g2_nand2_1 _10728_ (.Y(_04768_),
    .A(net1496),
    .B(net1711));
 sg13g2_xor2_1 _10729_ (.B(_04768_),
    .A(_04648_),
    .X(_04769_));
 sg13g2_nand2_1 _10730_ (.Y(_04770_),
    .A(_04766_),
    .B(_04769_));
 sg13g2_xor2_1 _10731_ (.B(_04769_),
    .A(_04766_),
    .X(_04771_));
 sg13g2_inv_1 _10732_ (.Y(_04772_),
    .A(_04771_));
 sg13g2_o21ai_1 _10733_ (.B1(_04659_),
    .Y(_04773_),
    .A1(_04530_),
    .A2(_04657_));
 sg13g2_nand2_1 _10734_ (.Y(_04774_),
    .A(net1497),
    .B(net1705));
 sg13g2_nand2_1 _10735_ (.Y(_04775_),
    .A(net1502),
    .B(net1698));
 sg13g2_nand2_1 _10736_ (.Y(_04776_),
    .A(net1503),
    .B(net1697));
 sg13g2_xor2_1 _10737_ (.B(_04776_),
    .A(_04656_),
    .X(_04777_));
 sg13g2_nand2b_1 _10738_ (.Y(_04778_),
    .B(_04777_),
    .A_N(_04774_));
 sg13g2_xnor2_1 _10739_ (.Y(_04779_),
    .A(_04774_),
    .B(_04777_));
 sg13g2_nand2_1 _10740_ (.Y(_04780_),
    .A(_04773_),
    .B(_04779_));
 sg13g2_xnor2_1 _10741_ (.Y(_04781_),
    .A(_04773_),
    .B(_04779_));
 sg13g2_xnor2_1 _10742_ (.Y(_04782_),
    .A(_04772_),
    .B(_04781_));
 sg13g2_nor2_1 _10743_ (.A(_04765_),
    .B(_04782_),
    .Y(_04783_));
 sg13g2_xor2_1 _10744_ (.B(_04782_),
    .A(_04765_),
    .X(_04784_));
 sg13g2_xnor2_1 _10745_ (.Y(_04785_),
    .A(_04751_),
    .B(_04784_));
 sg13g2_nor2b_1 _10746_ (.A(_04785_),
    .B_N(_04750_),
    .Y(_04786_));
 sg13g2_xor2_1 _10747_ (.B(_04785_),
    .A(_04750_),
    .X(_04787_));
 sg13g2_xor2_1 _10748_ (.B(_04787_),
    .A(_04749_),
    .X(_04788_));
 sg13g2_nand2_1 _10749_ (.Y(_04789_),
    .A(_04718_),
    .B(_04788_));
 sg13g2_xnor2_1 _10750_ (.Y(_04790_),
    .A(_04718_),
    .B(_04788_));
 sg13g2_o21ai_1 _10751_ (.B1(_04688_),
    .Y(_04791_),
    .A1(_04689_),
    .A2(_04696_));
 sg13g2_a21o_2 _10752_ (.A2(_04664_),
    .A1(_04631_),
    .B1(_04666_),
    .X(_04792_));
 sg13g2_o21ai_1 _10753_ (.B1(_04690_),
    .Y(_04793_),
    .A1(_03809_),
    .A2(_04691_));
 sg13g2_nand2_1 _10754_ (.Y(_04794_),
    .A(_04431_),
    .B(_04435_));
 sg13g2_xnor2_1 _10755_ (.Y(_04795_),
    .A(_04431_),
    .B(_04435_));
 sg13g2_xnor2_1 _10756_ (.Y(_04796_),
    .A(_04041_),
    .B(_04795_));
 sg13g2_nand2_1 _10757_ (.Y(_04797_),
    .A(_04793_),
    .B(_04796_));
 sg13g2_xnor2_1 _10758_ (.Y(_04798_),
    .A(_04793_),
    .B(_04796_));
 sg13g2_xnor2_1 _10759_ (.Y(_04799_),
    .A(_03807_),
    .B(_04798_));
 sg13g2_inv_1 _10760_ (.Y(_04800_),
    .A(_04799_));
 sg13g2_o21ai_1 _10761_ (.B1(_04686_),
    .Y(_04801_),
    .A1(_04676_),
    .A2(_04684_));
 sg13g2_a21o_1 _10762_ (.A2(_04681_),
    .A1(_04678_),
    .B1(_04683_),
    .X(_04802_));
 sg13g2_o21ai_1 _10763_ (.B1(_04661_),
    .Y(_04803_),
    .A1(_04653_),
    .A2(_04662_));
 sg13g2_inv_1 _10764_ (.Y(_04804_),
    .A(_04803_));
 sg13g2_o21ai_1 _10765_ (.B1(_04679_),
    .Y(_04805_),
    .A1(_04275_),
    .A2(_04680_));
 sg13g2_a21o_1 _10766_ (.A2(_04651_),
    .A1(_04646_),
    .B1(_04649_),
    .X(_04806_));
 sg13g2_nand2_1 _10767_ (.Y(_04807_),
    .A(net1729),
    .B(_04521_));
 sg13g2_o21ai_1 _10768_ (.B1(_04807_),
    .Y(_04808_),
    .A1(_04521_),
    .A2(_04646_));
 sg13g2_xnor2_1 _10769_ (.Y(_04809_),
    .A(_04398_),
    .B(_04808_));
 sg13g2_xnor2_1 _10770_ (.Y(_04810_),
    .A(_04806_),
    .B(_04809_));
 sg13g2_nor2b_1 _10771_ (.A(_04810_),
    .B_N(_04805_),
    .Y(_04811_));
 sg13g2_xor2_1 _10772_ (.B(_04810_),
    .A(_04805_),
    .X(_04812_));
 sg13g2_xor2_1 _10773_ (.B(_04812_),
    .A(_04803_),
    .X(_04813_));
 sg13g2_nand2b_1 _10774_ (.Y(_04814_),
    .B(_04802_),
    .A_N(_04813_));
 sg13g2_xor2_1 _10775_ (.B(_04813_),
    .A(_04802_),
    .X(_04815_));
 sg13g2_nand2b_1 _10776_ (.Y(_04816_),
    .B(_04801_),
    .A_N(_04815_));
 sg13g2_xor2_1 _10777_ (.B(_04815_),
    .A(_04801_),
    .X(_04817_));
 sg13g2_xnor2_1 _10778_ (.Y(_04818_),
    .A(_04800_),
    .B(_04817_));
 sg13g2_nor2b_1 _10779_ (.A(_04818_),
    .B_N(_04792_),
    .Y(_04819_));
 sg13g2_xor2_1 _10780_ (.B(_04818_),
    .A(_04792_),
    .X(_04820_));
 sg13g2_nor2b_1 _10781_ (.A(_04820_),
    .B_N(_04791_),
    .Y(_04821_));
 sg13g2_xor2_1 _10782_ (.B(_04820_),
    .A(_04791_),
    .X(_04822_));
 sg13g2_xor2_1 _10783_ (.B(_04822_),
    .A(_04790_),
    .X(_04823_));
 sg13g2_xnor2_1 _10784_ (.Y(_04824_),
    .A(_04717_),
    .B(_04823_));
 sg13g2_nor2_1 _10785_ (.A(_04716_),
    .B(_04824_),
    .Y(_04825_));
 sg13g2_xor2_1 _10786_ (.B(_04824_),
    .A(_04716_),
    .X(_04826_));
 sg13g2_nand2b_1 _10787_ (.Y(_04827_),
    .B(_04826_),
    .A_N(_04713_));
 sg13g2_xnor2_1 _10788_ (.Y(_04828_),
    .A(_04713_),
    .B(_04826_));
 sg13g2_nand2_1 _10789_ (.Y(_04829_),
    .A(_04586_),
    .B(_04828_));
 sg13g2_xor2_1 _10790_ (.B(_04828_),
    .A(_04586_),
    .X(_04830_));
 sg13g2_and2_1 _10791_ (.A(_04706_),
    .B(_04830_),
    .X(_04831_));
 sg13g2_xor2_1 _10792_ (.B(_04830_),
    .A(_04706_),
    .X(_04832_));
 sg13g2_o21ai_1 _10793_ (.B1(_04708_),
    .Y(_04833_),
    .A1(_04583_),
    .A2(_04710_));
 sg13g2_and2_1 _10794_ (.A(_04832_),
    .B(_04833_),
    .X(_04834_));
 sg13g2_xor2_1 _10795_ (.B(_04833_),
    .A(_04832_),
    .X(_04835_));
 sg13g2_o21ai_1 _10796_ (.B1(net1759),
    .Y(_04836_),
    .A1(net1401),
    .A2(_04835_));
 sg13g2_a21oi_1 _10797_ (.A1(net1401),
    .A2(_05542_),
    .Y(_00332_),
    .B1(_04836_));
 sg13g2_a21oi_1 _10798_ (.A1(_04832_),
    .A2(_04833_),
    .Y(_04837_),
    .B1(_04831_));
 sg13g2_a21oi_1 _10799_ (.A1(_04717_),
    .A2(_04823_),
    .Y(_04838_),
    .B1(_04825_));
 sg13g2_nor2_1 _10800_ (.A(_04819_),
    .B(_04821_),
    .Y(_04839_));
 sg13g2_o21ai_1 _10801_ (.B1(_04797_),
    .Y(_04840_),
    .A1(_03808_),
    .A2(_04798_));
 sg13g2_o21ai_1 _10802_ (.B1(_04840_),
    .Y(_04841_),
    .A1(_04819_),
    .A2(_04821_));
 sg13g2_xor2_1 _10803_ (.B(_04840_),
    .A(_04839_),
    .X(_04842_));
 sg13g2_o21ai_1 _10804_ (.B1(_04789_),
    .Y(_04843_),
    .A1(_04790_),
    .A2(_04822_));
 sg13g2_o21ai_1 _10805_ (.B1(_04748_),
    .Y(_04844_),
    .A1(_04749_),
    .A2(_04787_));
 sg13g2_o21ai_1 _10806_ (.B1(_04724_),
    .Y(_04845_),
    .A1(_04725_),
    .A2(_04746_));
 sg13g2_nand2b_1 _10807_ (.Y(_04846_),
    .B(_04722_),
    .A_N(_04339_));
 sg13g2_mux2_1 _10808_ (.A0(_04340_),
    .A1(_04339_),
    .S(_04722_),
    .X(_04847_));
 sg13g2_inv_2 _10809_ (.Y(_04848_),
    .A(_04847_));
 sg13g2_o21ai_1 _10810_ (.B1(_04741_),
    .Y(_04849_),
    .A1(_04734_),
    .A2(_04742_));
 sg13g2_o21ai_1 _10811_ (.B1(_04596_),
    .Y(_04850_),
    .A1(_04598_),
    .A2(_04721_));
 sg13g2_nand2_1 _10812_ (.Y(_04851_),
    .A(net1568),
    .B(net1670));
 sg13g2_nand2_1 _10813_ (.Y(_04852_),
    .A(net1572),
    .B(net1662));
 sg13g2_nand2_1 _10814_ (.Y(_04853_),
    .A(net1576),
    .B(net1662));
 sg13g2_xor2_1 _10815_ (.B(_04853_),
    .A(_04729_),
    .X(_04854_));
 sg13g2_nand2b_1 _10816_ (.Y(_04855_),
    .B(_04854_),
    .A_N(_04851_));
 sg13g2_xnor2_1 _10817_ (.Y(_04856_),
    .A(_04851_),
    .B(_04854_));
 sg13g2_inv_1 _10818_ (.Y(_04857_),
    .A(_04856_));
 sg13g2_o21ai_1 _10819_ (.B1(_04739_),
    .Y(_04858_),
    .A1(_04616_),
    .A2(_04737_));
 sg13g2_o21ai_1 _10820_ (.B1(net1655),
    .Y(_04859_),
    .A1(net1584),
    .A2(net1591));
 sg13g2_nand3_1 _10821_ (.B(net1591),
    .C(net1655),
    .A(net1584),
    .Y(_04860_));
 sg13g2_nand2b_1 _10822_ (.Y(_04861_),
    .B(_04860_),
    .A_N(_04859_));
 sg13g2_nand2_1 _10823_ (.Y(_04862_),
    .A(net1579),
    .B(net1659));
 sg13g2_xor2_1 _10824_ (.B(_04862_),
    .A(_04861_),
    .X(_04863_));
 sg13g2_nand2_1 _10825_ (.Y(_04864_),
    .A(_04858_),
    .B(_04863_));
 sg13g2_xnor2_1 _10826_ (.Y(_04865_),
    .A(_04858_),
    .B(_04863_));
 sg13g2_xnor2_1 _10827_ (.Y(_04866_),
    .A(_04856_),
    .B(_04865_));
 sg13g2_xnor2_1 _10828_ (.Y(_04867_),
    .A(_04850_),
    .B(_04866_));
 sg13g2_nor2b_1 _10829_ (.A(_04867_),
    .B_N(_04849_),
    .Y(_04868_));
 sg13g2_xor2_1 _10830_ (.B(_04867_),
    .A(_04849_),
    .X(_04869_));
 sg13g2_or2_1 _10831_ (.X(_04870_),
    .B(_04869_),
    .A(_04848_));
 sg13g2_xnor2_1 _10832_ (.Y(_04871_),
    .A(_04847_),
    .B(_04869_));
 sg13g2_nand2_1 _10833_ (.Y(_04872_),
    .A(_04845_),
    .B(_04871_));
 sg13g2_xnor2_1 _10834_ (.Y(_04873_),
    .A(_04845_),
    .B(_04871_));
 sg13g2_a21oi_1 _10835_ (.A1(_04752_),
    .A2(_04764_),
    .Y(_04874_),
    .B1(_04783_));
 sg13g2_a21o_1 _10836_ (.A2(_04743_),
    .A1(_04727_),
    .B1(_04745_),
    .X(_04875_));
 sg13g2_a21o_1 _10837_ (.A2(_04760_),
    .A1(_04754_),
    .B1(_04762_),
    .X(_04876_));
 sg13g2_o21ai_1 _10838_ (.B1(_04758_),
    .Y(_04877_),
    .A1(_04755_),
    .A2(_04759_));
 sg13g2_o21ai_1 _10839_ (.B1(_04732_),
    .Y(_04878_),
    .A1(_04608_),
    .A2(_04730_));
 sg13g2_nand2_1 _10840_ (.Y(_04879_),
    .A(net1507),
    .B(net1684));
 sg13g2_nand2_1 _10841_ (.Y(_04880_),
    .A(net1512),
    .B(net1674));
 sg13g2_nand2_1 _10842_ (.Y(_04881_),
    .A(net1564),
    .B(net1678));
 sg13g2_or2_1 _10843_ (.X(_04882_),
    .B(_04880_),
    .A(_04757_));
 sg13g2_xnor2_1 _10844_ (.Y(_04883_),
    .A(_04756_),
    .B(_04881_));
 sg13g2_xor2_1 _10845_ (.B(_04883_),
    .A(_04879_),
    .X(_04884_));
 sg13g2_xnor2_1 _10846_ (.Y(_04885_),
    .A(_04878_),
    .B(_04884_));
 sg13g2_nor2b_1 _10847_ (.A(_04885_),
    .B_N(_04877_),
    .Y(_04886_));
 sg13g2_xnor2_1 _10848_ (.Y(_04887_),
    .A(_04877_),
    .B(_04885_));
 sg13g2_nand2_1 _10849_ (.Y(_04888_),
    .A(_04876_),
    .B(_04887_));
 sg13g2_xnor2_1 _10850_ (.Y(_04889_),
    .A(_04876_),
    .B(_04887_));
 sg13g2_nand2_1 _10851_ (.Y(_04890_),
    .A(net1485),
    .B(net1716));
 sg13g2_nand2_1 _10852_ (.Y(_04891_),
    .A(net1496),
    .B(net1705));
 sg13g2_xor2_1 _10853_ (.B(_04891_),
    .A(_04767_),
    .X(_04892_));
 sg13g2_nand2b_1 _10854_ (.Y(_04893_),
    .B(_04892_),
    .A_N(_04890_));
 sg13g2_xor2_1 _10855_ (.B(_04892_),
    .A(_04890_),
    .X(_04894_));
 sg13g2_o21ai_1 _10856_ (.B1(_04778_),
    .Y(_04895_),
    .A1(_04656_),
    .A2(_04776_));
 sg13g2_nand2_1 _10857_ (.Y(_04896_),
    .A(net1497),
    .B(net1702));
 sg13g2_nand2_2 _10858_ (.Y(_04897_),
    .A(net1503),
    .B(net1693));
 sg13g2_xor2_1 _10859_ (.B(_04897_),
    .A(_04775_),
    .X(_04898_));
 sg13g2_nand2b_1 _10860_ (.Y(_04899_),
    .B(_04898_),
    .A_N(_04896_));
 sg13g2_xnor2_1 _10861_ (.Y(_04900_),
    .A(_04896_),
    .B(_04898_));
 sg13g2_nand2_1 _10862_ (.Y(_04901_),
    .A(_04895_),
    .B(_04900_));
 sg13g2_xnor2_1 _10863_ (.Y(_04902_),
    .A(_04895_),
    .B(_04900_));
 sg13g2_xnor2_1 _10864_ (.Y(_04903_),
    .A(_04894_),
    .B(_04902_));
 sg13g2_xor2_1 _10865_ (.B(_04903_),
    .A(_04889_),
    .X(_04904_));
 sg13g2_nand2_1 _10866_ (.Y(_04905_),
    .A(_04875_),
    .B(_04904_));
 sg13g2_xnor2_1 _10867_ (.Y(_04906_),
    .A(_04875_),
    .B(_04904_));
 sg13g2_xnor2_1 _10868_ (.Y(_04907_),
    .A(_04874_),
    .B(_04906_));
 sg13g2_xor2_1 _10869_ (.B(_04907_),
    .A(_04873_),
    .X(_04908_));
 sg13g2_nand2_1 _10870_ (.Y(_04909_),
    .A(_04844_),
    .B(_04908_));
 sg13g2_xnor2_1 _10871_ (.Y(_04910_),
    .A(_04844_),
    .B(_04908_));
 sg13g2_o21ai_1 _10872_ (.B1(_04816_),
    .Y(_04911_),
    .A1(_04800_),
    .A2(_04817_));
 sg13g2_a21o_2 _10873_ (.A2(_04784_),
    .A1(_04751_),
    .B1(_04786_),
    .X(_04912_));
 sg13g2_nand2b_2 _10874_ (.Y(_04913_),
    .B(net1558),
    .A_N(_04037_));
 sg13g2_o21ai_1 _10875_ (.B1(_04913_),
    .Y(_04914_),
    .A1(_03566_),
    .A2(_04038_));
 sg13g2_o21ai_1 _10876_ (.B1(_04794_),
    .Y(_04915_),
    .A1(_04042_),
    .A2(_04795_));
 sg13g2_nand2_1 _10877_ (.Y(_04916_),
    .A(_04551_),
    .B(_04555_));
 sg13g2_xnor2_1 _10878_ (.Y(_04917_),
    .A(_04551_),
    .B(_04555_));
 sg13g2_xnor2_1 _10879_ (.Y(_04918_),
    .A(_04174_),
    .B(_04917_));
 sg13g2_nand2_1 _10880_ (.Y(_04919_),
    .A(_04915_),
    .B(_04918_));
 sg13g2_xnor2_1 _10881_ (.Y(_04920_),
    .A(_04915_),
    .B(_04918_));
 sg13g2_xor2_1 _10882_ (.B(_04920_),
    .A(_04914_),
    .X(_04921_));
 sg13g2_o21ai_1 _10883_ (.B1(_04814_),
    .Y(_04922_),
    .A1(_04804_),
    .A2(_04812_));
 sg13g2_a21o_1 _10884_ (.A2(_04809_),
    .A1(_04806_),
    .B1(_04811_),
    .X(_04923_));
 sg13g2_o21ai_1 _10885_ (.B1(_04780_),
    .Y(_04924_),
    .A1(_04772_),
    .A2(_04781_));
 sg13g2_o21ai_1 _10886_ (.B1(_04807_),
    .Y(_04925_),
    .A1(_04399_),
    .A2(_04808_));
 sg13g2_o21ai_1 _10887_ (.B1(_04770_),
    .Y(_04926_),
    .A1(_04648_),
    .A2(_04768_));
 sg13g2_nand2_1 _10888_ (.Y(_04927_),
    .A(net1722),
    .B(_04646_));
 sg13g2_o21ai_1 _10889_ (.B1(_04927_),
    .Y(_04928_),
    .A1(_04646_),
    .A2(_04766_));
 sg13g2_xnor2_1 _10890_ (.Y(_04929_),
    .A(_04521_),
    .B(_04928_));
 sg13g2_xnor2_1 _10891_ (.Y(_04930_),
    .A(_04926_),
    .B(_04929_));
 sg13g2_nor2b_1 _10892_ (.A(_04930_),
    .B_N(_04925_),
    .Y(_04931_));
 sg13g2_xnor2_1 _10893_ (.Y(_04932_),
    .A(_04925_),
    .B(_04930_));
 sg13g2_xnor2_1 _10894_ (.Y(_04933_),
    .A(_04924_),
    .B(_04932_));
 sg13g2_nor2b_1 _10895_ (.A(_04933_),
    .B_N(_04923_),
    .Y(_04934_));
 sg13g2_xor2_1 _10896_ (.B(_04933_),
    .A(_04923_),
    .X(_04935_));
 sg13g2_nor2b_1 _10897_ (.A(_04935_),
    .B_N(_04922_),
    .Y(_04936_));
 sg13g2_xor2_1 _10898_ (.B(_04935_),
    .A(_04922_),
    .X(_04937_));
 sg13g2_inv_1 _10899_ (.Y(_04938_),
    .A(_04937_));
 sg13g2_xor2_1 _10900_ (.B(_04937_),
    .A(_04921_),
    .X(_04939_));
 sg13g2_nor2b_1 _10901_ (.A(_04939_),
    .B_N(_04912_),
    .Y(_04940_));
 sg13g2_xor2_1 _10902_ (.B(_04939_),
    .A(_04912_),
    .X(_04941_));
 sg13g2_nor2b_1 _10903_ (.A(_04941_),
    .B_N(_04911_),
    .Y(_04942_));
 sg13g2_xor2_1 _10904_ (.B(_04941_),
    .A(_04911_),
    .X(_04943_));
 sg13g2_xor2_1 _10905_ (.B(_04943_),
    .A(_04910_),
    .X(_04944_));
 sg13g2_xnor2_1 _10906_ (.Y(_04945_),
    .A(_04843_),
    .B(_04944_));
 sg13g2_nor2_1 _10907_ (.A(_04842_),
    .B(_04945_),
    .Y(_04946_));
 sg13g2_xor2_1 _10908_ (.B(_04945_),
    .A(_04842_),
    .X(_04947_));
 sg13g2_nor2b_1 _10909_ (.A(_04838_),
    .B_N(_04947_),
    .Y(_04948_));
 sg13g2_xnor2_1 _10910_ (.Y(_04949_),
    .A(_04838_),
    .B(_04947_));
 sg13g2_xnor2_1 _10911_ (.Y(_04950_),
    .A(_04715_),
    .B(_04949_));
 sg13g2_and3_1 _10912_ (.X(_04951_),
    .A(_04827_),
    .B(_04829_),
    .C(_04950_));
 sg13g2_nand3_1 _10913_ (.B(_04829_),
    .C(_04950_),
    .A(_04827_),
    .Y(_04952_));
 sg13g2_a21oi_1 _10914_ (.A1(_04827_),
    .A2(_04829_),
    .Y(_04953_),
    .B1(_04950_));
 sg13g2_nor2_1 _10915_ (.A(_04951_),
    .B(_04953_),
    .Y(_04954_));
 sg13g2_xnor2_1 _10916_ (.Y(_04955_),
    .A(_04837_),
    .B(_04954_));
 sg13g2_o21ai_1 _10917_ (.B1(net1759),
    .Y(_04956_),
    .A1(net1401),
    .A2(_04955_));
 sg13g2_a21oi_1 _10918_ (.A1(net1400),
    .A2(_05541_),
    .Y(_00333_),
    .B1(_04956_));
 sg13g2_or2_1 _10919_ (.X(_04957_),
    .B(_04953_),
    .A(_04831_));
 sg13g2_a22oi_1 _10920_ (.Y(_04958_),
    .B1(_04957_),
    .B2(_04952_),
    .A2(_04954_),
    .A1(_04834_));
 sg13g2_a21o_1 _10921_ (.A2(_04949_),
    .A1(_04715_),
    .B1(_04948_),
    .X(_04959_));
 sg13g2_a21oi_1 _10922_ (.A1(_04843_),
    .A2(_04944_),
    .Y(_04960_),
    .B1(_04946_));
 sg13g2_o21ai_1 _10923_ (.B1(_04909_),
    .Y(_04961_),
    .A1(_04910_),
    .A2(_04943_));
 sg13g2_o21ai_1 _10924_ (.B1(_04872_),
    .Y(_04962_),
    .A1(_04873_),
    .A2(_04907_));
 sg13g2_and2_1 _10925_ (.A(_04846_),
    .B(_04870_),
    .X(_04963_));
 sg13g2_o21ai_1 _10926_ (.B1(_04864_),
    .Y(_04964_),
    .A1(_04857_),
    .A2(_04865_));
 sg13g2_nand2_1 _10927_ (.Y(_04965_),
    .A(net1568),
    .B(net1667));
 sg13g2_nand2_1 _10928_ (.Y(_04966_),
    .A(net1572),
    .B(net1658));
 sg13g2_nand2_1 _10929_ (.Y(_04967_),
    .A(net1576),
    .B(net1658));
 sg13g2_xor2_1 _10930_ (.B(_04967_),
    .A(_04852_),
    .X(_04968_));
 sg13g2_nand2b_1 _10931_ (.Y(_04969_),
    .B(_04968_),
    .A_N(_04965_));
 sg13g2_xnor2_1 _10932_ (.Y(_04970_),
    .A(_04965_),
    .B(_04968_));
 sg13g2_o21ai_1 _10933_ (.B1(_04860_),
    .Y(_04971_),
    .A1(_04859_),
    .A2(_04862_));
 sg13g2_nand2_1 _10934_ (.Y(_04972_),
    .A(net1579),
    .B(net1656));
 sg13g2_xnor2_1 _10935_ (.Y(_04973_),
    .A(_04861_),
    .B(_04972_));
 sg13g2_and4_1 _10936_ (.A(net1579),
    .B(net1584),
    .C(net1591),
    .D(net1656),
    .X(_04974_));
 sg13g2_xnor2_1 _10937_ (.Y(_04975_),
    .A(_04971_),
    .B(_04973_));
 sg13g2_xor2_1 _10938_ (.B(_04975_),
    .A(_04970_),
    .X(_04976_));
 sg13g2_xnor2_1 _10939_ (.Y(_04977_),
    .A(_04850_),
    .B(_04976_));
 sg13g2_nor2b_1 _10940_ (.A(_04977_),
    .B_N(_04964_),
    .Y(_04978_));
 sg13g2_xor2_1 _10941_ (.B(_04977_),
    .A(_04964_),
    .X(_04979_));
 sg13g2_xnor2_1 _10942_ (.Y(_04980_),
    .A(_04848_),
    .B(_04979_));
 sg13g2_nor2_1 _10943_ (.A(_04963_),
    .B(_04980_),
    .Y(_04981_));
 sg13g2_xor2_1 _10944_ (.B(_04980_),
    .A(_04963_),
    .X(_04982_));
 sg13g2_o21ai_1 _10945_ (.B1(_04888_),
    .Y(_04983_),
    .A1(_04889_),
    .A2(_04903_));
 sg13g2_a21oi_1 _10946_ (.A1(_04850_),
    .A2(_04866_),
    .Y(_04984_),
    .B1(_04868_));
 sg13g2_a21o_1 _10947_ (.A2(_04884_),
    .A1(_04878_),
    .B1(_04886_),
    .X(_04985_));
 sg13g2_o21ai_1 _10948_ (.B1(_04882_),
    .Y(_04986_),
    .A1(_04879_),
    .A2(_04883_));
 sg13g2_o21ai_1 _10949_ (.B1(_04855_),
    .Y(_04987_),
    .A1(_04729_),
    .A2(_04853_));
 sg13g2_nand2_1 _10950_ (.Y(_04988_),
    .A(net1507),
    .B(net1683));
 sg13g2_nand2_1 _10951_ (.Y(_04989_),
    .A(net1512),
    .B(\cordic_inst.MUX_cordic_state$write_1__VAL_1[75] ));
 sg13g2_nand2_1 _10952_ (.Y(_04990_),
    .A(net1564),
    .B(net1670));
 sg13g2_xor2_1 _10953_ (.B(_04990_),
    .A(_04880_),
    .X(_04991_));
 sg13g2_nand2b_1 _10954_ (.Y(_04992_),
    .B(_04991_),
    .A_N(_04988_));
 sg13g2_xnor2_1 _10955_ (.Y(_04993_),
    .A(_04988_),
    .B(_04991_));
 sg13g2_xnor2_1 _10956_ (.Y(_04994_),
    .A(_04987_),
    .B(_04993_));
 sg13g2_nor2b_1 _10957_ (.A(_04994_),
    .B_N(_04986_),
    .Y(_04995_));
 sg13g2_xnor2_1 _10958_ (.Y(_04996_),
    .A(_04986_),
    .B(_04994_));
 sg13g2_nand2_1 _10959_ (.Y(_04997_),
    .A(_04985_),
    .B(_04996_));
 sg13g2_xnor2_1 _10960_ (.Y(_04998_),
    .A(_04985_),
    .B(_04996_));
 sg13g2_nand2_1 _10961_ (.Y(_04999_),
    .A(net1485),
    .B(net1711));
 sg13g2_nand2_1 _10962_ (.Y(_05000_),
    .A(net1492),
    .B(net1702));
 sg13g2_nor2_1 _10963_ (.A(_04891_),
    .B(_05000_),
    .Y(_05001_));
 sg13g2_a22oi_1 _10964_ (.Y(_05002_),
    .B1(net1705),
    .B2(net1492),
    .A2(net1702),
    .A1(net1496));
 sg13g2_nor3_1 _10965_ (.A(_04999_),
    .B(_05001_),
    .C(_05002_),
    .Y(_05003_));
 sg13g2_o21ai_1 _10966_ (.B1(_04999_),
    .Y(_05004_),
    .A1(_05001_),
    .A2(_05002_));
 sg13g2_nand2b_1 _10967_ (.Y(_05005_),
    .B(_05004_),
    .A_N(_05003_));
 sg13g2_o21ai_1 _10968_ (.B1(_04899_),
    .Y(_05006_),
    .A1(_04775_),
    .A2(_04897_));
 sg13g2_nand2_1 _10969_ (.Y(_05007_),
    .A(net1497),
    .B(net1698));
 sg13g2_nand2_1 _10970_ (.Y(_05008_),
    .A(net1502),
    .B(net1684));
 sg13g2_nor2_1 _10971_ (.A(_04897_),
    .B(_05008_),
    .Y(_05009_));
 sg13g2_or2_1 _10972_ (.X(_05010_),
    .B(_05008_),
    .A(_04897_));
 sg13g2_a22oi_1 _10973_ (.Y(_05011_),
    .B1(net1693),
    .B2(net1502),
    .A2(net1684),
    .A1(net1503));
 sg13g2_nor2_1 _10974_ (.A(_05009_),
    .B(_05011_),
    .Y(_05012_));
 sg13g2_xnor2_1 _10975_ (.Y(_05013_),
    .A(_05007_),
    .B(_05012_));
 sg13g2_nand2_1 _10976_ (.Y(_05014_),
    .A(_05006_),
    .B(_05013_));
 sg13g2_xnor2_1 _10977_ (.Y(_05015_),
    .A(_05006_),
    .B(_05013_));
 sg13g2_xnor2_1 _10978_ (.Y(_05016_),
    .A(_05005_),
    .B(_05015_));
 sg13g2_xnor2_1 _10979_ (.Y(_05017_),
    .A(_04998_),
    .B(_05016_));
 sg13g2_nor2_1 _10980_ (.A(_04984_),
    .B(_05017_),
    .Y(_05018_));
 sg13g2_xor2_1 _10981_ (.B(_05017_),
    .A(_04984_),
    .X(_05019_));
 sg13g2_xnor2_1 _10982_ (.Y(_05020_),
    .A(_04983_),
    .B(_05019_));
 sg13g2_inv_1 _10983_ (.Y(_05021_),
    .A(_05020_));
 sg13g2_xnor2_1 _10984_ (.Y(_05022_),
    .A(_04982_),
    .B(_05020_));
 sg13g2_nand2_1 _10985_ (.Y(_05023_),
    .A(_04962_),
    .B(_05022_));
 sg13g2_xnor2_1 _10986_ (.Y(_05024_),
    .A(_04962_),
    .B(_05022_));
 sg13g2_a21oi_1 _10987_ (.A1(_04921_),
    .A2(_04938_),
    .Y(_05025_),
    .B1(_04936_));
 sg13g2_o21ai_1 _10988_ (.B1(_04905_),
    .Y(_05026_),
    .A1(_04874_),
    .A2(_04906_));
 sg13g2_nor2b_1 _10989_ (.A(_03809_),
    .B_N(_04303_),
    .Y(_05027_));
 sg13g2_xor2_1 _10990_ (.B(_04303_),
    .A(_03809_),
    .X(_05028_));
 sg13g2_o21ai_1 _10991_ (.B1(_04916_),
    .Y(_05029_),
    .A1(_04175_),
    .A2(_04917_));
 sg13g2_nand2_1 _10992_ (.Y(_05030_),
    .A(_04677_),
    .B(_04681_));
 sg13g2_xnor2_1 _10993_ (.Y(_05031_),
    .A(_04677_),
    .B(_04681_));
 sg13g2_xnor2_1 _10994_ (.Y(_05032_),
    .A(_04307_),
    .B(_05031_));
 sg13g2_xnor2_1 _10995_ (.Y(_05033_),
    .A(_05029_),
    .B(_05032_));
 sg13g2_nor2_1 _10996_ (.A(_05028_),
    .B(_05033_),
    .Y(_05034_));
 sg13g2_xnor2_1 _10997_ (.Y(_05035_),
    .A(_05028_),
    .B(_05033_));
 sg13g2_a21o_1 _10998_ (.A2(_04932_),
    .A1(_04924_),
    .B1(_04934_),
    .X(_05036_));
 sg13g2_a21o_1 _10999_ (.A2(_04929_),
    .A1(_04926_),
    .B1(_04931_),
    .X(_05037_));
 sg13g2_o21ai_1 _11000_ (.B1(_04901_),
    .Y(_05038_),
    .A1(_04894_),
    .A2(_04902_));
 sg13g2_o21ai_1 _11001_ (.B1(_04927_),
    .Y(_05039_),
    .A1(_04522_),
    .A2(_04928_));
 sg13g2_o21ai_1 _11002_ (.B1(_04893_),
    .Y(_05040_),
    .A1(_04767_),
    .A2(_04891_));
 sg13g2_o21ai_1 _11003_ (.B1(net1485),
    .Y(_05041_),
    .A1(net1716),
    .A2(net1722));
 sg13g2_nand2_1 _11004_ (.Y(_05042_),
    .A(net1716),
    .B(_04766_));
 sg13g2_nand2b_1 _11005_ (.Y(_05043_),
    .B(_05042_),
    .A_N(_05041_));
 sg13g2_xnor2_1 _11006_ (.Y(_05044_),
    .A(_04646_),
    .B(_05043_));
 sg13g2_xnor2_1 _11007_ (.Y(_05045_),
    .A(_05040_),
    .B(_05044_));
 sg13g2_nor2b_1 _11008_ (.A(_05045_),
    .B_N(_05039_),
    .Y(_05046_));
 sg13g2_xnor2_1 _11009_ (.Y(_05047_),
    .A(_05039_),
    .B(_05045_));
 sg13g2_xnor2_1 _11010_ (.Y(_05048_),
    .A(_05038_),
    .B(_05047_));
 sg13g2_nor2b_1 _11011_ (.A(_05048_),
    .B_N(_05037_),
    .Y(_05049_));
 sg13g2_xnor2_1 _11012_ (.Y(_05050_),
    .A(_05037_),
    .B(_05048_));
 sg13g2_xnor2_1 _11013_ (.Y(_05051_),
    .A(_05036_),
    .B(_05050_));
 sg13g2_nor2_1 _11014_ (.A(_05035_),
    .B(_05051_),
    .Y(_05052_));
 sg13g2_xor2_1 _11015_ (.B(_05051_),
    .A(_05035_),
    .X(_05053_));
 sg13g2_nand2_1 _11016_ (.Y(_05054_),
    .A(_05026_),
    .B(_05053_));
 sg13g2_xnor2_1 _11017_ (.Y(_05055_),
    .A(_05026_),
    .B(_05053_));
 sg13g2_xnor2_1 _11018_ (.Y(_05056_),
    .A(_05025_),
    .B(_05055_));
 sg13g2_xor2_1 _11019_ (.B(_05056_),
    .A(_05024_),
    .X(_05057_));
 sg13g2_and2_1 _11020_ (.A(_04961_),
    .B(_05057_),
    .X(_05058_));
 sg13g2_or2_1 _11021_ (.X(_05059_),
    .B(_05057_),
    .A(_04961_));
 sg13g2_nand2b_1 _11022_ (.Y(_05060_),
    .B(_05059_),
    .A_N(_05058_));
 sg13g2_nor2_1 _11023_ (.A(_04940_),
    .B(_04942_),
    .Y(_05061_));
 sg13g2_o21ai_1 _11024_ (.B1(_04919_),
    .Y(_05062_),
    .A1(_04914_),
    .A2(_04920_));
 sg13g2_o21ai_1 _11025_ (.B1(_05062_),
    .Y(_05063_),
    .A1(_04940_),
    .A2(_04942_));
 sg13g2_xnor2_1 _11026_ (.Y(_05064_),
    .A(_05061_),
    .B(_05062_));
 sg13g2_nand2b_1 _11027_ (.Y(_05065_),
    .B(_05064_),
    .A_N(_04913_));
 sg13g2_xnor2_1 _11028_ (.Y(_05066_),
    .A(_04913_),
    .B(_05064_));
 sg13g2_xnor2_1 _11029_ (.Y(_05067_),
    .A(_05060_),
    .B(_05066_));
 sg13g2_nand2b_1 _11030_ (.Y(_05068_),
    .B(_05067_),
    .A_N(_04960_));
 sg13g2_xnor2_1 _11031_ (.Y(_05069_),
    .A(_04960_),
    .B(_05067_));
 sg13g2_nand2b_1 _11032_ (.Y(_05070_),
    .B(_05069_),
    .A_N(_04841_));
 sg13g2_xnor2_1 _11033_ (.Y(_05071_),
    .A(_04841_),
    .B(_05069_));
 sg13g2_nand2_1 _11034_ (.Y(_05072_),
    .A(_04959_),
    .B(_05071_));
 sg13g2_xnor2_1 _11035_ (.Y(_05073_),
    .A(_04959_),
    .B(_05071_));
 sg13g2_xor2_1 _11036_ (.B(_05073_),
    .A(_04958_),
    .X(_05074_));
 sg13g2_o21ai_1 _11037_ (.B1(net1759),
    .Y(_05075_),
    .A1(net1400),
    .A2(_05074_));
 sg13g2_a21oi_1 _11038_ (.A1(net1401),
    .A2(_05540_),
    .Y(_00334_),
    .B1(_05075_));
 sg13g2_o21ai_1 _11039_ (.B1(_05072_),
    .Y(_05076_),
    .A1(_04958_),
    .A2(_05073_));
 sg13g2_nand2_1 _11040_ (.Y(_05077_),
    .A(_05068_),
    .B(_05070_));
 sg13g2_nand2_1 _11041_ (.Y(_05078_),
    .A(_05063_),
    .B(_05065_));
 sg13g2_a21oi_1 _11042_ (.A1(_05059_),
    .A2(_05066_),
    .Y(_05079_),
    .B1(_05058_));
 sg13g2_a21oi_1 _11043_ (.A1(_04983_),
    .A2(_05019_),
    .Y(_05080_),
    .B1(_05018_));
 sg13g2_a21oi_1 _11044_ (.A1(_05038_),
    .A2(_05047_),
    .Y(_05081_),
    .B1(_05049_));
 sg13g2_a21oi_1 _11045_ (.A1(_05040_),
    .A2(_05044_),
    .Y(_05082_),
    .B1(_05046_));
 sg13g2_xor2_1 _11046_ (.B(_05082_),
    .A(_05081_),
    .X(_05083_));
 sg13g2_o21ai_1 _11047_ (.B1(_05030_),
    .Y(_05084_),
    .A1(_04308_),
    .A2(_05031_));
 sg13g2_xor2_1 _11048_ (.B(_04805_),
    .A(_04435_),
    .X(_05085_));
 sg13g2_xnor2_1 _11049_ (.Y(_05086_),
    .A(_05084_),
    .B(_05085_));
 sg13g2_o21ai_1 _11050_ (.B1(_05042_),
    .Y(_05087_),
    .A1(_04647_),
    .A2(_05041_));
 sg13g2_or2_1 _11051_ (.X(_05088_),
    .B(_05003_),
    .A(_05001_));
 sg13g2_xnor2_1 _11052_ (.Y(_05089_),
    .A(_04999_),
    .B(_05043_));
 sg13g2_xnor2_1 _11053_ (.Y(_05090_),
    .A(_05088_),
    .B(_05089_));
 sg13g2_xnor2_1 _11054_ (.Y(_05091_),
    .A(_05087_),
    .B(_05090_));
 sg13g2_xor2_1 _11055_ (.B(_04431_),
    .A(_04426_),
    .X(_05092_));
 sg13g2_xnor2_1 _11056_ (.Y(_05093_),
    .A(_05091_),
    .B(_05092_));
 sg13g2_o21ai_1 _11057_ (.B1(_05014_),
    .Y(_05094_),
    .A1(_05005_),
    .A2(_05015_));
 sg13g2_xor2_1 _11058_ (.B(_05094_),
    .A(_04809_),
    .X(_05095_));
 sg13g2_xnor2_1 _11059_ (.Y(_05096_),
    .A(_05093_),
    .B(_05095_));
 sg13g2_xnor2_1 _11060_ (.Y(_05097_),
    .A(_05086_),
    .B(_05096_));
 sg13g2_xnor2_1 _11061_ (.Y(_05098_),
    .A(_05083_),
    .B(_05097_));
 sg13g2_xnor2_1 _11062_ (.Y(_05099_),
    .A(_05080_),
    .B(_05098_));
 sg13g2_o21ai_1 _11063_ (.B1(_04992_),
    .Y(_05100_),
    .A1(_04880_),
    .A2(_04990_));
 sg13g2_a21oi_1 _11064_ (.A1(_04987_),
    .A2(_04993_),
    .Y(_05101_),
    .B1(_04995_));
 sg13g2_xnor2_1 _11065_ (.Y(_05102_),
    .A(_05100_),
    .B(_05101_));
 sg13g2_o21ai_1 _11066_ (.B1(_04969_),
    .Y(_05103_),
    .A1(_04852_),
    .A2(_04967_));
 sg13g2_nand2_1 _11067_ (.Y(_05104_),
    .A(net1486),
    .B(net1705));
 sg13g2_xnor2_1 _11068_ (.Y(_05105_),
    .A(_05103_),
    .B(_05104_));
 sg13g2_nand2_1 _11069_ (.Y(_05106_),
    .A(net1497),
    .B(net1693));
 sg13g2_nand2_1 _11070_ (.Y(_05107_),
    .A(net1496),
    .B(net1698));
 sg13g2_xnor2_1 _11071_ (.Y(_05108_),
    .A(_05000_),
    .B(_05107_));
 sg13g2_nand2_1 _11072_ (.Y(_05109_),
    .A(net1503),
    .B(net1679));
 sg13g2_xor2_1 _11073_ (.B(_05109_),
    .A(_05008_),
    .X(_05110_));
 sg13g2_xnor2_1 _11074_ (.Y(_05111_),
    .A(_05108_),
    .B(_05110_));
 sg13g2_xnor2_1 _11075_ (.Y(_05112_),
    .A(_05106_),
    .B(_05111_));
 sg13g2_o21ai_1 _11076_ (.B1(_05010_),
    .Y(_05113_),
    .A1(_05007_),
    .A2(_05011_));
 sg13g2_nand2_1 _11077_ (.Y(_05114_),
    .A(net1507),
    .B(net1678));
 sg13g2_nand2_1 _11078_ (.Y(_05115_),
    .A(net1565),
    .B(net1666));
 sg13g2_xor2_1 _11079_ (.B(_05115_),
    .A(_04989_),
    .X(_05116_));
 sg13g2_xnor2_1 _11080_ (.Y(_05117_),
    .A(_05114_),
    .B(_05116_));
 sg13g2_xnor2_1 _11081_ (.Y(_05118_),
    .A(_05113_),
    .B(_05117_));
 sg13g2_xnor2_1 _11082_ (.Y(_05119_),
    .A(_05112_),
    .B(_05118_));
 sg13g2_xnor2_1 _11083_ (.Y(_05120_),
    .A(_05105_),
    .B(_05119_));
 sg13g2_xnor2_1 _11084_ (.Y(_05121_),
    .A(_05102_),
    .B(_05120_));
 sg13g2_nand2_1 _11085_ (.Y(_05122_),
    .A(net1568),
    .B(net1665));
 sg13g2_nand2_1 _11086_ (.Y(_05123_),
    .A(net1576),
    .B(net1655));
 sg13g2_xnor2_1 _11087_ (.Y(_05124_),
    .A(_04966_),
    .B(_05123_));
 sg13g2_xnor2_1 _11088_ (.Y(_05125_),
    .A(_05122_),
    .B(_05124_));
 sg13g2_a21oi_1 _11089_ (.A1(_04970_),
    .A2(_04975_),
    .Y(_05126_),
    .B1(_04974_));
 sg13g2_xnor2_1 _11090_ (.Y(_05127_),
    .A(_05125_),
    .B(_05126_));
 sg13g2_a21oi_1 _11091_ (.A1(_04859_),
    .A2(_04972_),
    .Y(_05128_),
    .B1(_04974_));
 sg13g2_xor2_1 _11092_ (.B(_05128_),
    .A(_04850_),
    .X(_05129_));
 sg13g2_xnor2_1 _11093_ (.Y(_05130_),
    .A(_05127_),
    .B(_05129_));
 sg13g2_xnor2_1 _11094_ (.Y(_05131_),
    .A(_05121_),
    .B(_05130_));
 sg13g2_a21oi_1 _11095_ (.A1(_04850_),
    .A2(_04976_),
    .Y(_05132_),
    .B1(_04978_));
 sg13g2_xnor2_1 _11096_ (.Y(_05133_),
    .A(_04848_),
    .B(_05132_));
 sg13g2_xnor2_1 _11097_ (.Y(_05134_),
    .A(_05131_),
    .B(_05133_));
 sg13g2_o21ai_1 _11098_ (.B1(_04846_),
    .Y(_05135_),
    .A1(_04848_),
    .A2(_04979_));
 sg13g2_o21ai_1 _11099_ (.B1(_04997_),
    .Y(_05136_),
    .A1(_04998_),
    .A2(_05016_));
 sg13g2_xnor2_1 _11100_ (.Y(_05137_),
    .A(_05135_),
    .B(_05136_));
 sg13g2_xnor2_1 _11101_ (.Y(_05138_),
    .A(_05134_),
    .B(_05137_));
 sg13g2_xnor2_1 _11102_ (.Y(_05139_),
    .A(_05099_),
    .B(_05138_));
 sg13g2_a21oi_1 _11103_ (.A1(_05036_),
    .A2(_05050_),
    .Y(_05140_),
    .B1(_05052_));
 sg13g2_a21oi_1 _11104_ (.A1(_05029_),
    .A2(_05032_),
    .Y(_05141_),
    .B1(_05034_));
 sg13g2_a21oi_1 _11105_ (.A1(_04982_),
    .A2(_05021_),
    .Y(_05142_),
    .B1(_04981_));
 sg13g2_o21ai_1 _11106_ (.B1(_05054_),
    .Y(_05143_),
    .A1(_05025_),
    .A2(_05055_));
 sg13g2_xnor2_1 _11107_ (.Y(_05144_),
    .A(_05140_),
    .B(_05142_));
 sg13g2_xnor2_1 _11108_ (.Y(_05145_),
    .A(_05139_),
    .B(_05144_));
 sg13g2_xnor2_1 _11109_ (.Y(_05146_),
    .A(_05141_),
    .B(_05143_));
 sg13g2_xnor2_1 _11110_ (.Y(_05147_),
    .A(_05145_),
    .B(_05146_));
 sg13g2_o21ai_1 _11111_ (.B1(_05023_),
    .Y(_05148_),
    .A1(_05024_),
    .A2(_05056_));
 sg13g2_xnor2_1 _11112_ (.Y(_05149_),
    .A(_05027_),
    .B(_05148_));
 sg13g2_xnor2_1 _11113_ (.Y(_05150_),
    .A(_05147_),
    .B(_05149_));
 sg13g2_xnor2_1 _11114_ (.Y(_05151_),
    .A(_05079_),
    .B(_05150_));
 sg13g2_xnor2_1 _11115_ (.Y(_05152_),
    .A(_05078_),
    .B(_05151_));
 sg13g2_xnor2_1 _11116_ (.Y(_05153_),
    .A(_05077_),
    .B(_05152_));
 sg13g2_xnor2_1 _11117_ (.Y(_05154_),
    .A(_05076_),
    .B(_05153_));
 sg13g2_o21ai_1 _11118_ (.B1(net1759),
    .Y(_05155_),
    .A1(net658),
    .A2(net1472));
 sg13g2_a21oi_1 _11119_ (.A1(net1472),
    .A2(_05154_),
    .Y(_00335_),
    .B1(net659));
 sg13g2_nand2_1 _11120_ (.Y(_05156_),
    .A(net733),
    .B(_02447_));
 sg13g2_xor2_1 _11121_ (.B(_02447_),
    .A(net733),
    .X(_05157_));
 sg13g2_nor3_2 _11122_ (.A(net1466),
    .B(mac_en_mac),
    .C(mac_en_clear),
    .Y(_05158_));
 sg13g2_or3_1 _11123_ (.A(net1466),
    .B(mac_en_mac),
    .C(mac_en_clear),
    .X(_05159_));
 sg13g2_a22oi_1 _11124_ (.Y(_05160_),
    .B1(net1340),
    .B2(net476),
    .A2(_05157_),
    .A1(net1466));
 sg13g2_nor2_1 _11125_ (.A(net1741),
    .B(net477),
    .Y(_00336_));
 sg13g2_nor2b_1 _11126_ (.A(net733),
    .B_N(_02447_),
    .Y(_05161_));
 sg13g2_nand2b_1 _11127_ (.Y(_05162_),
    .B(\mac_inst.accumulator[1] ),
    .A_N(_02527_));
 sg13g2_nand2_1 _11128_ (.Y(_05163_),
    .A(\mac_inst.accumulator[1] ),
    .B(_02527_));
 sg13g2_xnor2_1 _11129_ (.Y(_05164_),
    .A(\mac_inst.accumulator[1] ),
    .B(_02527_));
 sg13g2_xor2_1 _11130_ (.B(_02527_),
    .A(\mac_inst.accumulator[1] ),
    .X(_05165_));
 sg13g2_o21ai_1 _11131_ (.B1(net1466),
    .Y(_05166_),
    .A1(_05161_),
    .A2(_05164_));
 sg13g2_a21o_1 _11132_ (.A2(_05164_),
    .A1(_05161_),
    .B1(_05166_),
    .X(_05167_));
 sg13g2_nand2_1 _11133_ (.Y(_05168_),
    .A(net365),
    .B(net1340));
 sg13g2_a21oi_1 _11134_ (.A1(_05167_),
    .A2(net366),
    .Y(_00337_),
    .B1(net1744));
 sg13g2_o21ai_1 _11135_ (.B1(_05163_),
    .Y(_05169_),
    .A1(_05161_),
    .A2(_05164_));
 sg13g2_nor2b_1 _11136_ (.A(_02619_),
    .B_N(\mac_inst.accumulator[2] ),
    .Y(_05170_));
 sg13g2_and2_1 _11137_ (.A(\mac_inst.accumulator[2] ),
    .B(_02619_),
    .X(_05171_));
 sg13g2_xnor2_1 _11138_ (.Y(_05172_),
    .A(net726),
    .B(_02619_));
 sg13g2_xor2_1 _11139_ (.B(_02619_),
    .A(\mac_inst.accumulator[2] ),
    .X(_05173_));
 sg13g2_a21oi_1 _11140_ (.A1(_05169_),
    .A2(_05172_),
    .Y(_05174_),
    .B1(net1384));
 sg13g2_o21ai_1 _11141_ (.B1(_05174_),
    .Y(_05175_),
    .A1(_05169_),
    .A2(_05172_));
 sg13g2_nand2_1 _11142_ (.Y(_05176_),
    .A(net408),
    .B(net1337));
 sg13g2_a21oi_1 _11143_ (.A1(_05175_),
    .A2(net409),
    .Y(_00338_),
    .B1(net1739));
 sg13g2_a21oi_1 _11144_ (.A1(_05169_),
    .A2(_05172_),
    .Y(_05177_),
    .B1(_05170_));
 sg13g2_nor2_1 _11145_ (.A(_05538_),
    .B(_02711_),
    .Y(_05178_));
 sg13g2_nand2_1 _11146_ (.Y(_05179_),
    .A(\mac_inst.accumulator[3] ),
    .B(_02711_));
 sg13g2_xnor2_1 _11147_ (.Y(_05180_),
    .A(\mac_inst.accumulator[3] ),
    .B(_02711_));
 sg13g2_a21oi_1 _11148_ (.A1(_05177_),
    .A2(_05180_),
    .Y(_05181_),
    .B1(net1384));
 sg13g2_o21ai_1 _11149_ (.B1(_05181_),
    .Y(_05182_),
    .A1(_05177_),
    .A2(_05180_));
 sg13g2_nand2_1 _11150_ (.Y(_05183_),
    .A(net522),
    .B(net1334));
 sg13g2_a21oi_1 _11151_ (.A1(_05182_),
    .A2(_05183_),
    .Y(_00339_),
    .B1(net1743));
 sg13g2_o21ai_1 _11152_ (.B1(_05179_),
    .Y(_05184_),
    .A1(_05177_),
    .A2(_05180_));
 sg13g2_nor2_1 _11153_ (.A(_05537_),
    .B(_02820_),
    .Y(_05185_));
 sg13g2_and2_1 _11154_ (.A(\mac_inst.accumulator[4] ),
    .B(_02820_),
    .X(_05186_));
 sg13g2_xnor2_1 _11155_ (.Y(_05187_),
    .A(_05537_),
    .B(_02820_));
 sg13g2_inv_1 _11156_ (.Y(_05188_),
    .A(_05187_));
 sg13g2_a21oi_1 _11157_ (.A1(_05184_),
    .A2(_05187_),
    .Y(_05189_),
    .B1(net1383));
 sg13g2_o21ai_1 _11158_ (.B1(_05189_),
    .Y(_05190_),
    .A1(_05184_),
    .A2(_05187_));
 sg13g2_nand2_1 _11159_ (.Y(_05191_),
    .A(net420),
    .B(net1335));
 sg13g2_a21oi_1 _11160_ (.A1(_05190_),
    .A2(net421),
    .Y(_00340_),
    .B1(net1737));
 sg13g2_a21oi_1 _11161_ (.A1(_05184_),
    .A2(_05187_),
    .Y(_05192_),
    .B1(_05186_));
 sg13g2_or2_1 _11162_ (.X(_05193_),
    .B(_02926_),
    .A(_05536_));
 sg13g2_nand2_1 _11163_ (.Y(_05194_),
    .A(\mac_inst.accumulator[5] ),
    .B(_02926_));
 sg13g2_xnor2_1 _11164_ (.Y(_05195_),
    .A(\mac_inst.accumulator[5] ),
    .B(_02926_));
 sg13g2_xnor2_1 _11165_ (.Y(_05196_),
    .A(_05536_),
    .B(_02926_));
 sg13g2_o21ai_1 _11166_ (.B1(net1468),
    .Y(_05197_),
    .A1(_05192_),
    .A2(_05195_));
 sg13g2_a21oi_1 _11167_ (.A1(_05192_),
    .A2(_05195_),
    .Y(_05198_),
    .B1(_05197_));
 sg13g2_a21oi_1 _11168_ (.A1(net487),
    .A2(net1331),
    .Y(_05199_),
    .B1(_05198_));
 sg13g2_nor2_1 _11169_ (.A(net1737),
    .B(net488),
    .Y(_00341_));
 sg13g2_o21ai_1 _11170_ (.B1(_05194_),
    .Y(_05200_),
    .A1(_05192_),
    .A2(_05195_));
 sg13g2_nor2b_1 _11171_ (.A(_03043_),
    .B_N(\mac_inst.accumulator[6] ),
    .Y(_05201_));
 sg13g2_and2_1 _11172_ (.A(\mac_inst.accumulator[6] ),
    .B(_03043_),
    .X(_05202_));
 sg13g2_xnor2_1 _11173_ (.Y(_05203_),
    .A(\mac_inst.accumulator[6] ),
    .B(_03043_));
 sg13g2_inv_1 _11174_ (.Y(_05204_),
    .A(_05203_));
 sg13g2_a21oi_1 _11175_ (.A1(_05200_),
    .A2(_05203_),
    .Y(_05205_),
    .B1(net1383));
 sg13g2_o21ai_1 _11176_ (.B1(_05205_),
    .Y(_05206_),
    .A1(_05200_),
    .A2(_05203_));
 sg13g2_nand2_1 _11177_ (.Y(_05207_),
    .A(net371),
    .B(net1335));
 sg13g2_a21oi_1 _11178_ (.A1(_05206_),
    .A2(net372),
    .Y(_00342_),
    .B1(net1735));
 sg13g2_a21o_2 _11179_ (.A2(_05203_),
    .A1(_05200_),
    .B1(_05201_),
    .X(_05208_));
 sg13g2_and2_1 _11180_ (.A(\mac_inst.accumulator[7] ),
    .B(_03153_),
    .X(_05209_));
 sg13g2_nand2_1 _11181_ (.Y(_05210_),
    .A(\mac_inst.accumulator[7] ),
    .B(_03154_));
 sg13g2_xor2_1 _11182_ (.B(_03153_),
    .A(\mac_inst.accumulator[7] ),
    .X(_05211_));
 sg13g2_a21oi_1 _11183_ (.A1(_05208_),
    .A2(_05211_),
    .Y(_05212_),
    .B1(net1383));
 sg13g2_o21ai_1 _11184_ (.B1(_05212_),
    .Y(_05213_),
    .A1(_05208_),
    .A2(_05211_));
 sg13g2_nand2_1 _11185_ (.Y(_05214_),
    .A(net377),
    .B(net1332));
 sg13g2_a21oi_1 _11186_ (.A1(_05213_),
    .A2(_05214_),
    .Y(_00343_),
    .B1(net1735));
 sg13g2_a21oi_2 _11187_ (.B1(_05209_),
    .Y(_05215_),
    .A2(_05211_),
    .A1(_05208_));
 sg13g2_and2_1 _11188_ (.A(\mac_inst.accumulator[8] ),
    .B(_03282_),
    .X(_05216_));
 sg13g2_xnor2_1 _11189_ (.Y(_05217_),
    .A(\mac_inst.accumulator[8] ),
    .B(_03282_));
 sg13g2_nand2_1 _11190_ (.Y(_05218_),
    .A(_05215_),
    .B(_05217_));
 sg13g2_nor2_1 _11191_ (.A(_05215_),
    .B(_05217_),
    .Y(_05219_));
 sg13g2_nand3b_1 _11192_ (.B(net1468),
    .C(_05218_),
    .Y(_05220_),
    .A_N(_05219_));
 sg13g2_nand2_1 _11193_ (.Y(_05221_),
    .A(net595),
    .B(net1330));
 sg13g2_a21oi_1 _11194_ (.A1(_05220_),
    .A2(_05221_),
    .Y(_00344_),
    .B1(net1734));
 sg13g2_nor2_1 _11195_ (.A(_05535_),
    .B(_03408_),
    .Y(_05222_));
 sg13g2_and2_1 _11196_ (.A(\mac_inst.accumulator[9] ),
    .B(_03408_),
    .X(_05223_));
 sg13g2_xnor2_1 _11197_ (.Y(_05224_),
    .A(_05535_),
    .B(_03408_));
 sg13g2_nor3_1 _11198_ (.A(_05216_),
    .B(_05219_),
    .C(net1201),
    .Y(_05225_));
 sg13g2_nand2_1 _11199_ (.Y(_05226_),
    .A(_05219_),
    .B(net1201));
 sg13g2_a21oi_1 _11200_ (.A1(_05216_),
    .A2(net1201),
    .Y(_05227_),
    .B1(_05225_));
 sg13g2_nand3_1 _11201_ (.B(_05226_),
    .C(_05227_),
    .A(net1468),
    .Y(_05228_));
 sg13g2_nand2_1 _11202_ (.Y(_05229_),
    .A(net586),
    .B(net1330));
 sg13g2_a21oi_1 _11203_ (.A1(_05228_),
    .A2(_05229_),
    .Y(_00345_),
    .B1(net1734));
 sg13g2_a21oi_1 _11204_ (.A1(_05216_),
    .A2(net1201),
    .Y(_05230_),
    .B1(_05223_));
 sg13g2_nand2_1 _11205_ (.Y(_05231_),
    .A(_05226_),
    .B(_05230_));
 sg13g2_nand2_1 _11206_ (.Y(_05232_),
    .A(\mac_inst.accumulator[10] ),
    .B(_03544_));
 sg13g2_nor2b_1 _11207_ (.A(_03544_),
    .B_N(\mac_inst.accumulator[10] ),
    .Y(_05233_));
 sg13g2_xor2_1 _11208_ (.B(_03544_),
    .A(\mac_inst.accumulator[10] ),
    .X(_05234_));
 sg13g2_inv_1 _11209_ (.Y(_05235_),
    .A(_05234_));
 sg13g2_a21oi_1 _11210_ (.A1(_05226_),
    .A2(_05230_),
    .Y(_05236_),
    .B1(_05234_));
 sg13g2_nor2_1 _11211_ (.A(net1383),
    .B(_05236_),
    .Y(_05237_));
 sg13g2_o21ai_1 _11212_ (.B1(_05237_),
    .Y(_05238_),
    .A1(_05231_),
    .A2(_05235_));
 sg13g2_nand2_1 _11213_ (.Y(_05239_),
    .A(net557),
    .B(net1331));
 sg13g2_a21oi_1 _11214_ (.A1(_05238_),
    .A2(_05239_),
    .Y(_00346_),
    .B1(net1734));
 sg13g2_nand2_1 _11215_ (.Y(_05240_),
    .A(_05534_),
    .B(_03673_));
 sg13g2_xnor2_1 _11216_ (.Y(_05241_),
    .A(\mac_inst.accumulator[11] ),
    .B(_03673_));
 sg13g2_nor2_1 _11217_ (.A(_05233_),
    .B(_05236_),
    .Y(_05242_));
 sg13g2_a21oi_1 _11218_ (.A1(_05241_),
    .A2(_05242_),
    .Y(_05243_),
    .B1(net1383));
 sg13g2_o21ai_1 _11219_ (.B1(_05243_),
    .Y(_05244_),
    .A1(_05241_),
    .A2(_05242_));
 sg13g2_nand2_1 _11220_ (.Y(_05245_),
    .A(net405),
    .B(net1333));
 sg13g2_a21oi_1 _11221_ (.A1(_05244_),
    .A2(_05245_),
    .Y(_00347_),
    .B1(net1735));
 sg13g2_nor2_1 _11222_ (.A(_05234_),
    .B(_05241_),
    .Y(_05246_));
 sg13g2_nand3b_1 _11223_ (.B(net1201),
    .C(_05246_),
    .Y(_05247_),
    .A_N(_05217_));
 sg13g2_or2_1 _11224_ (.X(_05248_),
    .B(_05247_),
    .A(_05215_));
 sg13g2_and2_1 _11225_ (.A(\mac_inst.accumulator[11] ),
    .B(_03673_),
    .X(_05249_));
 sg13g2_nor3_1 _11226_ (.A(_05230_),
    .B(_05234_),
    .C(_05241_),
    .Y(_05250_));
 sg13g2_nor2b_1 _11227_ (.A(_05241_),
    .B_N(_05233_),
    .Y(_05251_));
 sg13g2_or2_1 _11228_ (.X(_05252_),
    .B(_05251_),
    .A(_05250_));
 sg13g2_nor3_1 _11229_ (.A(_05249_),
    .B(_05250_),
    .C(_05251_),
    .Y(_05253_));
 sg13g2_o21ai_1 _11230_ (.B1(_05253_),
    .Y(_05254_),
    .A1(_05215_),
    .A2(_05247_));
 sg13g2_or2_1 _11231_ (.X(_05255_),
    .B(_03803_),
    .A(_05533_));
 sg13g2_and2_1 _11232_ (.A(net552),
    .B(_03803_),
    .X(_05256_));
 sg13g2_xnor2_1 _11233_ (.Y(_05257_),
    .A(_05533_),
    .B(_03803_));
 sg13g2_inv_1 _11234_ (.Y(_05258_),
    .A(_05257_));
 sg13g2_a21oi_1 _11235_ (.A1(_05254_),
    .A2(_05257_),
    .Y(_05259_),
    .B1(net1383));
 sg13g2_o21ai_1 _11236_ (.B1(_05259_),
    .Y(_05260_),
    .A1(_05254_),
    .A2(_05257_));
 sg13g2_nand2_1 _11237_ (.Y(_05261_),
    .A(net433),
    .B(net1333));
 sg13g2_a21oi_1 _11238_ (.A1(_05260_),
    .A2(_05261_),
    .Y(_00348_),
    .B1(net1738));
 sg13g2_nor2b_1 _11239_ (.A(\mac_inst.accumulator[13] ),
    .B_N(_03934_),
    .Y(_05262_));
 sg13g2_nor2b_2 _11240_ (.A(_03934_),
    .B_N(\mac_inst.accumulator[13] ),
    .Y(_05263_));
 sg13g2_xnor2_1 _11241_ (.Y(_05264_),
    .A(\mac_inst.accumulator[13] ),
    .B(_03934_));
 sg13g2_or2_1 _11242_ (.X(_05265_),
    .B(_05263_),
    .A(_05262_));
 sg13g2_a21oi_1 _11243_ (.A1(_05254_),
    .A2(_05257_),
    .Y(_05266_),
    .B1(_05256_));
 sg13g2_nor2_1 _11244_ (.A(_05265_),
    .B(_05266_),
    .Y(_05267_));
 sg13g2_a21oi_1 _11245_ (.A1(_05265_),
    .A2(_05266_),
    .Y(_05268_),
    .B1(net1383));
 sg13g2_nand2b_1 _11246_ (.Y(_05269_),
    .B(_05268_),
    .A_N(_05267_));
 sg13g2_nand2_1 _11247_ (.Y(_05270_),
    .A(net461),
    .B(net1333));
 sg13g2_a21oi_1 _11248_ (.A1(_05269_),
    .A2(_05270_),
    .Y(_00349_),
    .B1(net1742));
 sg13g2_nand2_1 _11249_ (.Y(_05271_),
    .A(\mac_inst.accumulator[14] ),
    .B(_04068_));
 sg13g2_nand2b_1 _11250_ (.Y(_05272_),
    .B(\mac_inst.accumulator[14] ),
    .A_N(_04068_));
 sg13g2_xor2_1 _11251_ (.B(_04068_),
    .A(\mac_inst.accumulator[14] ),
    .X(_05273_));
 sg13g2_inv_1 _11252_ (.Y(_05274_),
    .A(_05273_));
 sg13g2_or3_1 _11253_ (.A(_05263_),
    .B(_05267_),
    .C(_05274_),
    .X(_05275_));
 sg13g2_o21ai_1 _11254_ (.B1(_05274_),
    .Y(_05276_),
    .A1(_05263_),
    .A2(_05267_));
 sg13g2_nand3_1 _11255_ (.B(_05275_),
    .C(_05276_),
    .A(net1468),
    .Y(_05277_));
 sg13g2_nand2_1 _11256_ (.Y(_05278_),
    .A(net534),
    .B(net1333));
 sg13g2_a21oi_1 _11257_ (.A1(_05277_),
    .A2(_05278_),
    .Y(_00350_),
    .B1(net1738));
 sg13g2_nor2_1 _11258_ (.A(\mac_inst.accumulator[15] ),
    .B(_04200_),
    .Y(_05279_));
 sg13g2_xor2_1 _11259_ (.B(_04200_),
    .A(\mac_inst.accumulator[15] ),
    .X(_05280_));
 sg13g2_and2_1 _11260_ (.A(_05272_),
    .B(_05276_),
    .X(_05281_));
 sg13g2_o21ai_1 _11261_ (.B1(net1466),
    .Y(_05282_),
    .A1(net1200),
    .A2(_05281_));
 sg13g2_a21oi_1 _11262_ (.A1(net1200),
    .A2(_05281_),
    .Y(_05283_),
    .B1(_05282_));
 sg13g2_a21oi_1 _11263_ (.A1(net573),
    .A2(net1336),
    .Y(_05284_),
    .B1(_05283_));
 sg13g2_nor2_1 _11264_ (.A(net1738),
    .B(_05284_),
    .Y(_00351_));
 sg13g2_nor2_1 _11265_ (.A(_05256_),
    .B(_05263_),
    .Y(_05285_));
 sg13g2_nor4_1 _11266_ (.A(_05262_),
    .B(_05273_),
    .C(net1200),
    .D(_05285_),
    .Y(_05286_));
 sg13g2_nand2b_1 _11267_ (.Y(_05287_),
    .B(\mac_inst.accumulator[15] ),
    .A_N(_04200_));
 sg13g2_o21ai_1 _11268_ (.B1(_05287_),
    .Y(_05288_),
    .A1(_05272_),
    .A2(net1200));
 sg13g2_nor4_1 _11269_ (.A(_05249_),
    .B(_05252_),
    .C(_05286_),
    .D(_05288_),
    .Y(_05289_));
 sg13g2_nor4_1 _11270_ (.A(_05258_),
    .B(_05265_),
    .C(_05273_),
    .D(net1200),
    .Y(_05290_));
 sg13g2_nor3_1 _11271_ (.A(_05286_),
    .B(_05288_),
    .C(_05290_),
    .Y(_05291_));
 sg13g2_a21o_2 _11272_ (.A2(_05289_),
    .A1(_05248_),
    .B1(_05291_),
    .X(_05292_));
 sg13g2_nand2_1 _11273_ (.Y(_05293_),
    .A(\mac_inst.accumulator[16] ),
    .B(_04331_));
 sg13g2_and2_1 _11274_ (.A(\mac_inst.accumulator[16] ),
    .B(_04330_),
    .X(_05294_));
 sg13g2_xor2_1 _11275_ (.B(_04330_),
    .A(\mac_inst.accumulator[16] ),
    .X(_05295_));
 sg13g2_nand2b_1 _11276_ (.Y(_05296_),
    .B(_05292_),
    .A_N(_05295_));
 sg13g2_nand2b_1 _11277_ (.Y(_05297_),
    .B(_05295_),
    .A_N(_05292_));
 sg13g2_and3_1 _11278_ (.X(_05298_),
    .A(net1466),
    .B(_05296_),
    .C(_05297_));
 sg13g2_a21oi_1 _11279_ (.A1(net592),
    .A2(net1336),
    .Y(_05299_),
    .B1(_05298_));
 sg13g2_nor2_1 _11280_ (.A(net1738),
    .B(_05299_),
    .Y(_00352_));
 sg13g2_and2_1 _11281_ (.A(\mac_inst.accumulator[17] ),
    .B(_04457_),
    .X(_05300_));
 sg13g2_inv_1 _11282_ (.Y(_05301_),
    .A(_05300_));
 sg13g2_nor2b_1 _11283_ (.A(_04457_),
    .B_N(\mac_inst.accumulator[17] ),
    .Y(_05302_));
 sg13g2_xnor2_1 _11284_ (.Y(_05303_),
    .A(\mac_inst.accumulator[17] ),
    .B(_04457_));
 sg13g2_nor2_1 _11285_ (.A(_05294_),
    .B(_05303_),
    .Y(_05304_));
 sg13g2_nand2_1 _11286_ (.Y(_05305_),
    .A(_05297_),
    .B(_05304_));
 sg13g2_nand2_1 _11287_ (.Y(_05306_),
    .A(_05295_),
    .B(_05303_));
 sg13g2_nor2_1 _11288_ (.A(_05292_),
    .B(_05306_),
    .Y(_05307_));
 sg13g2_or2_1 _11289_ (.X(_05308_),
    .B(_05306_),
    .A(_05292_));
 sg13g2_a21oi_1 _11290_ (.A1(_05294_),
    .A2(_05303_),
    .Y(_05309_),
    .B1(net1384));
 sg13g2_nand3_1 _11291_ (.B(_05308_),
    .C(_05309_),
    .A(_05305_),
    .Y(_05310_));
 sg13g2_nand2_1 _11292_ (.Y(_05311_),
    .A(net496),
    .B(net1336));
 sg13g2_a21oi_1 _11293_ (.A1(_05310_),
    .A2(_05311_),
    .Y(_00353_),
    .B1(net1740));
 sg13g2_nor2_2 _11294_ (.A(_05532_),
    .B(_04581_),
    .Y(_05312_));
 sg13g2_and2_1 _11295_ (.A(_05532_),
    .B(_04581_),
    .X(_05313_));
 sg13g2_nor2_1 _11296_ (.A(_05312_),
    .B(_05313_),
    .Y(_05314_));
 sg13g2_or2_1 _11297_ (.X(_05315_),
    .B(_05313_),
    .A(_05312_));
 sg13g2_a21oi_1 _11298_ (.A1(_05294_),
    .A2(_05303_),
    .Y(_05316_),
    .B1(_05302_));
 sg13g2_nand3_1 _11299_ (.B(_05314_),
    .C(_05316_),
    .A(_05308_),
    .Y(_05317_));
 sg13g2_a21oi_1 _11300_ (.A1(_05308_),
    .A2(_05316_),
    .Y(_05318_),
    .B1(_05314_));
 sg13g2_nand3b_1 _11301_ (.B(net1467),
    .C(_05317_),
    .Y(_05319_),
    .A_N(_05318_));
 sg13g2_nand2_1 _11302_ (.Y(_05320_),
    .A(net506),
    .B(net1338));
 sg13g2_a21oi_1 _11303_ (.A1(_05319_),
    .A2(_05320_),
    .Y(_00354_),
    .B1(net1741));
 sg13g2_nand2b_1 _11304_ (.Y(_05321_),
    .B(\mac_inst.accumulator[19] ),
    .A_N(_04711_));
 sg13g2_nor2b_1 _11305_ (.A(\mac_inst.accumulator[19] ),
    .B_N(_04711_),
    .Y(_05322_));
 sg13g2_xnor2_1 _11306_ (.Y(_05323_),
    .A(\mac_inst.accumulator[19] ),
    .B(_04711_));
 sg13g2_inv_1 _11307_ (.Y(_05324_),
    .A(_05323_));
 sg13g2_nand2_1 _11308_ (.Y(_05325_),
    .A(\mac_inst.accumulator[18] ),
    .B(_04581_));
 sg13g2_nand2b_1 _11309_ (.Y(_05326_),
    .B(_05325_),
    .A_N(_05318_));
 sg13g2_a21oi_1 _11310_ (.A1(_05323_),
    .A2(_05326_),
    .Y(_05327_),
    .B1(net1384));
 sg13g2_o21ai_1 _11311_ (.B1(_05327_),
    .Y(_05328_),
    .A1(_05323_),
    .A2(_05326_));
 sg13g2_nand2_1 _11312_ (.Y(_05329_),
    .A(net548),
    .B(net1336));
 sg13g2_a21oi_1 _11313_ (.A1(_05328_),
    .A2(_05329_),
    .Y(_00355_),
    .B1(net1742));
 sg13g2_and2_1 _11314_ (.A(_05321_),
    .B(_05325_),
    .X(_05330_));
 sg13g2_o21ai_1 _11315_ (.B1(_05316_),
    .Y(_05331_),
    .A1(_05322_),
    .A2(_05330_));
 sg13g2_a21oi_1 _11316_ (.A1(_05314_),
    .A2(_05330_),
    .Y(_05332_),
    .B1(_05322_));
 sg13g2_o21ai_1 _11317_ (.B1(_05332_),
    .Y(_05333_),
    .A1(_05307_),
    .A2(_05331_));
 sg13g2_nand2_1 _11318_ (.Y(_05334_),
    .A(\mac_inst.accumulator[20] ),
    .B(_04835_));
 sg13g2_nor2b_1 _11319_ (.A(_04835_),
    .B_N(\mac_inst.accumulator[20] ),
    .Y(_05335_));
 sg13g2_xnor2_1 _11320_ (.Y(_05336_),
    .A(\mac_inst.accumulator[20] ),
    .B(_04835_));
 sg13g2_nor2b_1 _11321_ (.A(_05336_),
    .B_N(_05333_),
    .Y(_05337_));
 sg13g2_nand2b_1 _11322_ (.Y(_05338_),
    .B(_05336_),
    .A_N(_05333_));
 sg13g2_nand3b_1 _11323_ (.B(_05338_),
    .C(net1467),
    .Y(_05339_),
    .A_N(_05337_));
 sg13g2_nand2_1 _11324_ (.Y(_05340_),
    .A(net553),
    .B(net1338));
 sg13g2_a21oi_1 _11325_ (.A1(_05339_),
    .A2(_05340_),
    .Y(_00356_),
    .B1(net1740));
 sg13g2_nor2_1 _11326_ (.A(_05531_),
    .B(_04955_),
    .Y(_05341_));
 sg13g2_nand2_1 _11327_ (.Y(_05342_),
    .A(\mac_inst.accumulator[21] ),
    .B(_04955_));
 sg13g2_xnor2_1 _11328_ (.Y(_05343_),
    .A(\mac_inst.accumulator[21] ),
    .B(_04955_));
 sg13g2_nor2_1 _11329_ (.A(_05335_),
    .B(_05343_),
    .Y(_05344_));
 sg13g2_nand2_1 _11330_ (.Y(_05345_),
    .A(_05338_),
    .B(_05344_));
 sg13g2_nand3b_1 _11331_ (.B(_05336_),
    .C(_05343_),
    .Y(_05346_),
    .A_N(_05333_));
 sg13g2_a21oi_1 _11332_ (.A1(_05335_),
    .A2(_05343_),
    .Y(_05347_),
    .B1(net1384));
 sg13g2_nand3_1 _11333_ (.B(_05346_),
    .C(_05347_),
    .A(_05345_),
    .Y(_05348_));
 sg13g2_nand2_1 _11334_ (.Y(_05349_),
    .A(net510),
    .B(net1339));
 sg13g2_a21oi_1 _11335_ (.A1(_05348_),
    .A2(_05349_),
    .Y(_00357_),
    .B1(net1740));
 sg13g2_a21oi_1 _11336_ (.A1(_05335_),
    .A2(_05343_),
    .Y(_05350_),
    .B1(_05341_));
 sg13g2_nor2b_1 _11337_ (.A(_05074_),
    .B_N(\mac_inst.accumulator[22] ),
    .Y(_05351_));
 sg13g2_nand2_1 _11338_ (.Y(_05352_),
    .A(\mac_inst.accumulator[22] ),
    .B(_05074_));
 sg13g2_xor2_1 _11339_ (.B(_05074_),
    .A(\mac_inst.accumulator[22] ),
    .X(_05353_));
 sg13g2_nand3_1 _11340_ (.B(_05350_),
    .C(_05353_),
    .A(_05346_),
    .Y(_05354_));
 sg13g2_a21oi_1 _11341_ (.A1(_05346_),
    .A2(_05350_),
    .Y(_05355_),
    .B1(_05353_));
 sg13g2_nand3b_1 _11342_ (.B(net1467),
    .C(_05354_),
    .Y(_05356_),
    .A_N(_05355_));
 sg13g2_nand2_1 _11343_ (.Y(_05357_),
    .A(net448),
    .B(net1338));
 sg13g2_a21oi_1 _11344_ (.A1(_05356_),
    .A2(_05357_),
    .Y(_00358_),
    .B1(net1741));
 sg13g2_xor2_1 _11345_ (.B(_05154_),
    .A(\mac_inst.accumulator[23] ),
    .X(_05358_));
 sg13g2_or3_1 _11346_ (.A(_05351_),
    .B(_05355_),
    .C(_05358_),
    .X(_05359_));
 sg13g2_o21ai_1 _11347_ (.B1(_05358_),
    .Y(_05360_),
    .A1(_05351_),
    .A2(_05355_));
 sg13g2_nand3_1 _11348_ (.B(_05359_),
    .C(_05360_),
    .A(net1467),
    .Y(_05361_));
 sg13g2_nand2_1 _11349_ (.Y(_05362_),
    .A(net406),
    .B(net1340));
 sg13g2_a21oi_1 _11350_ (.A1(_05361_),
    .A2(net407),
    .Y(_00359_),
    .B1(net1742));
 sg13g2_nor2b_2 _11351_ (.A(net1466),
    .B_N(mac_en_mac),
    .Y(_05363_));
 sg13g2_nand2_2 _11352_ (.Y(_05364_),
    .A(net1383),
    .B(mac_en_mac));
 sg13g2_a22oi_1 _11353_ (.Y(_05365_),
    .B1(net1329),
    .B2(_05157_),
    .A2(net1337),
    .A1(net598));
 sg13g2_nor2_1 _11354_ (.A(net1741),
    .B(net599),
    .Y(_00360_));
 sg13g2_o21ai_1 _11355_ (.B1(net1329),
    .Y(_05366_),
    .A1(_05156_),
    .A2(_05165_));
 sg13g2_a21oi_1 _11356_ (.A1(_05156_),
    .A2(_05165_),
    .Y(_05367_),
    .B1(_05366_));
 sg13g2_a21oi_1 _11357_ (.A1(net538),
    .A2(net1340),
    .Y(_05368_),
    .B1(_05367_));
 sg13g2_nor2_1 _11358_ (.A(net1744),
    .B(net539),
    .Y(_00361_));
 sg13g2_o21ai_1 _11359_ (.B1(_05162_),
    .Y(_05369_),
    .A1(_05156_),
    .A2(_05165_));
 sg13g2_o21ai_1 _11360_ (.B1(net1328),
    .Y(_05370_),
    .A1(_05173_),
    .A2(_05369_));
 sg13g2_a21oi_1 _11361_ (.A1(_05173_),
    .A2(_05369_),
    .Y(_05371_),
    .B1(_05370_));
 sg13g2_a21oi_1 _11362_ (.A1(net543),
    .A2(net1337),
    .Y(_05372_),
    .B1(_05371_));
 sg13g2_nor2_1 _11363_ (.A(net1743),
    .B(net544),
    .Y(_00362_));
 sg13g2_a21o_1 _11364_ (.A2(_05369_),
    .A1(_05173_),
    .B1(_05171_),
    .X(_05373_));
 sg13g2_a21oi_1 _11365_ (.A1(_05180_),
    .A2(_05373_),
    .Y(_05374_),
    .B1(net1319));
 sg13g2_o21ai_1 _11366_ (.B1(_05374_),
    .Y(_05375_),
    .A1(_05180_),
    .A2(_05373_));
 sg13g2_nand2_1 _11367_ (.Y(_05376_),
    .A(net369),
    .B(net1334));
 sg13g2_a21oi_1 _11368_ (.A1(_05375_),
    .A2(_05376_),
    .Y(_00363_),
    .B1(net1743));
 sg13g2_a21o_1 _11369_ (.A2(_05373_),
    .A1(_05180_),
    .B1(_05178_),
    .X(_05377_));
 sg13g2_a21oi_1 _11370_ (.A1(_05188_),
    .A2(_05377_),
    .Y(_05378_),
    .B1(net1319));
 sg13g2_o21ai_1 _11371_ (.B1(_05378_),
    .Y(_05379_),
    .A1(_05188_),
    .A2(_05377_));
 sg13g2_nand2_1 _11372_ (.Y(_05380_),
    .A(net515),
    .B(net1334));
 sg13g2_a21oi_1 _11373_ (.A1(_05379_),
    .A2(_05380_),
    .Y(_00364_),
    .B1(net1737));
 sg13g2_a21oi_1 _11374_ (.A1(_05188_),
    .A2(_05377_),
    .Y(_05381_),
    .B1(_05185_));
 sg13g2_a21oi_1 _11375_ (.A1(_05196_),
    .A2(_05381_),
    .Y(_05382_),
    .B1(net1319));
 sg13g2_o21ai_1 _11376_ (.B1(_05382_),
    .Y(_05383_),
    .A1(_05196_),
    .A2(_05381_));
 sg13g2_nand2_1 _11377_ (.Y(_05384_),
    .A(net378),
    .B(net1332));
 sg13g2_a21oi_1 _11378_ (.A1(_05383_),
    .A2(_05384_),
    .Y(_00365_),
    .B1(net1737));
 sg13g2_o21ai_1 _11379_ (.B1(_05193_),
    .Y(_05385_),
    .A1(_05196_),
    .A2(_05381_));
 sg13g2_a21oi_1 _11380_ (.A1(_05204_),
    .A2(_05385_),
    .Y(_05386_),
    .B1(net1319));
 sg13g2_o21ai_1 _11381_ (.B1(_05386_),
    .Y(_05387_),
    .A1(_05204_),
    .A2(_05385_));
 sg13g2_nand2_1 _11382_ (.Y(_05388_),
    .A(net537),
    .B(net1331));
 sg13g2_a21oi_1 _11383_ (.A1(_05387_),
    .A2(_05388_),
    .Y(_00366_),
    .B1(net1735));
 sg13g2_a21oi_1 _11384_ (.A1(_05204_),
    .A2(_05385_),
    .Y(_05389_),
    .B1(_05202_));
 sg13g2_a21oi_1 _11385_ (.A1(_05211_),
    .A2(_05389_),
    .Y(_05390_),
    .B1(net1319));
 sg13g2_o21ai_1 _11386_ (.B1(_05390_),
    .Y(_05391_),
    .A1(_05211_),
    .A2(_05389_));
 sg13g2_nand2_1 _11387_ (.Y(_05392_),
    .A(net550),
    .B(net1331));
 sg13g2_a21oi_1 _11388_ (.A1(_05391_),
    .A2(_05392_),
    .Y(_00367_),
    .B1(net1735));
 sg13g2_o21ai_1 _11389_ (.B1(_05210_),
    .Y(_05393_),
    .A1(_05211_),
    .A2(_05389_));
 sg13g2_or2_1 _11390_ (.X(_05394_),
    .B(_05393_),
    .A(_05217_));
 sg13g2_nand2_1 _11391_ (.Y(_05395_),
    .A(_05217_),
    .B(_05393_));
 sg13g2_nand3_1 _11392_ (.B(_05394_),
    .C(_05395_),
    .A(net1328),
    .Y(_05396_));
 sg13g2_nand2_1 _11393_ (.Y(_05397_),
    .A(net560),
    .B(net1330));
 sg13g2_a21oi_1 _11394_ (.A1(_05396_),
    .A2(_05397_),
    .Y(_00368_),
    .B1(net1734));
 sg13g2_nand2_1 _11395_ (.Y(_05398_),
    .A(\mac_inst.accumulator[8] ),
    .B(_03283_));
 sg13g2_nand3_1 _11396_ (.B(_05395_),
    .C(_05398_),
    .A(net1201),
    .Y(_05399_));
 sg13g2_nor2_1 _11397_ (.A(net1201),
    .B(_05398_),
    .Y(_05400_));
 sg13g2_nor2_1 _11398_ (.A(net1201),
    .B(_05395_),
    .Y(_05401_));
 sg13g2_nor3_1 _11399_ (.A(net1319),
    .B(_05400_),
    .C(_05401_),
    .Y(_05402_));
 sg13g2_nand2_1 _11400_ (.Y(_05403_),
    .A(_05399_),
    .B(_05402_));
 sg13g2_nand2_1 _11401_ (.Y(_05404_),
    .A(net561),
    .B(net1330));
 sg13g2_a21oi_1 _11402_ (.A1(_05403_),
    .A2(_05404_),
    .Y(_00369_),
    .B1(net1734));
 sg13g2_or2_1 _11403_ (.X(_05405_),
    .B(_05400_),
    .A(_05222_));
 sg13g2_or2_1 _11404_ (.X(_05406_),
    .B(_05405_),
    .A(_05401_));
 sg13g2_nand2b_1 _11405_ (.Y(_05407_),
    .B(_05235_),
    .A_N(_05406_));
 sg13g2_nand2_1 _11406_ (.Y(_05408_),
    .A(_05234_),
    .B(_05406_));
 sg13g2_nand3_1 _11407_ (.B(_05407_),
    .C(_05408_),
    .A(net1328),
    .Y(_05409_));
 sg13g2_nand2_1 _11408_ (.Y(_05410_),
    .A(net588),
    .B(net1330));
 sg13g2_a21oi_1 _11409_ (.A1(_05409_),
    .A2(_05410_),
    .Y(_00370_),
    .B1(net1734));
 sg13g2_nand2_1 _11410_ (.Y(_05411_),
    .A(_05232_),
    .B(_05408_));
 sg13g2_xor2_1 _11411_ (.B(_05411_),
    .A(_05241_),
    .X(_05412_));
 sg13g2_nand2_1 _11412_ (.Y(_05413_),
    .A(net1328),
    .B(_05412_));
 sg13g2_nand2_1 _11413_ (.Y(_05414_),
    .A(net607),
    .B(net1331));
 sg13g2_a21oi_1 _11414_ (.A1(_05413_),
    .A2(_05414_),
    .Y(_00371_),
    .B1(net1734));
 sg13g2_and2_1 _11415_ (.A(_05234_),
    .B(_05241_),
    .X(_05415_));
 sg13g2_nor2b_1 _11416_ (.A(_05224_),
    .B_N(_05217_),
    .Y(_05416_));
 sg13g2_nand3_1 _11417_ (.B(_05415_),
    .C(_05416_),
    .A(_05393_),
    .Y(_05417_));
 sg13g2_o21ai_1 _11418_ (.B1(_05232_),
    .Y(_05418_),
    .A1(_05534_),
    .A2(_03673_));
 sg13g2_a22oi_1 _11419_ (.Y(_05419_),
    .B1(_05418_),
    .B2(_05240_),
    .A2(_05415_),
    .A1(_05405_));
 sg13g2_a21oi_1 _11420_ (.A1(_05417_),
    .A2(_05419_),
    .Y(_05420_),
    .B1(_05257_));
 sg13g2_nand3_1 _11421_ (.B(_05417_),
    .C(_05419_),
    .A(_05257_),
    .Y(_05421_));
 sg13g2_nand3b_1 _11422_ (.B(_05421_),
    .C(net1328),
    .Y(_05422_),
    .A_N(_05420_));
 sg13g2_nand2_1 _11423_ (.Y(_05423_),
    .A(net563),
    .B(net1333));
 sg13g2_a21oi_1 _11424_ (.A1(_05422_),
    .A2(_05423_),
    .Y(_00372_),
    .B1(net1738));
 sg13g2_and2_1 _11425_ (.A(_05265_),
    .B(_05420_),
    .X(_05424_));
 sg13g2_nand2_1 _11426_ (.Y(_05425_),
    .A(_05255_),
    .B(_05264_));
 sg13g2_nor2_1 _11427_ (.A(_05420_),
    .B(_05425_),
    .Y(_05426_));
 sg13g2_o21ai_1 _11428_ (.B1(net1328),
    .Y(_05427_),
    .A1(_05255_),
    .A2(_05264_));
 sg13g2_nor3_1 _11429_ (.A(_05424_),
    .B(_05426_),
    .C(_05427_),
    .Y(_05428_));
 sg13g2_a21oi_1 _11430_ (.A1(net602),
    .A2(net1333),
    .Y(_05429_),
    .B1(_05428_));
 sg13g2_nor2_1 _11431_ (.A(net1739),
    .B(_05429_),
    .Y(_00373_));
 sg13g2_nand2_1 _11432_ (.Y(_05430_),
    .A(\mac_inst.accumulator[13] ),
    .B(_03934_));
 sg13g2_o21ai_1 _11433_ (.B1(_05430_),
    .Y(_05431_),
    .A1(_05255_),
    .A2(_05264_));
 sg13g2_or2_1 _11434_ (.X(_05432_),
    .B(_05431_),
    .A(_05424_));
 sg13g2_nand2_1 _11435_ (.Y(_05433_),
    .A(_05273_),
    .B(_05432_));
 sg13g2_o21ai_1 _11436_ (.B1(net1328),
    .Y(_05434_),
    .A1(_05273_),
    .A2(_05432_));
 sg13g2_nand2b_1 _11437_ (.Y(_05435_),
    .B(_05433_),
    .A_N(_05434_));
 sg13g2_nand2_1 _11438_ (.Y(_05436_),
    .A(net570),
    .B(net1334));
 sg13g2_a21oi_1 _11439_ (.A1(_05435_),
    .A2(_05436_),
    .Y(_00374_),
    .B1(net1739));
 sg13g2_nand2_1 _11440_ (.Y(_05437_),
    .A(_05271_),
    .B(_05433_));
 sg13g2_a21oi_1 _11441_ (.A1(net1200),
    .A2(_05437_),
    .Y(_05438_),
    .B1(net1319));
 sg13g2_o21ai_1 _11442_ (.B1(_05438_),
    .Y(_05439_),
    .A1(_05280_),
    .A2(_05437_));
 sg13g2_nand2_1 _11443_ (.Y(_05440_),
    .A(net589),
    .B(net1337));
 sg13g2_a21oi_1 _11444_ (.A1(_05439_),
    .A2(net590),
    .Y(_00375_),
    .B1(net1739));
 sg13g2_nand3_1 _11445_ (.B(net1200),
    .C(_05431_),
    .A(_05273_),
    .Y(_05441_));
 sg13g2_a22oi_1 _11446_ (.Y(_05442_),
    .B1(_04200_),
    .B2(\mac_inst.accumulator[15] ),
    .A2(_04068_),
    .A1(\mac_inst.accumulator[14] ));
 sg13g2_or2_1 _11447_ (.X(_05443_),
    .B(_05442_),
    .A(_05279_));
 sg13g2_and2_1 _11448_ (.A(_05441_),
    .B(_05443_),
    .X(_05444_));
 sg13g2_nand4_1 _11449_ (.B(_05265_),
    .C(_05273_),
    .A(_05258_),
    .Y(_05445_),
    .D(net1200));
 sg13g2_and3_1 _11450_ (.X(_05446_),
    .A(_05419_),
    .B(_05441_),
    .C(_05443_));
 sg13g2_a22oi_1 _11451_ (.Y(_05447_),
    .B1(_05446_),
    .B2(_05417_),
    .A2(_05445_),
    .A1(_05444_));
 sg13g2_inv_1 _11452_ (.Y(_05448_),
    .A(_05447_));
 sg13g2_nand2_1 _11453_ (.Y(_05449_),
    .A(_05295_),
    .B(_05448_));
 sg13g2_nand2b_1 _11454_ (.Y(_05450_),
    .B(_05447_),
    .A_N(_05295_));
 sg13g2_nand3_1 _11455_ (.B(_05449_),
    .C(_05450_),
    .A(net1329),
    .Y(_05451_));
 sg13g2_nand2_1 _11456_ (.Y(_05452_),
    .A(net581),
    .B(net1336));
 sg13g2_a21oi_1 _11457_ (.A1(_05451_),
    .A2(_05452_),
    .Y(_00376_),
    .B1(net1738));
 sg13g2_a21o_1 _11458_ (.A2(_05450_),
    .A1(_05293_),
    .B1(_05303_),
    .X(_05453_));
 sg13g2_nand3_1 _11459_ (.B(_05303_),
    .C(_05450_),
    .A(_05293_),
    .Y(_05454_));
 sg13g2_nand3_1 _11460_ (.B(_05453_),
    .C(_05454_),
    .A(net1329),
    .Y(_05455_));
 sg13g2_nand2_1 _11461_ (.Y(_05456_),
    .A(net600),
    .B(net1336));
 sg13g2_a21oi_1 _11462_ (.A1(_05455_),
    .A2(_05456_),
    .Y(_00377_),
    .B1(net1740));
 sg13g2_nand3_1 _11463_ (.B(_05315_),
    .C(_05453_),
    .A(_05301_),
    .Y(_05457_));
 sg13g2_a21oi_1 _11464_ (.A1(_05301_),
    .A2(_05453_),
    .Y(_05458_),
    .B1(_05315_));
 sg13g2_nand3b_1 _11465_ (.B(net1329),
    .C(_05457_),
    .Y(_05459_),
    .A_N(_05458_));
 sg13g2_nand2_1 _11466_ (.Y(_05460_),
    .A(net558),
    .B(net1337));
 sg13g2_a21oi_1 _11467_ (.A1(_05459_),
    .A2(net559),
    .Y(_00378_),
    .B1(net1740));
 sg13g2_nor3_1 _11468_ (.A(_05312_),
    .B(_05324_),
    .C(_05458_),
    .Y(_05461_));
 sg13g2_o21ai_1 _11469_ (.B1(_05324_),
    .Y(_05462_),
    .A1(_05312_),
    .A2(_05458_));
 sg13g2_nor2_1 _11470_ (.A(net1319),
    .B(_05461_),
    .Y(_05463_));
 sg13g2_a21oi_1 _11471_ (.A1(_05462_),
    .A2(_05463_),
    .Y(_05464_),
    .B1(net1339));
 sg13g2_o21ai_1 _11472_ (.B1(net1757),
    .Y(_05465_),
    .A1(net643),
    .A2(_05159_));
 sg13g2_nor2_1 _11473_ (.A(_05464_),
    .B(_05465_),
    .Y(_00379_));
 sg13g2_nor4_1 _11474_ (.A(_05295_),
    .B(_05303_),
    .C(_05315_),
    .D(_05323_),
    .Y(_05466_));
 sg13g2_nor2_1 _11475_ (.A(_05300_),
    .B(_05312_),
    .Y(_05467_));
 sg13g2_or2_1 _11476_ (.X(_05468_),
    .B(_05303_),
    .A(_05293_));
 sg13g2_a221oi_1 _11477_ (.B2(_05468_),
    .C1(_05323_),
    .B1(_05467_),
    .A1(_05532_),
    .Y(_05469_),
    .A2(_04581_));
 sg13g2_a221oi_1 _11478_ (.B2(_05466_),
    .C1(_05469_),
    .B1(_05447_),
    .A1(\mac_inst.accumulator[19] ),
    .Y(_05470_),
    .A2(_04711_));
 sg13g2_a21oi_1 _11479_ (.A1(_05336_),
    .A2(_05470_),
    .Y(_05471_),
    .B1(_05364_));
 sg13g2_o21ai_1 _11480_ (.B1(_05471_),
    .Y(_05472_),
    .A1(_05336_),
    .A2(_05470_));
 sg13g2_nand2_1 _11481_ (.Y(_05473_),
    .A(net593),
    .B(net1338));
 sg13g2_a21oi_1 _11482_ (.A1(_05472_),
    .A2(_05473_),
    .Y(_00380_),
    .B1(net1741));
 sg13g2_o21ai_1 _11483_ (.B1(_05343_),
    .Y(_05474_),
    .A1(_05336_),
    .A2(_05470_));
 sg13g2_nand2b_1 _11484_ (.Y(_05475_),
    .B(_05334_),
    .A_N(_05474_));
 sg13g2_nor3_1 _11485_ (.A(_05336_),
    .B(_05343_),
    .C(_05470_),
    .Y(_05476_));
 sg13g2_o21ai_1 _11486_ (.B1(net1329),
    .Y(_05477_),
    .A1(_05334_),
    .A2(_05343_));
 sg13g2_nor2_1 _11487_ (.A(_05476_),
    .B(_05477_),
    .Y(_05478_));
 sg13g2_a21oi_1 _11488_ (.A1(_05475_),
    .A2(_05478_),
    .Y(_05479_),
    .B1(net1338));
 sg13g2_o21ai_1 _11489_ (.B1(net1759),
    .Y(_05480_),
    .A1(net639),
    .A2(_05159_));
 sg13g2_nor2_1 _11490_ (.A(_05479_),
    .B(_05480_),
    .Y(_00381_));
 sg13g2_o21ai_1 _11491_ (.B1(_05342_),
    .Y(_05481_),
    .A1(_05334_),
    .A2(_05343_));
 sg13g2_nor3_1 _11492_ (.A(_05353_),
    .B(_05476_),
    .C(_05481_),
    .Y(_05482_));
 sg13g2_o21ai_1 _11493_ (.B1(_05353_),
    .Y(_05483_),
    .A1(_05476_),
    .A2(_05481_));
 sg13g2_nand2_1 _11494_ (.Y(_05484_),
    .A(net1329),
    .B(_05483_));
 sg13g2_nor2_1 _11495_ (.A(_05482_),
    .B(_05484_),
    .Y(_05485_));
 sg13g2_a21oi_1 _11496_ (.A1(net551),
    .A2(net1339),
    .Y(_05486_),
    .B1(_05485_));
 sg13g2_nor2_1 _11497_ (.A(net1742),
    .B(_05486_),
    .Y(_00382_));
 sg13g2_nand3_1 _11498_ (.B(_05358_),
    .C(_05483_),
    .A(_05352_),
    .Y(_05487_));
 sg13g2_a21oi_1 _11499_ (.A1(_05352_),
    .A2(_05483_),
    .Y(_05488_),
    .B1(_05358_));
 sg13g2_nor2_1 _11500_ (.A(_05364_),
    .B(_05488_),
    .Y(_05489_));
 sg13g2_a21oi_1 _11501_ (.A1(_05487_),
    .A2(_05489_),
    .Y(_05490_),
    .B1(net1338));
 sg13g2_o21ai_1 _11502_ (.B1(net1760),
    .Y(_05491_),
    .A1(net666),
    .A2(_05159_));
 sg13g2_nor2_1 _11503_ (.A(_05490_),
    .B(_05491_),
    .Y(_00383_));
 sg13g2_o21ai_1 _11504_ (.B1(net1769),
    .Y(_05492_),
    .A1(\mac_inst.RDY_get_multiply ),
    .A2(net1473));
 sg13g2_nor2_1 _11505_ (.A(net278),
    .B(_05492_),
    .Y(_00384_));
 sg13g2_o21ai_1 _11506_ (.B1(net1776),
    .Y(_05493_),
    .A1(\mac_inst.RDY_get_msu ),
    .A2(mac_en_msu));
 sg13g2_nor2_1 _11507_ (.A(net274),
    .B(_05493_),
    .Y(_00385_));
 sg13g2_o21ai_1 _11508_ (.B1(net1769),
    .Y(_05494_),
    .A1(\mac_inst.RDY_get_mac ),
    .A2(mac_en_mac));
 sg13g2_nor2_1 _11509_ (.A(net276),
    .B(_05494_),
    .Y(_00386_));
 sg13g2_o21ai_1 _11510_ (.B1(_05157_),
    .Y(_05495_),
    .A1(net1466),
    .A2(mac_en_mac));
 sg13g2_o21ai_1 _11511_ (.B1(net1758),
    .Y(_05496_),
    .A1(net733),
    .A2(_05159_));
 sg13g2_a21oi_1 _11512_ (.A1(_05159_),
    .A2(_05495_),
    .Y(_00387_),
    .B1(_05496_));
 sg13g2_a21oi_1 _11513_ (.A1(net735),
    .A2(net1340),
    .Y(_05497_),
    .B1(_05367_));
 sg13g2_a21oi_1 _11514_ (.A1(_05167_),
    .A2(net736),
    .Y(_00388_),
    .B1(net1741));
 sg13g2_a21oi_1 _11515_ (.A1(net726),
    .A2(net1337),
    .Y(_05498_),
    .B1(_05371_));
 sg13g2_a21oi_1 _11516_ (.A1(_05175_),
    .A2(net727),
    .Y(_00389_),
    .B1(net1739));
 sg13g2_nand2_1 _11517_ (.Y(_05499_),
    .A(net830),
    .B(net1334));
 sg13g2_nand3_1 _11518_ (.B(_05375_),
    .C(_05499_),
    .A(_05182_),
    .Y(_05500_));
 sg13g2_and2_1 _11519_ (.A(net1752),
    .B(_05500_),
    .X(_00390_));
 sg13g2_nand2_1 _11520_ (.Y(_05501_),
    .A(net796),
    .B(net1334));
 sg13g2_nand3_1 _11521_ (.B(_05379_),
    .C(_05501_),
    .A(_05190_),
    .Y(_05502_));
 sg13g2_and2_1 _11522_ (.A(net1752),
    .B(_05502_),
    .X(_00391_));
 sg13g2_a21oi_1 _11523_ (.A1(net721),
    .A2(net1331),
    .Y(_05503_),
    .B1(_05198_));
 sg13g2_a21oi_1 _11524_ (.A1(_05383_),
    .A2(_05503_),
    .Y(_00392_),
    .B1(net1737));
 sg13g2_nand2_1 _11525_ (.Y(_05504_),
    .A(net836),
    .B(net1332));
 sg13g2_nand3_1 _11526_ (.B(_05387_),
    .C(_05504_),
    .A(_05206_),
    .Y(_05505_));
 sg13g2_and2_1 _11527_ (.A(net1752),
    .B(_05505_),
    .X(_00393_));
 sg13g2_nand2_1 _11528_ (.Y(_05506_),
    .A(net826),
    .B(net1332));
 sg13g2_nand3_1 _11529_ (.B(_05391_),
    .C(_05506_),
    .A(_05213_),
    .Y(_05507_));
 sg13g2_and2_1 _11530_ (.A(net1752),
    .B(_05507_),
    .X(_00394_));
 sg13g2_nand2_1 _11531_ (.Y(_05508_),
    .A(net805),
    .B(net1330));
 sg13g2_nand3_1 _11532_ (.B(_05396_),
    .C(_05508_),
    .A(_05220_),
    .Y(_05509_));
 sg13g2_and2_1 _11533_ (.A(net1753),
    .B(_05509_),
    .X(_00395_));
 sg13g2_nand2_1 _11534_ (.Y(_05510_),
    .A(_05228_),
    .B(_05403_));
 sg13g2_a21oi_1 _11535_ (.A1(net554),
    .A2(net1330),
    .Y(_05511_),
    .B1(_05510_));
 sg13g2_nor2_1 _11536_ (.A(net1734),
    .B(_05511_),
    .Y(_00396_));
 sg13g2_nand2_1 _11537_ (.Y(_05512_),
    .A(net814),
    .B(net1330));
 sg13g2_nand3_1 _11538_ (.B(_05409_),
    .C(_05512_),
    .A(_05238_),
    .Y(_05513_));
 sg13g2_and2_1 _11539_ (.A(net1751),
    .B(_05513_),
    .X(_00397_));
 sg13g2_a22oi_1 _11540_ (.Y(_05514_),
    .B1(net1328),
    .B2(_05412_),
    .A2(net1331),
    .A1(net746));
 sg13g2_a21oi_1 _11541_ (.A1(_05244_),
    .A2(_05514_),
    .Y(_00398_),
    .B1(net1735));
 sg13g2_nand2_1 _11542_ (.Y(_05515_),
    .A(_05260_),
    .B(_05422_));
 sg13g2_a21oi_1 _11543_ (.A1(net552),
    .A2(net1333),
    .Y(_05516_),
    .B1(_05515_));
 sg13g2_nor2_1 _11544_ (.A(net1738),
    .B(_05516_),
    .Y(_00399_));
 sg13g2_a21oi_1 _11545_ (.A1(net720),
    .A2(net1333),
    .Y(_05517_),
    .B1(_05428_));
 sg13g2_a21oi_1 _11546_ (.A1(_05269_),
    .A2(_05517_),
    .Y(_00400_),
    .B1(net1738));
 sg13g2_nand2_1 _11547_ (.Y(_05518_),
    .A(net827),
    .B(net1334));
 sg13g2_nand3_1 _11548_ (.B(_05435_),
    .C(_05518_),
    .A(_05277_),
    .Y(_05519_));
 sg13g2_and2_1 _11549_ (.A(net1757),
    .B(_05519_),
    .X(_00401_));
 sg13g2_a21oi_1 _11550_ (.A1(net747),
    .A2(net1336),
    .Y(_05520_),
    .B1(_05283_));
 sg13g2_a21oi_1 _11551_ (.A1(_05439_),
    .A2(_05520_),
    .Y(_00402_),
    .B1(net1739));
 sg13g2_a21oi_1 _11552_ (.A1(net712),
    .A2(net1336),
    .Y(_05521_),
    .B1(_05298_));
 sg13g2_a21oi_1 _11553_ (.A1(_05451_),
    .A2(_05521_),
    .Y(_00403_),
    .B1(net1739));
 sg13g2_nand2_1 _11554_ (.Y(_05522_),
    .A(_05310_),
    .B(_05455_));
 sg13g2_a21oi_1 _11555_ (.A1(net610),
    .A2(net1337),
    .Y(_05523_),
    .B1(_05522_));
 sg13g2_nor2_1 _11556_ (.A(net1740),
    .B(net611),
    .Y(_00404_));
 sg13g2_nand2_1 _11557_ (.Y(_05524_),
    .A(net788),
    .B(net1339));
 sg13g2_and2_1 _11558_ (.A(_05319_),
    .B(_05524_),
    .X(_05525_));
 sg13g2_a21oi_1 _11559_ (.A1(_05459_),
    .A2(_05525_),
    .Y(_00405_),
    .B1(net1740));
 sg13g2_o21ai_1 _11560_ (.B1(net1757),
    .Y(_05526_),
    .A1(net713),
    .A2(_05159_));
 sg13g2_a21oi_1 _11561_ (.A1(_05328_),
    .A2(_05464_),
    .Y(_00406_),
    .B1(_05526_));
 sg13g2_nand2_1 _11562_ (.Y(_05527_),
    .A(net819),
    .B(net1338));
 sg13g2_nand3_1 _11563_ (.B(_05472_),
    .C(_05527_),
    .A(_05339_),
    .Y(_05528_));
 sg13g2_and2_1 _11564_ (.A(net1759),
    .B(_05528_),
    .X(_00407_));
 sg13g2_a221oi_1 _11565_ (.B2(_05479_),
    .C1(net1740),
    .B1(_05348_),
    .A1(_05531_),
    .Y(_00408_),
    .A2(net1338));
 sg13g2_a21oi_1 _11566_ (.A1(net704),
    .A2(net1339),
    .Y(_05529_),
    .B1(_05485_));
 sg13g2_a21oi_1 _11567_ (.A1(_05356_),
    .A2(_05529_),
    .Y(_00409_),
    .B1(net1741));
 sg13g2_o21ai_1 _11568_ (.B1(net1759),
    .Y(_05530_),
    .A1(net651),
    .A2(_05159_));
 sg13g2_a21oi_1 _11569_ (.A1(_05361_),
    .A2(_05490_),
    .Y(_00410_),
    .B1(_05530_));
 sg13g2_dfrbpq_2 _11570_ (.RESET_B(net28),
    .D(_00030_),
    .Q(\cordic_inst.CASE_cordic_state_BITS_7_TO_3_0_262144_1_13107_ETC__q2[19] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_1 _11571_ (.RESET_B(net29),
    .D(_00022_),
    .Q(\cordic_inst.current_op[0] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 _11572_ (.RESET_B(net30),
    .D(_00023_),
    .Q(\cordic_inst.current_op[1] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 _11573_ (.RESET_B(net43),
    .D(_00024_),
    .Q(\cordic_inst.current_op[2] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 _11574_ (.RESET_B(net27),
    .D(_00025_),
    .Q(\cordic_inst.current_op[3] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 _11575_ (.RESET_B(net1788),
    .D(_00031_),
    .Q(\cordic_inst.MUX_cordic_state$write_1__VAL_1[64] ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_1 _11576_ (.RESET_B(net1761),
    .D(_00032_),
    .Q(\cordic_inst.MUX_cordic_state$write_1__VAL_1[65] ),
    .CLK(clknet_leaf_43_clk));
 sg13g2_dfrbpq_1 _11577_ (.RESET_B(net1788),
    .D(_00033_),
    .Q(\cordic_inst.MUX_cordic_state$write_1__VAL_1[66] ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_1 _11578_ (.RESET_B(net1755),
    .D(_00034_),
    .Q(\cordic_inst.MUX_cordic_state$write_1__VAL_1[67] ),
    .CLK(clknet_leaf_57_clk));
 sg13g2_dfrbpq_1 _11579_ (.RESET_B(net1762),
    .D(_00035_),
    .Q(\cordic_inst.MUX_cordic_state$write_1__VAL_1[68] ),
    .CLK(clknet_leaf_44_clk));
 sg13g2_dfrbpq_1 _11580_ (.RESET_B(net1761),
    .D(_00036_),
    .Q(\cordic_inst.MUX_cordic_state$write_1__VAL_1[69] ),
    .CLK(clknet_leaf_56_clk));
 sg13g2_dfrbpq_2 _11581_ (.RESET_B(net1788),
    .D(_00037_),
    .Q(\cordic_inst.MUX_cordic_state$write_1__VAL_1[70] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_2 _11582_ (.RESET_B(net1762),
    .D(_00038_),
    .Q(\cordic_inst.MUX_cordic_state$write_1__VAL_1[71] ),
    .CLK(clknet_leaf_44_clk));
 sg13g2_dfrbpq_1 _11583_ (.RESET_B(net1780),
    .D(_00039_),
    .Q(\cordic_inst.MUX_cordic_state$write_1__VAL_1[72] ),
    .CLK(clknet_leaf_40_clk));
 sg13g2_dfrbpq_1 _11584_ (.RESET_B(net1762),
    .D(_00040_),
    .Q(\cordic_inst.MUX_cordic_state$write_1__VAL_1[73] ),
    .CLK(clknet_leaf_43_clk));
 sg13g2_dfrbpq_1 _11585_ (.RESET_B(net1781),
    .D(_00041_),
    .Q(\cordic_inst.MUX_cordic_state$write_1__VAL_1[74] ),
    .CLK(clknet_leaf_40_clk));
 sg13g2_dfrbpq_2 _11586_ (.RESET_B(net1762),
    .D(_00042_),
    .Q(\cordic_inst.MUX_cordic_state$write_1__VAL_1[75] ),
    .CLK(clknet_leaf_43_clk));
 sg13g2_dfrbpq_2 _11587_ (.RESET_B(net1783),
    .D(_00043_),
    .Q(\cordic_inst.MUX_cordic_state$write_1__VAL_1[76] ),
    .CLK(clknet_leaf_39_clk));
 sg13g2_dfrbpq_1 _11588_ (.RESET_B(net1762),
    .D(_00044_),
    .Q(\cordic_inst.MUX_cordic_state$write_1__VAL_1[77] ),
    .CLK(clknet_leaf_46_clk));
 sg13g2_dfrbpq_1 _11589_ (.RESET_B(net1783),
    .D(_00045_),
    .Q(\cordic_inst.MUX_cordic_state$write_1__VAL_1[78] ),
    .CLK(clknet_leaf_39_clk));
 sg13g2_dfrbpq_2 _11590_ (.RESET_B(net1762),
    .D(_00046_),
    .Q(\cordic_inst.MUX_cordic_state$write_1__VAL_1[79] ),
    .CLK(clknet_leaf_46_clk));
 sg13g2_dfrbpq_1 _11591_ (.RESET_B(net1790),
    .D(_00047_),
    .Q(\cordic_inst.MUX_cordic_state$write_1__VAL_1[32] ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_2 _11592_ (.RESET_B(net1792),
    .D(_00048_),
    .Q(\cordic_inst.MUX_cordic_state$write_1__VAL_1[33] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_1 _11593_ (.RESET_B(net1781),
    .D(_00049_),
    .Q(\cordic_inst.MUX_cordic_state$write_1__VAL_1[34] ),
    .CLK(clknet_leaf_38_clk));
 sg13g2_dfrbpq_2 _11594_ (.RESET_B(net1792),
    .D(_00050_),
    .Q(\cordic_inst.MUX_cordic_state$write_1__VAL_1[35] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_1 _11595_ (.RESET_B(net1783),
    .D(_00051_),
    .Q(\cordic_inst.MUX_cordic_state$write_1__VAL_1[36] ),
    .CLK(clknet_leaf_38_clk));
 sg13g2_dfrbpq_1 _11596_ (.RESET_B(net1792),
    .D(_00052_),
    .Q(\cordic_inst.MUX_cordic_state$write_1__VAL_1[37] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_1 _11597_ (.RESET_B(net1787),
    .D(_00053_),
    .Q(\cordic_inst.MUX_cordic_state$write_1__VAL_1[38] ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_1 _11598_ (.RESET_B(net1783),
    .D(_00054_),
    .Q(\cordic_inst.MUX_cordic_state$write_1__VAL_1[39] ),
    .CLK(clknet_leaf_38_clk));
 sg13g2_dfrbpq_1 _11599_ (.RESET_B(net1790),
    .D(_00055_),
    .Q(\cordic_inst.MUX_cordic_state$write_1__VAL_1[40] ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_1 _11600_ (.RESET_B(net1790),
    .D(_00056_),
    .Q(\cordic_inst.MUX_cordic_state$write_1__VAL_1[41] ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_1 _11601_ (.RESET_B(net1781),
    .D(_00057_),
    .Q(\cordic_inst.MUX_cordic_state$write_1__VAL_1[42] ),
    .CLK(clknet_leaf_37_clk));
 sg13g2_dfrbpq_1 _11602_ (.RESET_B(net1791),
    .D(_00058_),
    .Q(\cordic_inst.MUX_cordic_state$write_1__VAL_1[43] ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_1 _11603_ (.RESET_B(net1791),
    .D(_00059_),
    .Q(\cordic_inst.MUX_cordic_state$write_1__VAL_1[44] ),
    .CLK(clknet_leaf_37_clk));
 sg13g2_dfrbpq_1 _11604_ (.RESET_B(net1790),
    .D(_00060_),
    .Q(\cordic_inst.MUX_cordic_state$write_1__VAL_1[45] ),
    .CLK(clknet_leaf_37_clk));
 sg13g2_dfrbpq_1 _11605_ (.RESET_B(net1779),
    .D(_00061_),
    .Q(\cordic_inst.MUX_cordic_state$write_1__VAL_1[46] ),
    .CLK(clknet_leaf_40_clk));
 sg13g2_dfrbpq_1 _11606_ (.RESET_B(net1781),
    .D(_00062_),
    .Q(\cordic_inst.MUX_cordic_state$write_1__VAL_1[47] ),
    .CLK(clknet_leaf_37_clk));
 sg13g2_dfrbpq_1 _11607_ (.RESET_B(net1773),
    .D(net351),
    .Q(\result_reg[24] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_1 _11608_ (.RESET_B(net1791),
    .D(net341),
    .Q(\result_reg[25] ),
    .CLK(clknet_leaf_36_clk));
 sg13g2_dfrbpq_1 _11609_ (.RESET_B(net1786),
    .D(net293),
    .Q(\result_reg[26] ),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_1 _11610_ (.RESET_B(net1773),
    .D(net301),
    .Q(\result_reg[27] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_1 _11611_ (.RESET_B(net1782),
    .D(net303),
    .Q(\result_reg[28] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_1 _11612_ (.RESET_B(net1773),
    .D(net283),
    .Q(\result_reg[29] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_1 _11613_ (.RESET_B(net1784),
    .D(net325),
    .Q(\result_reg[30] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_1 _11614_ (.RESET_B(net1778),
    .D(net411),
    .Q(\result_reg[31] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_2 _11615_ (.RESET_B(net1768),
    .D(net525),
    .Q(\result_reg[32] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_2 _11616_ (.RESET_B(net1767),
    .D(net479),
    .Q(\result_reg[33] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 _11617_ (.RESET_B(net1767),
    .D(net533),
    .Q(\result_reg[34] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 _11618_ (.RESET_B(net1767),
    .D(net403),
    .Q(\result_reg[35] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_2 _11619_ (.RESET_B(net1767),
    .D(net505),
    .Q(\result_reg[36] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_2 _11620_ (.RESET_B(net1767),
    .D(net432),
    .Q(\result_reg[37] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 _11621_ (.RESET_B(net1767),
    .D(net452),
    .Q(\result_reg[38] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 _11622_ (.RESET_B(net1772),
    .D(net390),
    .Q(\result_reg[39] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_1 _11623_ (.RESET_B(net1768),
    .D(net531),
    .Q(\result_reg[40] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 _11624_ (.RESET_B(net1784),
    .D(net317),
    .Q(\result_reg[41] ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_1 _11625_ (.RESET_B(net1772),
    .D(net321),
    .Q(\result_reg[42] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 _11626_ (.RESET_B(net1772),
    .D(net345),
    .Q(\result_reg[43] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 _11627_ (.RESET_B(net1782),
    .D(net382),
    .Q(\result_reg[44] ),
    .CLK(clknet_leaf_36_clk));
 sg13g2_dfrbpq_1 _11628_ (.RESET_B(net1782),
    .D(net481),
    .Q(\result_reg[45] ),
    .CLK(clknet_leaf_41_clk));
 sg13g2_dfrbpq_1 _11629_ (.RESET_B(net1778),
    .D(net333),
    .Q(\result_reg[46] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_1 _11630_ (.RESET_B(net1778),
    .D(net361),
    .Q(\result_reg[47] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_1 _11631_ (.RESET_B(net1786),
    .D(net419),
    .Q(\result_reg[48] ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_dfrbpq_1 _11632_ (.RESET_B(net1784),
    .D(net396),
    .Q(\result_reg[49] ),
    .CLK(clknet_leaf_31_clk));
 sg13g2_dfrbpq_1 _11633_ (.RESET_B(net1786),
    .D(net291),
    .Q(\result_reg[50] ),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_1 _11634_ (.RESET_B(net1786),
    .D(net467),
    .Q(\result_reg[51] ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_dfrbpq_1 _11635_ (.RESET_B(net1791),
    .D(_00091_),
    .Q(\result_reg[52] ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_1 _11636_ (.RESET_B(net1772),
    .D(net289),
    .Q(\result_reg[53] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_1 _11637_ (.RESET_B(net1772),
    .D(net331),
    .Q(\result_reg[54] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_1 _11638_ (.RESET_B(net1785),
    .D(net323),
    .Q(\result_reg[55] ),
    .CLK(clknet_leaf_31_clk));
 sg13g2_dfrbpq_1 _11639_ (.RESET_B(net1772),
    .D(_00095_),
    .Q(\result_reg[56] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 _11640_ (.RESET_B(net1785),
    .D(net384),
    .Q(\result_reg[57] ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_1 _11641_ (.RESET_B(net1786),
    .D(_00097_),
    .Q(\result_reg[58] ),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_1 _11642_ (.RESET_B(net1772),
    .D(net349),
    .Q(\result_reg[59] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 _11643_ (.RESET_B(net1773),
    .D(net309),
    .Q(\result_reg[60] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_1 _11644_ (.RESET_B(net1785),
    .D(net347),
    .Q(\result_reg[61] ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_1 _11645_ (.RESET_B(net1791),
    .D(_00101_),
    .Q(\result_reg[62] ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_1 _11646_ (.RESET_B(net1790),
    .D(net364),
    .Q(\result_reg[63] ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_1 _11647_ (.RESET_B(net1791),
    .D(net394),
    .Q(\result_reg[64] ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_1 _11648_ (.RESET_B(net1790),
    .D(net441),
    .Q(\result_reg[65] ),
    .CLK(clknet_leaf_36_clk));
 sg13g2_dfrbpq_1 _11649_ (.RESET_B(net1790),
    .D(_00105_),
    .Q(\result_reg[66] ),
    .CLK(clknet_leaf_36_clk));
 sg13g2_dfrbpq_1 _11650_ (.RESET_B(net1765),
    .D(net285),
    .Q(\result_reg[67] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_1 _11651_ (.RESET_B(net1778),
    .D(net327),
    .Q(\result_reg[68] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_2 _11652_ (.RESET_B(net1781),
    .D(net475),
    .Q(\result_reg[69] ),
    .CLK(clknet_leaf_36_clk));
 sg13g2_dfrbpq_2 _11653_ (.RESET_B(net1782),
    .D(_00109_),
    .Q(\result_reg[70] ),
    .CLK(clknet_leaf_37_clk));
 sg13g2_dfrbpq_2 _11654_ (.RESET_B(net1781),
    .D(net380),
    .Q(\result_reg[71] ),
    .CLK(clknet_leaf_37_clk));
 sg13g2_dfrbpq_2 _11655_ (.RESET_B(net92),
    .D(_00001_),
    .Q(\cordic_inst.CASE_cordic_state_BITS_7_TO_3_0_3217_1_1901_2__ETC__q3[1] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_1 _11656_ (.RESET_B(net93),
    .D(_00002_),
    .Q(\cordic_inst.CASE_cordic_state_BITS_7_TO_3_0_3217_1_1901_2__ETC__q3[3] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_1 _11657_ (.RESET_B(net94),
    .D(_00003_),
    .Q(\cordic_inst.CASE_cordic_state_BITS_7_TO_3_0_3217_1_1901_2__ETC__q3[5] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_1 _11658_ (.RESET_B(net95),
    .D(_00004_),
    .Q(\cordic_inst.CASE_cordic_state_BITS_7_TO_3_0_3217_1_1901_2__ETC__q3[7] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_1 _11659_ (.RESET_B(net164),
    .D(_00005_),
    .Q(\cordic_inst.CASE_cordic_state_BITS_7_TO_3_0_3217_1_1901_2__ETC__q3[9] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_1 _11660_ (.RESET_B(net273),
    .D(_00000_),
    .Q(\cordic_inst.CASE_cordic_state_BITS_7_TO_3_0_3217_1_1901_2__ETC__q3[11] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_1 _11661_ (.RESET_B(net272),
    .D(_00111_),
    .Q(\cordic_inst.CASE_cordic_state_BITS_7_TO_3_0_3217_1_1901_2__ETC__q3[6] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_1 _11662_ (.RESET_B(net271),
    .D(_00112_),
    .Q(\cordic_inst.CASE_cordic_state_BITS_7_TO_3_0_3217_1_1901_2__ETC__q3[8] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_2 _11663_ (.RESET_B(net270),
    .D(_00113_),
    .Q(\cordic_inst.CASE_cordic_state_BITS_7_TO_3_0_3217_1_1901_2__ETC__q3[0] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_1 _11664_ (.RESET_B(net269),
    .D(_00114_),
    .Q(\cordic_inst.CASE_cordic_state_BITS_7_TO_3_0_3217_1_1901_2__ETC__q3[2] ),
    .CLK(clknet_leaf_68_clk));
 sg13g2_dfrbpq_1 _11665_ (.RESET_B(net268),
    .D(_00115_),
    .Q(\cordic_inst.CASE_cordic_state_BITS_7_TO_3_0_3217_1_1901_2__ETC__q3[4] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_1 _11666_ (.RESET_B(net267),
    .D(_00116_),
    .Q(\cordic_inst.CASE_cordic_state_BITS_7_TO_3_0_3217_1_1901_2__ETC__q3[10] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_2 _11667_ (.RESET_B(net1774),
    .D(_00118_),
    .Q(uo_out[0]),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_2 _11668_ (.RESET_B(net1776),
    .D(_00119_),
    .Q(uo_out[1]),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_2 _11669_ (.RESET_B(net1774),
    .D(_00120_),
    .Q(uo_out[2]),
    .CLK(clknet_leaf_28_clk));
 sg13g2_dfrbpq_1 _11670_ (.RESET_B(net1776),
    .D(_00121_),
    .Q(uo_out[3]),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_2 _11671_ (.RESET_B(net1774),
    .D(_00122_),
    .Q(uo_out[4]),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_1 _11672_ (.RESET_B(net1776),
    .D(_00123_),
    .Q(uo_out[5]),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_2 _11673_ (.RESET_B(net1776),
    .D(_00124_),
    .Q(uo_out[6]),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_2 _11674_ (.RESET_B(net1774),
    .D(net756),
    .Q(uo_out[7]),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_2 _11675_ (.RESET_B(net1774),
    .D(net725),
    .Q(\state[0] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_2 _11676_ (.RESET_B(net1775),
    .D(_00127_),
    .Q(\state[1] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_1 _11677_ (.RESET_B(net1774),
    .D(_00128_),
    .Q(\state[2] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_2 _11678_ (.RESET_B(net1787),
    .D(_00129_),
    .Q(\cmd_reg[0] ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_dfrbpq_2 _11679_ (.RESET_B(net1787),
    .D(net694),
    .Q(\cmd_reg[1] ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_dfrbpq_2 _11680_ (.RESET_B(net1787),
    .D(net719),
    .Q(\cmd_reg[2] ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_2 _11681_ (.RESET_B(net1775),
    .D(net692),
    .Q(\cmd_reg[3] ),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_1 _11682_ (.RESET_B(net1787),
    .D(net626),
    .Q(\cmd_reg[4] ),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_1 _11683_ (.RESET_B(net1787),
    .D(net620),
    .Q(\cmd_reg[5] ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_dfrbpq_1 _11684_ (.RESET_B(net1787),
    .D(net583),
    .Q(\cmd_reg[6] ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_1 _11685_ (.RESET_B(net1787),
    .D(net569),
    .Q(\cmd_reg[7] ),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_1 _11686_ (.RESET_B(net1792),
    .D(_00137_),
    .Q(\cordic_inst.MUX_cordic_state$write_1__VAL_1[56] ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_2 _11687_ (.RESET_B(net1763),
    .D(_00138_),
    .Q(\cordic_inst.MUX_cordic_state$write_1__VAL_1[57] ),
    .CLK(clknet_leaf_40_clk));
 sg13g2_dfrbpq_2 _11688_ (.RESET_B(net1790),
    .D(_00139_),
    .Q(\cordic_inst.MUX_cordic_state$write_1__VAL_1[58] ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_1 _11689_ (.RESET_B(net1755),
    .D(_00140_),
    .Q(\cordic_inst.MUX_cordic_state$write_1__VAL_1[59] ),
    .CLK(clknet_leaf_57_clk));
 sg13g2_dfrbpq_1 _11690_ (.RESET_B(net1788),
    .D(_00141_),
    .Q(\cordic_inst.MUX_cordic_state$write_1__VAL_1[60] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_2 _11691_ (.RESET_B(net1763),
    .D(_00142_),
    .Q(\cordic_inst.MUX_cordic_state$write_1__VAL_1[61] ),
    .CLK(clknet_leaf_40_clk));
 sg13g2_dfrbpq_1 _11692_ (.RESET_B(net1792),
    .D(_00143_),
    .Q(\cordic_inst.MUX_cordic_state$write_1__VAL_1[62] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_2 _11693_ (.RESET_B(net1761),
    .D(_00144_),
    .Q(\cordic_inst.MUX_cordic_state$write_1__VAL_1[63] ),
    .CLK(clknet_leaf_44_clk));
 sg13g2_dfrbpq_1 _11694_ (.RESET_B(net1779),
    .D(_00145_),
    .Q(\cordic_inst.MUX_cordic_state$write_1__VAL_1[48] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_2 _11695_ (.RESET_B(net1782),
    .D(_00146_),
    .Q(\cordic_inst.MUX_cordic_state$write_1__VAL_1[49] ),
    .CLK(clknet_leaf_37_clk));
 sg13g2_dfrbpq_1 _11696_ (.RESET_B(net1782),
    .D(_00147_),
    .Q(\cordic_inst.MUX_cordic_state$write_1__VAL_1[50] ),
    .CLK(clknet_leaf_38_clk));
 sg13g2_dfrbpq_1 _11697_ (.RESET_B(net1781),
    .D(_00148_),
    .Q(\cordic_inst.MUX_cordic_state$write_1__VAL_1[51] ),
    .CLK(clknet_leaf_38_clk));
 sg13g2_dfrbpq_1 _11698_ (.RESET_B(net1781),
    .D(_00149_),
    .Q(\cordic_inst.MUX_cordic_state$write_1__VAL_1[52] ),
    .CLK(clknet_leaf_39_clk));
 sg13g2_dfrbpq_2 _11699_ (.RESET_B(net1783),
    .D(_00150_),
    .Q(\cordic_inst.MUX_cordic_state$write_1__VAL_1[53] ),
    .CLK(clknet_leaf_39_clk));
 sg13g2_dfrbpq_2 _11700_ (.RESET_B(net1783),
    .D(_00151_),
    .Q(\cordic_inst.MUX_cordic_state$write_1__VAL_1[54] ),
    .CLK(clknet_leaf_39_clk));
 sg13g2_dfrbpq_1 _11701_ (.RESET_B(net1783),
    .D(_00152_),
    .Q(\cordic_inst.MUX_cordic_state$write_1__VAL_1[55] ),
    .CLK(clknet_leaf_39_clk));
 sg13g2_dfrbpq_1 _11702_ (.RESET_B(net1785),
    .D(net329),
    .Q(\result_reg[0] ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_1 _11703_ (.RESET_B(net1784),
    .D(net335),
    .Q(\result_reg[1] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_1 _11704_ (.RESET_B(net1786),
    .D(net386),
    .Q(\result_reg[2] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_1 _11705_ (.RESET_B(net1766),
    .D(net313),
    .Q(\result_reg[3] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_1 _11706_ (.RESET_B(net1779),
    .D(net305),
    .Q(\result_reg[4] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_1 _11707_ (.RESET_B(net1779),
    .D(net319),
    .Q(\result_reg[5] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_1 _11708_ (.RESET_B(net1766),
    .D(net281),
    .Q(\result_reg[6] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_1 _11709_ (.RESET_B(net1778),
    .D(net307),
    .Q(\result_reg[7] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_1 _11710_ (.RESET_B(net1766),
    .D(net343),
    .Q(\result_reg[8] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_1 _11711_ (.RESET_B(net1772),
    .D(net357),
    .Q(\result_reg[9] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_1 _11712_ (.RESET_B(net1779),
    .D(net295),
    .Q(\result_reg[10] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_1 _11713_ (.RESET_B(net1773),
    .D(net297),
    .Q(\result_reg[11] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_1 _11714_ (.RESET_B(net1773),
    .D(net577),
    .Q(\result_reg[12] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_1 _11715_ (.RESET_B(net1779),
    .D(net287),
    .Q(\result_reg[13] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_1 _11716_ (.RESET_B(net1777),
    .D(net567),
    .Q(\result_reg[14] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_1 _11717_ (.RESET_B(net1778),
    .D(net572),
    .Q(\result_reg[15] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_1 _11718_ (.RESET_B(net1786),
    .D(net606),
    .Q(\result_reg[16] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_1 _11719_ (.RESET_B(net1784),
    .D(net388),
    .Q(\result_reg[17] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_1 _11720_ (.RESET_B(net1779),
    .D(net299),
    .Q(\result_reg[18] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_1 _11721_ (.RESET_B(net1766),
    .D(net339),
    .Q(\result_reg[19] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_1 _11722_ (.RESET_B(net1778),
    .D(net315),
    .Q(\result_reg[20] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_1 _11723_ (.RESET_B(net1784),
    .D(net311),
    .Q(\result_reg[21] ),
    .CLK(clknet_leaf_31_clk));
 sg13g2_dfrbpq_1 _11724_ (.RESET_B(net1784),
    .D(net337),
    .Q(\result_reg[22] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_1 _11725_ (.RESET_B(net1784),
    .D(net353),
    .Q(\result_reg[23] ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_1 _11726_ (.RESET_B(net1774),
    .D(net9),
    .Q(wr_prev),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_1 _11727_ (.RESET_B(net1774),
    .D(net10),
    .Q(rd_prev),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_2 _11728_ (.RESET_B(net1768),
    .D(_00013_),
    .Q(cordic_en_sin_cos),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 _11729_ (.RESET_B(net1773),
    .D(_00007_),
    .Q(cordic_en_atan2),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_2 _11730_ (.RESET_B(net1770),
    .D(_00014_),
    .Q(cordic_en_sqrt),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_2 _11731_ (.RESET_B(net1767),
    .D(_00012_),
    .Q(cordic_en_normalize),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 _11732_ (.RESET_B(net1770),
    .D(_00010_),
    .Q(cordic_en_get_sin_cos),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 _11733_ (.RESET_B(net1770),
    .D(_00008_),
    .Q(cordic_en_get_atan2),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 _11734_ (.RESET_B(net1770),
    .D(_00011_),
    .Q(cordic_en_get_sqrt),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 _11735_ (.RESET_B(net1770),
    .D(_00009_),
    .Q(cordic_en_get_normalize),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 _11736_ (.RESET_B(net1769),
    .D(_00021_),
    .Q(mac_en_multiply),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 _11737_ (.RESET_B(net1770),
    .D(_00018_),
    .Q(mac_en_get_multiply),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_2 _11738_ (.RESET_B(net1771),
    .D(_00019_),
    .Q(mac_en_mac),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 _11739_ (.RESET_B(net1769),
    .D(_00016_),
    .Q(mac_en_get_mac),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_2 _11740_ (.RESET_B(net1776),
    .D(_00020_),
    .Q(mac_en_msu),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_1 _11741_ (.RESET_B(net1769),
    .D(_00017_),
    .Q(mac_en_get_msu),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_2 _11742_ (.RESET_B(net1751),
    .D(_00015_),
    .Q(mac_en_clear),
    .CLK(clknet_leaf_64_clk));
 sg13g2_dfrbpq_1 _11743_ (.RESET_B(net1775),
    .D(_00177_),
    .Q(\byte_counter[0] ),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_2 _11744_ (.RESET_B(net1775),
    .D(net775),
    .Q(\byte_counter[1] ),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_2 _11745_ (.RESET_B(net1775),
    .D(net669),
    .Q(\byte_counter[2] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_2 _11746_ (.RESET_B(net1775),
    .D(net773),
    .Q(\byte_counter[3] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_1 _11747_ (.RESET_B(net266),
    .D(_00181_),
    .Q(\cordic_inst.IF_IF_cordic_state_BITS_2_TO_1_EQ_1_THEN_NOT_c_ETC___d36[1] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_2 _11748_ (.RESET_B(net264),
    .D(_00182_),
    .Q(cordic_busy),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_2 _11749_ (.RESET_B(net262),
    .D(net717),
    .Q(\cordic_inst.cordic_state[0] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 _11750_ (.RESET_B(net260),
    .D(_00184_),
    .Q(\cordic_inst.cordic_state[3] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_2 _11751_ (.RESET_B(net258),
    .D(_00185_),
    .Q(\cordic_inst.cordic_state[4] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _11752_ (.RESET_B(net256),
    .D(_00186_),
    .Q(\cordic_inst.cordic_state[5] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_2 _11753_ (.RESET_B(net254),
    .D(_00187_),
    .Q(\cordic_inst.cordic_state[6] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_1 _11754_ (.RESET_B(net252),
    .D(_00188_),
    .Q(\cordic_inst.cordic_state[7] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_2 _11755_ (.RESET_B(net250),
    .D(net673),
    .Q(\cordic_atan2_result[0] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_2 _11756_ (.RESET_B(net248),
    .D(_00190_),
    .Q(\cordic_atan2_result[1] ),
    .CLK(clknet_leaf_55_clk));
 sg13g2_dfrbpq_2 _11757_ (.RESET_B(net246),
    .D(_00191_),
    .Q(\cordic_atan2_result[2] ),
    .CLK(clknet_leaf_58_clk));
 sg13g2_dfrbpq_2 _11758_ (.RESET_B(net244),
    .D(_00192_),
    .Q(\cordic_atan2_result[3] ),
    .CLK(clknet_leaf_57_clk));
 sg13g2_dfrbpq_2 _11759_ (.RESET_B(net242),
    .D(_00193_),
    .Q(\cordic_atan2_result[4] ),
    .CLK(clknet_leaf_58_clk));
 sg13g2_dfrbpq_2 _11760_ (.RESET_B(net240),
    .D(_00194_),
    .Q(\cordic_atan2_result[5] ),
    .CLK(clknet_leaf_59_clk));
 sg13g2_dfrbpq_2 _11761_ (.RESET_B(net238),
    .D(_00195_),
    .Q(\cordic_atan2_result[6] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_2 _11762_ (.RESET_B(net236),
    .D(_00196_),
    .Q(\cordic_atan2_result[7] ),
    .CLK(clknet_leaf_60_clk));
 sg13g2_dfrbpq_2 _11763_ (.RESET_B(net234),
    .D(_00197_),
    .Q(\cordic_atan2_result[8] ),
    .CLK(clknet_leaf_68_clk));
 sg13g2_dfrbpq_2 _11764_ (.RESET_B(net232),
    .D(_00198_),
    .Q(\cordic_atan2_result[9] ),
    .CLK(clknet_leaf_68_clk));
 sg13g2_dfrbpq_1 _11765_ (.RESET_B(net230),
    .D(net585),
    .Q(\cordic_atan2_result[10] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_2 _11766_ (.RESET_B(net228),
    .D(_00200_),
    .Q(\cordic_atan2_result[11] ),
    .CLK(clknet_leaf_59_clk));
 sg13g2_dfrbpq_2 _11767_ (.RESET_B(net226),
    .D(_00201_),
    .Q(\cordic_atan2_result[12] ),
    .CLK(clknet_leaf_57_clk));
 sg13g2_dfrbpq_2 _11768_ (.RESET_B(net224),
    .D(_00202_),
    .Q(\cordic_atan2_result[13] ),
    .CLK(clknet_leaf_56_clk));
 sg13g2_dfrbpq_2 _11769_ (.RESET_B(net222),
    .D(_00203_),
    .Q(\cordic_atan2_result[14] ),
    .CLK(clknet_leaf_56_clk));
 sg13g2_dfrbpq_1 _11770_ (.RESET_B(net220),
    .D(_00204_),
    .Q(\cordic_atan2_result[15] ),
    .CLK(clknet_leaf_56_clk));
 sg13g2_dfrbpq_2 _11771_ (.RESET_B(net218),
    .D(_00205_),
    .Q(\cordic_atan2_result[16] ),
    .CLK(clknet_leaf_56_clk));
 sg13g2_dfrbpq_2 _11772_ (.RESET_B(net216),
    .D(_00206_),
    .Q(\cordic_atan2_result[17] ),
    .CLK(clknet_leaf_55_clk));
 sg13g2_dfrbpq_2 _11773_ (.RESET_B(net214),
    .D(_00207_),
    .Q(\cordic_atan2_result[18] ),
    .CLK(clknet_leaf_55_clk));
 sg13g2_dfrbpq_2 _11774_ (.RESET_B(net212),
    .D(_00208_),
    .Q(\cordic_atan2_result[19] ),
    .CLK(clknet_leaf_55_clk));
 sg13g2_dfrbpq_2 _11775_ (.RESET_B(net210),
    .D(_00209_),
    .Q(\cordic_atan2_result[20] ),
    .CLK(clknet_leaf_45_clk));
 sg13g2_dfrbpq_2 _11776_ (.RESET_B(net208),
    .D(_00210_),
    .Q(\cordic_atan2_result[21] ),
    .CLK(clknet_leaf_44_clk));
 sg13g2_dfrbpq_2 _11777_ (.RESET_B(net206),
    .D(_00211_),
    .Q(\cordic_atan2_result[22] ),
    .CLK(clknet_leaf_45_clk));
 sg13g2_dfrbpq_2 _11778_ (.RESET_B(net204),
    .D(_00212_),
    .Q(\cordic_atan2_result[23] ),
    .CLK(clknet_leaf_45_clk));
 sg13g2_dfrbpq_2 _11779_ (.RESET_B(net202),
    .D(net787),
    .Q(\cordic_inst.cordic_state[32] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_2 _11780_ (.RESET_B(net200),
    .D(_00214_),
    .Q(\cordic_inst.cordic_state[33] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_2 _11781_ (.RESET_B(net198),
    .D(net700),
    .Q(\cordic_inst.cordic_state[34] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_2 _11782_ (.RESET_B(net196),
    .D(_00216_),
    .Q(\cordic_inst.cordic_state[35] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_2 _11783_ (.RESET_B(net194),
    .D(_00217_),
    .Q(\cordic_inst.cordic_state[36] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_1 _11784_ (.RESET_B(net192),
    .D(_00218_),
    .Q(\cordic_inst.cordic_state[37] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_1 _11785_ (.RESET_B(net190),
    .D(net702),
    .Q(\cordic_inst.cordic_state[38] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_1 _11786_ (.RESET_B(net188),
    .D(_00220_),
    .Q(\cordic_inst.cordic_state[39] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_1 _11787_ (.RESET_B(net186),
    .D(net829),
    .Q(\cordic_inst.cordic_state[40] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_1 _11788_ (.RESET_B(net184),
    .D(_00222_),
    .Q(\cordic_inst.cordic_state[41] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_2 _11789_ (.RESET_B(net182),
    .D(_00223_),
    .Q(\cordic_inst.cordic_state[42] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_2 _11790_ (.RESET_B(net180),
    .D(_00224_),
    .Q(\cordic_inst.cordic_state[43] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 _11791_ (.RESET_B(net178),
    .D(_00225_),
    .Q(\cordic_inst.cordic_state[44] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_2 _11792_ (.RESET_B(net176),
    .D(_00226_),
    .Q(\cordic_inst.cordic_state[45] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_1 _11793_ (.RESET_B(net174),
    .D(_00227_),
    .Q(\cordic_inst.cordic_state[46] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 _11794_ (.RESET_B(net172),
    .D(_00228_),
    .Q(\cordic_inst.cordic_state[47] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 _11795_ (.RESET_B(net170),
    .D(_00229_),
    .Q(\cordic_inst.cordic_state[48] ),
    .CLK(clknet_4_8_0_clk));
 sg13g2_dfrbpq_2 _11796_ (.RESET_B(net168),
    .D(_00230_),
    .Q(\cordic_inst.cordic_state[49] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 _11797_ (.RESET_B(net166),
    .D(net706),
    .Q(\cordic_inst.cordic_state[50] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_2 _11798_ (.RESET_B(net163),
    .D(_00232_),
    .Q(\cordic_inst.cordic_state[51] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_1 _11799_ (.RESET_B(net161),
    .D(_00233_),
    .Q(\cordic_inst.cordic_state[52] ),
    .CLK(clknet_leaf_42_clk));
 sg13g2_dfrbpq_2 _11800_ (.RESET_B(net159),
    .D(_00234_),
    .Q(\cordic_inst.cordic_state[53] ),
    .CLK(clknet_leaf_41_clk));
 sg13g2_dfrbpq_1 _11801_ (.RESET_B(net157),
    .D(_00235_),
    .Q(\cordic_inst.cordic_state[54] ),
    .CLK(clknet_leaf_41_clk));
 sg13g2_dfrbpq_1 _11802_ (.RESET_B(net155),
    .D(_00236_),
    .Q(\cordic_inst.cordic_state[55] ),
    .CLK(clknet_leaf_42_clk));
 sg13g2_dfrbpq_2 _11803_ (.RESET_B(net153),
    .D(net765),
    .Q(\cordic_inst.cordic_state[56] ),
    .CLK(clknet_leaf_41_clk));
 sg13g2_dfrbpq_2 _11804_ (.RESET_B(net151),
    .D(net723),
    .Q(\cordic_inst.cordic_state[57] ),
    .CLK(clknet_leaf_41_clk));
 sg13g2_dfrbpq_2 _11805_ (.RESET_B(net149),
    .D(net780),
    .Q(\cordic_inst.cordic_state[58] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_2 _11806_ (.RESET_B(net147),
    .D(_00240_),
    .Q(\cordic_inst.cordic_state[59] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_2 _11807_ (.RESET_B(net145),
    .D(_00241_),
    .Q(\cordic_inst.cordic_state[60] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_2 _11808_ (.RESET_B(net143),
    .D(net750),
    .Q(\cordic_inst.cordic_state[61] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_2 _11809_ (.RESET_B(net141),
    .D(_00243_),
    .Q(\cordic_inst.cordic_state[62] ),
    .CLK(clknet_4_3_0_clk));
 sg13g2_dfrbpq_2 _11810_ (.RESET_B(net139),
    .D(net763),
    .Q(\cordic_inst.cordic_state[63] ),
    .CLK(clknet_leaf_42_clk));
 sg13g2_dfrbpq_2 _11811_ (.RESET_B(net137),
    .D(net770),
    .Q(\cordic_inst.cordic_state[64] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_2 _11812_ (.RESET_B(net135),
    .D(_00246_),
    .Q(\cordic_inst.cordic_state[65] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_2 _11813_ (.RESET_B(net133),
    .D(_00247_),
    .Q(\cordic_inst.cordic_state[66] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_2 _11814_ (.RESET_B(net131),
    .D(_00248_),
    .Q(\cordic_inst.cordic_state[67] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_2 _11815_ (.RESET_B(net129),
    .D(_00249_),
    .Q(\cordic_inst.cordic_state[68] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_2 _11816_ (.RESET_B(net127),
    .D(_00250_),
    .Q(\cordic_inst.cordic_state[69] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_2 _11817_ (.RESET_B(net125),
    .D(net753),
    .Q(\cordic_inst.cordic_state[70] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_2 _11818_ (.RESET_B(net123),
    .D(_00252_),
    .Q(\cordic_inst.cordic_state[71] ),
    .CLK(clknet_leaf_57_clk));
 sg13g2_dfrbpq_2 _11819_ (.RESET_B(net121),
    .D(_00253_),
    .Q(\cordic_inst.cordic_state[72] ),
    .CLK(clknet_leaf_43_clk));
 sg13g2_dfrbpq_2 _11820_ (.RESET_B(net119),
    .D(net778),
    .Q(\cordic_inst.cordic_state[73] ),
    .CLK(clknet_leaf_43_clk));
 sg13g2_dfrbpq_2 _11821_ (.RESET_B(net117),
    .D(_00255_),
    .Q(\cordic_inst.cordic_state[74] ),
    .CLK(clknet_leaf_57_clk));
 sg13g2_dfrbpq_2 _11822_ (.RESET_B(net115),
    .D(net785),
    .Q(\cordic_inst.cordic_state[75] ),
    .CLK(clknet_leaf_57_clk));
 sg13g2_dfrbpq_2 _11823_ (.RESET_B(net113),
    .D(net794),
    .Q(\cordic_inst.cordic_state[76] ),
    .CLK(clknet_leaf_43_clk));
 sg13g2_dfrbpq_2 _11824_ (.RESET_B(net111),
    .D(_00258_),
    .Q(\cordic_inst.cordic_state[77] ),
    .CLK(clknet_leaf_43_clk));
 sg13g2_dfrbpq_2 _11825_ (.RESET_B(net109),
    .D(net783),
    .Q(\cordic_inst.cordic_state[78] ),
    .CLK(clknet_leaf_43_clk));
 sg13g2_dfrbpq_1 _11826_ (.RESET_B(net107),
    .D(_00260_),
    .Q(\cordic_inst.cordic_state[79] ),
    .CLK(clknet_leaf_42_clk));
 sg13g2_dfrbpq_2 _11827_ (.RESET_B(net1769),
    .D(_00029_),
    .Q(_00028_),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 _11828_ (.RESET_B(net1769),
    .D(net665),
    .Q(\exec_phase[1] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_2 _11829_ (.RESET_B(net1769),
    .D(net575),
    .Q(\exec_phase[2] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 _11830_ (.RESET_B(net104),
    .D(_00261_),
    .Q(\cordic_inst.operation_pending ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 _11831_ (.RESET_B(net102),
    .D(net485),
    .Q(\cordic_inst.operation_started ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_2 _11832_ (.RESET_B(net100),
    .D(_00263_),
    .Q(\cordic_inst.result_ready ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 _11833_ (.RESET_B(net98),
    .D(_00264_),
    .Q(\cordic_inst.get_normalize[48] ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_dfrbpq_1 _11834_ (.RESET_B(net96),
    .D(_00265_),
    .Q(\cordic_inst.get_normalize[49] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_1 _11835_ (.RESET_B(net90),
    .D(_00266_),
    .Q(\cordic_inst.get_normalize[50] ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_1 _11836_ (.RESET_B(net88),
    .D(_00267_),
    .Q(\cordic_inst.get_normalize[51] ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_dfrbpq_1 _11837_ (.RESET_B(net86),
    .D(_00268_),
    .Q(\cordic_inst.get_normalize[52] ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_1 _11838_ (.RESET_B(net84),
    .D(_00269_),
    .Q(\cordic_inst.get_normalize[53] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_1 _11839_ (.RESET_B(net82),
    .D(_00270_),
    .Q(\cordic_inst.get_normalize[54] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_1 _11840_ (.RESET_B(net80),
    .D(_00271_),
    .Q(\cordic_inst.get_normalize[55] ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_1 _11841_ (.RESET_B(net78),
    .D(_00272_),
    .Q(\cordic_inst.get_normalize[56] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 _11842_ (.RESET_B(net76),
    .D(_00273_),
    .Q(\cordic_inst.get_normalize[57] ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_1 _11843_ (.RESET_B(net74),
    .D(_00274_),
    .Q(\cordic_inst.get_normalize[58] ),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_1 _11844_ (.RESET_B(net72),
    .D(_00275_),
    .Q(\cordic_inst.get_normalize[59] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 _11845_ (.RESET_B(net70),
    .D(_00276_),
    .Q(\cordic_inst.get_normalize[60] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_1 _11846_ (.RESET_B(net68),
    .D(_00277_),
    .Q(\cordic_inst.get_normalize[61] ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_1 _11847_ (.RESET_B(net66),
    .D(_00278_),
    .Q(\cordic_inst.get_normalize[62] ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_1 _11848_ (.RESET_B(net64),
    .D(_00279_),
    .Q(\cordic_inst.get_normalize[63] ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_1 _11849_ (.RESET_B(net62),
    .D(_00280_),
    .Q(\cordic_inst.get_normalize[64] ),
    .CLK(clknet_leaf_31_clk));
 sg13g2_dfrbpq_1 _11850_ (.RESET_B(net60),
    .D(_00281_),
    .Q(\cordic_inst.get_normalize[65] ),
    .CLK(clknet_leaf_36_clk));
 sg13g2_dfrbpq_1 _11851_ (.RESET_B(net58),
    .D(_00282_),
    .Q(\cordic_inst.get_normalize[66] ),
    .CLK(clknet_leaf_40_clk));
 sg13g2_dfrbpq_1 _11852_ (.RESET_B(net56),
    .D(_00283_),
    .Q(\cordic_inst.get_normalize[67] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_1 _11853_ (.RESET_B(net55),
    .D(_00284_),
    .Q(\cordic_inst.get_normalize[68] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_1 _11854_ (.RESET_B(net53),
    .D(_00285_),
    .Q(\cordic_inst.get_normalize[69] ),
    .CLK(clknet_leaf_37_clk));
 sg13g2_dfrbpq_1 _11855_ (.RESET_B(net51),
    .D(_00286_),
    .Q(\cordic_inst.get_normalize[70] ),
    .CLK(clknet_leaf_40_clk));
 sg13g2_dfrbpq_1 _11856_ (.RESET_B(net49),
    .D(_00287_),
    .Q(\cordic_inst.get_normalize[71] ),
    .CLK(clknet_leaf_38_clk));
 sg13g2_dfrbpq_1 _11857_ (.RESET_B(net47),
    .D(_00288_),
    .Q(\cordic_inst.get_normalize[24] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_1 _11858_ (.RESET_B(net45),
    .D(_00289_),
    .Q(\cordic_inst.get_normalize[25] ),
    .CLK(clknet_leaf_41_clk));
 sg13g2_dfrbpq_1 _11859_ (.RESET_B(net42),
    .D(_00290_),
    .Q(\cordic_inst.get_normalize[26] ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_1 _11860_ (.RESET_B(net40),
    .D(_00291_),
    .Q(\cordic_inst.get_normalize[27] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_1 _11861_ (.RESET_B(net38),
    .D(_00292_),
    .Q(\cordic_inst.get_normalize[28] ),
    .CLK(clknet_leaf_38_clk));
 sg13g2_dfrbpq_1 _11862_ (.RESET_B(net36),
    .D(_00293_),
    .Q(\cordic_inst.get_normalize[29] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 _11863_ (.RESET_B(net34),
    .D(_00294_),
    .Q(\cordic_inst.get_normalize[30] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_1 _11864_ (.RESET_B(net32),
    .D(_00295_),
    .Q(\cordic_inst.get_normalize[31] ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_1 _11865_ (.RESET_B(net265),
    .D(_00296_),
    .Q(\cordic_inst.get_normalize[32] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 _11866_ (.RESET_B(net261),
    .D(_00297_),
    .Q(\cordic_inst.get_normalize[33] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 _11867_ (.RESET_B(net257),
    .D(_00298_),
    .Q(\cordic_inst.get_normalize[34] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 _11868_ (.RESET_B(net253),
    .D(_00299_),
    .Q(\cordic_inst.get_normalize[35] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 _11869_ (.RESET_B(net249),
    .D(_00300_),
    .Q(\cordic_inst.get_normalize[36] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 _11870_ (.RESET_B(net245),
    .D(_00301_),
    .Q(\cordic_inst.get_normalize[37] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 _11871_ (.RESET_B(net241),
    .D(_00302_),
    .Q(\cordic_inst.get_normalize[38] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 _11872_ (.RESET_B(net237),
    .D(_00303_),
    .Q(\cordic_inst.get_normalize[39] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_1 _11873_ (.RESET_B(net233),
    .D(_00304_),
    .Q(\cordic_inst.get_normalize[40] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 _11874_ (.RESET_B(net229),
    .D(_00305_),
    .Q(\cordic_inst.get_normalize[41] ),
    .CLK(clknet_leaf_31_clk));
 sg13g2_dfrbpq_1 _11875_ (.RESET_B(net225),
    .D(_00306_),
    .Q(\cordic_inst.get_normalize[42] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 _11876_ (.RESET_B(net221),
    .D(_00307_),
    .Q(\cordic_inst.get_normalize[43] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_1 _11877_ (.RESET_B(net217),
    .D(_00308_),
    .Q(\cordic_inst.get_normalize[44] ),
    .CLK(clknet_leaf_38_clk));
 sg13g2_dfrbpq_1 _11878_ (.RESET_B(net213),
    .D(_00309_),
    .Q(\cordic_inst.get_normalize[45] ),
    .CLK(clknet_leaf_40_clk));
 sg13g2_dfrbpq_1 _11879_ (.RESET_B(net209),
    .D(_00310_),
    .Q(\cordic_inst.get_normalize[46] ),
    .CLK(clknet_leaf_41_clk));
 sg13g2_dfrbpq_1 _11880_ (.RESET_B(net205),
    .D(_00311_),
    .Q(\cordic_inst.get_normalize[47] ),
    .CLK(clknet_leaf_41_clk));
 sg13g2_dfrbpq_1 _11881_ (.RESET_B(net201),
    .D(_00312_),
    .Q(\mac_inst.get_multiply[0] ),
    .CLK(clknet_leaf_47_clk));
 sg13g2_dfrbpq_1 _11882_ (.RESET_B(net197),
    .D(net617),
    .Q(\mac_inst.get_multiply[1] ),
    .CLK(clknet_leaf_47_clk));
 sg13g2_dfrbpq_1 _11883_ (.RESET_B(net193),
    .D(_00314_),
    .Q(\mac_inst.get_multiply[2] ),
    .CLK(clknet_leaf_54_clk));
 sg13g2_dfrbpq_1 _11884_ (.RESET_B(net189),
    .D(_00315_),
    .Q(\mac_inst.get_multiply[3] ),
    .CLK(clknet_leaf_56_clk));
 sg13g2_dfrbpq_1 _11885_ (.RESET_B(net185),
    .D(net604),
    .Q(\mac_inst.get_multiply[4] ),
    .CLK(clknet_leaf_61_clk));
 sg13g2_dfrbpq_1 _11886_ (.RESET_B(net181),
    .D(_00317_),
    .Q(\mac_inst.get_multiply[5] ),
    .CLK(clknet_leaf_58_clk));
 sg13g2_dfrbpq_1 _11887_ (.RESET_B(net177),
    .D(_00318_),
    .Q(\mac_inst.get_multiply[6] ),
    .CLK(clknet_leaf_61_clk));
 sg13g2_dfrbpq_1 _11888_ (.RESET_B(net173),
    .D(_00319_),
    .Q(\mac_inst.get_multiply[7] ),
    .CLK(clknet_leaf_61_clk));
 sg13g2_dfrbpq_1 _11889_ (.RESET_B(net169),
    .D(_00320_),
    .Q(\mac_inst.get_multiply[8] ),
    .CLK(clknet_leaf_68_clk));
 sg13g2_dfrbpq_1 _11890_ (.RESET_B(net165),
    .D(_00321_),
    .Q(\mac_inst.get_multiply[9] ),
    .CLK(clknet_leaf_68_clk));
 sg13g2_dfrbpq_1 _11891_ (.RESET_B(net160),
    .D(_00322_),
    .Q(\mac_inst.get_multiply[10] ),
    .CLK(clknet_leaf_65_clk));
 sg13g2_dfrbpq_1 _11892_ (.RESET_B(net156),
    .D(_00323_),
    .Q(\mac_inst.get_multiply[11] ),
    .CLK(clknet_leaf_61_clk));
 sg13g2_dfrbpq_1 _11893_ (.RESET_B(net152),
    .D(_00324_),
    .Q(\mac_inst.get_multiply[12] ),
    .CLK(clknet_leaf_61_clk));
 sg13g2_dfrbpq_1 _11894_ (.RESET_B(net148),
    .D(_00325_),
    .Q(\mac_inst.get_multiply[13] ),
    .CLK(clknet_leaf_54_clk));
 sg13g2_dfrbpq_1 _11895_ (.RESET_B(net144),
    .D(_00326_),
    .Q(\mac_inst.get_multiply[14] ),
    .CLK(clknet_leaf_54_clk));
 sg13g2_dfrbpq_1 _11896_ (.RESET_B(net140),
    .D(_00327_),
    .Q(\mac_inst.get_multiply[15] ),
    .CLK(clknet_leaf_54_clk));
 sg13g2_dfrbpq_1 _11897_ (.RESET_B(net136),
    .D(net623),
    .Q(\mac_inst.get_multiply[16] ),
    .CLK(clknet_leaf_52_clk));
 sg13g2_dfrbpq_1 _11898_ (.RESET_B(net132),
    .D(_00329_),
    .Q(\mac_inst.get_multiply[17] ),
    .CLK(clknet_leaf_50_clk));
 sg13g2_dfrbpq_1 _11899_ (.RESET_B(net128),
    .D(net630),
    .Q(\mac_inst.get_multiply[18] ),
    .CLK(clknet_leaf_50_clk));
 sg13g2_dfrbpq_1 _11900_ (.RESET_B(net124),
    .D(_00331_),
    .Q(\mac_inst.get_multiply[19] ),
    .CLK(clknet_leaf_51_clk));
 sg13g2_dfrbpq_1 _11901_ (.RESET_B(net120),
    .D(_00332_),
    .Q(\mac_inst.get_multiply[20] ),
    .CLK(clknet_leaf_48_clk));
 sg13g2_dfrbpq_1 _11902_ (.RESET_B(net116),
    .D(_00333_),
    .Q(\mac_inst.get_multiply[21] ),
    .CLK(clknet_leaf_48_clk));
 sg13g2_dfrbpq_1 _11903_ (.RESET_B(net112),
    .D(_00334_),
    .Q(\mac_inst.get_multiply[22] ),
    .CLK(clknet_leaf_48_clk));
 sg13g2_dfrbpq_1 _11904_ (.RESET_B(net108),
    .D(net660),
    .Q(\mac_inst.get_multiply[23] ),
    .CLK(clknet_leaf_48_clk));
 sg13g2_dfrbpq_1 _11905_ (.RESET_B(net105),
    .D(_00336_),
    .Q(\mac_inst.get_msu[0] ),
    .CLK(clknet_leaf_50_clk));
 sg13g2_dfrbpq_1 _11906_ (.RESET_B(net101),
    .D(net367),
    .Q(\mac_inst.get_msu[1] ),
    .CLK(clknet_leaf_51_clk));
 sg13g2_dfrbpq_1 _11907_ (.RESET_B(net97),
    .D(_00338_),
    .Q(\mac_inst.get_msu[2] ),
    .CLK(clknet_leaf_54_clk));
 sg13g2_dfrbpq_1 _11908_ (.RESET_B(net89),
    .D(_00339_),
    .Q(\mac_inst.get_msu[3] ),
    .CLK(clknet_leaf_56_clk));
 sg13g2_dfrbpq_1 _11909_ (.RESET_B(net85),
    .D(_00340_),
    .Q(\mac_inst.get_msu[4] ),
    .CLK(clknet_leaf_61_clk));
 sg13g2_dfrbpq_1 _11910_ (.RESET_B(net81),
    .D(_00341_),
    .Q(\mac_inst.get_msu[5] ),
    .CLK(clknet_leaf_58_clk));
 sg13g2_dfrbpq_1 _11911_ (.RESET_B(net77),
    .D(net373),
    .Q(\mac_inst.get_msu[6] ),
    .CLK(clknet_leaf_61_clk));
 sg13g2_dfrbpq_1 _11912_ (.RESET_B(net73),
    .D(_00343_),
    .Q(\mac_inst.get_msu[7] ),
    .CLK(clknet_leaf_61_clk));
 sg13g2_dfrbpq_1 _11913_ (.RESET_B(net69),
    .D(net596),
    .Q(\mac_inst.get_msu[8] ),
    .CLK(clknet_leaf_67_clk));
 sg13g2_dfrbpq_1 _11914_ (.RESET_B(net65),
    .D(net587),
    .Q(\mac_inst.get_msu[9] ),
    .CLK(clknet_leaf_67_clk));
 sg13g2_dfrbpq_1 _11915_ (.RESET_B(net61),
    .D(_00346_),
    .Q(\mac_inst.get_msu[10] ),
    .CLK(clknet_leaf_63_clk));
 sg13g2_dfrbpq_1 _11916_ (.RESET_B(net57),
    .D(_00347_),
    .Q(\mac_inst.get_msu[11] ),
    .CLK(clknet_leaf_63_clk));
 sg13g2_dfrbpq_1 _11917_ (.RESET_B(net54),
    .D(_00348_),
    .Q(\mac_inst.get_msu[12] ),
    .CLK(clknet_leaf_62_clk));
 sg13g2_dfrbpq_1 _11918_ (.RESET_B(net50),
    .D(net462),
    .Q(\mac_inst.get_msu[13] ),
    .CLK(clknet_leaf_62_clk));
 sg13g2_dfrbpq_1 _11919_ (.RESET_B(net46),
    .D(net535),
    .Q(\mac_inst.get_msu[14] ),
    .CLK(clknet_leaf_53_clk));
 sg13g2_dfrbpq_1 _11920_ (.RESET_B(net41),
    .D(_00351_),
    .Q(\mac_inst.get_msu[15] ),
    .CLK(clknet_leaf_52_clk));
 sg13g2_dfrbpq_1 _11921_ (.RESET_B(net37),
    .D(_00352_),
    .Q(\mac_inst.get_msu[16] ),
    .CLK(clknet_leaf_53_clk));
 sg13g2_dfrbpq_1 _11922_ (.RESET_B(net33),
    .D(net497),
    .Q(\mac_inst.get_msu[17] ),
    .CLK(clknet_leaf_52_clk));
 sg13g2_dfrbpq_1 _11923_ (.RESET_B(net263),
    .D(_00354_),
    .Q(\mac_inst.get_msu[18] ),
    .CLK(clknet_leaf_49_clk));
 sg13g2_dfrbpq_1 _11924_ (.RESET_B(net255),
    .D(net549),
    .Q(\mac_inst.get_msu[19] ),
    .CLK(clknet_leaf_52_clk));
 sg13g2_dfrbpq_1 _11925_ (.RESET_B(net247),
    .D(_00356_),
    .Q(\mac_inst.get_msu[20] ),
    .CLK(clknet_leaf_48_clk));
 sg13g2_dfrbpq_1 _11926_ (.RESET_B(net239),
    .D(_00357_),
    .Q(\mac_inst.get_msu[21] ),
    .CLK(clknet_leaf_48_clk));
 sg13g2_dfrbpq_1 _11927_ (.RESET_B(net231),
    .D(_00358_),
    .Q(\mac_inst.get_msu[22] ),
    .CLK(clknet_leaf_49_clk));
 sg13g2_dfrbpq_1 _11928_ (.RESET_B(net223),
    .D(_00359_),
    .Q(\mac_inst.get_msu[23] ),
    .CLK(clknet_leaf_50_clk));
 sg13g2_dfrbpq_1 _11929_ (.RESET_B(net215),
    .D(_00360_),
    .Q(\mac_inst.get_mac[0] ),
    .CLK(clknet_leaf_50_clk));
 sg13g2_dfrbpq_1 _11930_ (.RESET_B(net207),
    .D(_00361_),
    .Q(\mac_inst.get_mac[1] ),
    .CLK(clknet_leaf_55_clk));
 sg13g2_dfrbpq_1 _11931_ (.RESET_B(net199),
    .D(_00362_),
    .Q(\mac_inst.get_mac[2] ),
    .CLK(clknet_leaf_55_clk));
 sg13g2_dfrbpq_1 _11932_ (.RESET_B(net191),
    .D(_00363_),
    .Q(\mac_inst.get_mac[3] ),
    .CLK(clknet_leaf_56_clk));
 sg13g2_dfrbpq_1 _11933_ (.RESET_B(net183),
    .D(_00364_),
    .Q(\mac_inst.get_mac[4] ),
    .CLK(clknet_leaf_58_clk));
 sg13g2_dfrbpq_1 _11934_ (.RESET_B(net175),
    .D(_00365_),
    .Q(\mac_inst.get_mac[5] ),
    .CLK(clknet_leaf_59_clk));
 sg13g2_dfrbpq_1 _11935_ (.RESET_B(net167),
    .D(_00366_),
    .Q(\mac_inst.get_mac[6] ),
    .CLK(clknet_leaf_60_clk));
 sg13g2_dfrbpq_1 _11936_ (.RESET_B(net158),
    .D(_00367_),
    .Q(\mac_inst.get_mac[7] ),
    .CLK(clknet_4_0_0_clk));
 sg13g2_dfrbpq_1 _11937_ (.RESET_B(net150),
    .D(_00368_),
    .Q(\mac_inst.get_mac[8] ),
    .CLK(clknet_leaf_67_clk));
 sg13g2_dfrbpq_1 _11938_ (.RESET_B(net142),
    .D(net562),
    .Q(\mac_inst.get_mac[9] ),
    .CLK(clknet_leaf_67_clk));
 sg13g2_dfrbpq_1 _11939_ (.RESET_B(net134),
    .D(_00370_),
    .Q(\mac_inst.get_mac[10] ),
    .CLK(clknet_leaf_64_clk));
 sg13g2_dfrbpq_1 _11940_ (.RESET_B(net126),
    .D(net608),
    .Q(\mac_inst.get_mac[11] ),
    .CLK(clknet_leaf_63_clk));
 sg13g2_dfrbpq_2 _11941_ (.RESET_B(net118),
    .D(_00372_),
    .Q(\mac_inst.get_mac[12] ),
    .CLK(clknet_leaf_62_clk));
 sg13g2_dfrbpq_1 _11942_ (.RESET_B(net110),
    .D(_00373_),
    .Q(\mac_inst.get_mac[13] ),
    .CLK(clknet_leaf_53_clk));
 sg13g2_dfrbpq_1 _11943_ (.RESET_B(net103),
    .D(_00374_),
    .Q(\mac_inst.get_mac[14] ),
    .CLK(clknet_leaf_54_clk));
 sg13g2_dfrbpq_2 _11944_ (.RESET_B(net91),
    .D(net591),
    .Q(\mac_inst.get_mac[15] ),
    .CLK(clknet_leaf_53_clk));
 sg13g2_dfrbpq_2 _11945_ (.RESET_B(net83),
    .D(_00376_),
    .Q(\mac_inst.get_mac[16] ),
    .CLK(clknet_leaf_53_clk));
 sg13g2_dfrbpq_1 _11946_ (.RESET_B(net75),
    .D(net601),
    .Q(\mac_inst.get_mac[17] ),
    .CLK(clknet_leaf_52_clk));
 sg13g2_dfrbpq_1 _11947_ (.RESET_B(net67),
    .D(_00378_),
    .Q(\mac_inst.get_mac[18] ),
    .CLK(clknet_leaf_52_clk));
 sg13g2_dfrbpq_1 _11948_ (.RESET_B(net59),
    .D(_00379_),
    .Q(\mac_inst.get_mac[19] ),
    .CLK(clknet_leaf_52_clk));
 sg13g2_dfrbpq_2 _11949_ (.RESET_B(net52),
    .D(_00380_),
    .Q(\mac_inst.get_mac[20] ),
    .CLK(clknet_leaf_49_clk));
 sg13g2_dfrbpq_1 _11950_ (.RESET_B(net44),
    .D(net640),
    .Q(\mac_inst.get_mac[21] ),
    .CLK(clknet_leaf_47_clk));
 sg13g2_dfrbpq_1 _11951_ (.RESET_B(net35),
    .D(_00382_),
    .Q(\mac_inst.get_mac[22] ),
    .CLK(clknet_leaf_49_clk));
 sg13g2_dfrbpq_1 _11952_ (.RESET_B(net259),
    .D(net667),
    .Q(\mac_inst.get_mac[23] ),
    .CLK(clknet_leaf_47_clk));
 sg13g2_dfrbpq_1 _11953_ (.RESET_B(net243),
    .D(net279),
    .Q(\mac_inst.RDY_get_multiply ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 _11954_ (.RESET_B(net227),
    .D(net275),
    .Q(\mac_inst.RDY_get_msu ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 _11955_ (.RESET_B(net211),
    .D(net277),
    .Q(\mac_inst.RDY_get_mac ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_2 _11956_ (.RESET_B(net195),
    .D(net734),
    .Q(\mac_inst.accumulator[0] ),
    .CLK(clknet_leaf_51_clk));
 sg13g2_dfrbpq_2 _11957_ (.RESET_B(net179),
    .D(_00388_),
    .Q(\mac_inst.accumulator[1] ),
    .CLK(clknet_leaf_55_clk));
 sg13g2_dfrbpq_2 _11958_ (.RESET_B(net162),
    .D(_00389_),
    .Q(\mac_inst.accumulator[2] ),
    .CLK(clknet_leaf_55_clk));
 sg13g2_dfrbpq_2 _11959_ (.RESET_B(net146),
    .D(_00390_),
    .Q(\mac_inst.accumulator[3] ),
    .CLK(clknet_leaf_54_clk));
 sg13g2_dfrbpq_1 _11960_ (.RESET_B(net130),
    .D(_00391_),
    .Q(\mac_inst.accumulator[4] ),
    .CLK(clknet_leaf_54_clk));
 sg13g2_dfrbpq_2 _11961_ (.RESET_B(net114),
    .D(_00392_),
    .Q(\mac_inst.accumulator[5] ),
    .CLK(clknet_leaf_60_clk));
 sg13g2_dfrbpq_1 _11962_ (.RESET_B(net99),
    .D(_00393_),
    .Q(\mac_inst.accumulator[6] ),
    .CLK(clknet_leaf_60_clk));
 sg13g2_dfrbpq_2 _11963_ (.RESET_B(net79),
    .D(_00394_),
    .Q(\mac_inst.accumulator[7] ),
    .CLK(clknet_leaf_65_clk));
 sg13g2_dfrbpq_2 _11964_ (.RESET_B(net63),
    .D(_00395_),
    .Q(\mac_inst.accumulator[8] ),
    .CLK(clknet_leaf_64_clk));
 sg13g2_dfrbpq_1 _11965_ (.RESET_B(net48),
    .D(_00396_),
    .Q(\mac_inst.accumulator[9] ),
    .CLK(clknet_leaf_67_clk));
 sg13g2_dfrbpq_2 _11966_ (.RESET_B(net31),
    .D(_00397_),
    .Q(\mac_inst.accumulator[10] ),
    .CLK(clknet_leaf_63_clk));
 sg13g2_dfrbpq_2 _11967_ (.RESET_B(net235),
    .D(_00398_),
    .Q(\mac_inst.accumulator[11] ),
    .CLK(clknet_leaf_63_clk));
 sg13g2_dfrbpq_1 _11968_ (.RESET_B(net203),
    .D(_00399_),
    .Q(\mac_inst.accumulator[12] ),
    .CLK(clknet_leaf_62_clk));
 sg13g2_dfrbpq_2 _11969_ (.RESET_B(net171),
    .D(_00400_),
    .Q(\mac_inst.accumulator[13] ),
    .CLK(clknet_leaf_62_clk));
 sg13g2_dfrbpq_2 _11970_ (.RESET_B(net138),
    .D(_00401_),
    .Q(\mac_inst.accumulator[14] ),
    .CLK(clknet_leaf_53_clk));
 sg13g2_dfrbpq_2 _11971_ (.RESET_B(net106),
    .D(net748),
    .Q(\mac_inst.accumulator[15] ),
    .CLK(clknet_leaf_53_clk));
 sg13g2_dfrbpq_2 _11972_ (.RESET_B(net71),
    .D(_00403_),
    .Q(\mac_inst.accumulator[16] ),
    .CLK(clknet_leaf_52_clk));
 sg13g2_dfrbpq_2 _11973_ (.RESET_B(net39),
    .D(_00404_),
    .Q(\mac_inst.accumulator[17] ),
    .CLK(clknet_leaf_49_clk));
 sg13g2_dfrbpq_1 _11974_ (.RESET_B(net219),
    .D(_00405_),
    .Q(\mac_inst.accumulator[18] ),
    .CLK(clknet_leaf_49_clk));
 sg13g2_dfrbpq_2 _11975_ (.RESET_B(net154),
    .D(net714),
    .Q(\mac_inst.accumulator[19] ),
    .CLK(clknet_leaf_49_clk));
 sg13g2_dfrbpq_2 _11976_ (.RESET_B(net87),
    .D(_00407_),
    .Q(\mac_inst.accumulator[20] ),
    .CLK(clknet_leaf_48_clk));
 sg13g2_dfrbpq_1 _11977_ (.RESET_B(net251),
    .D(_00408_),
    .Q(\mac_inst.accumulator[21] ),
    .CLK(clknet_leaf_48_clk));
 sg13g2_dfrbpq_2 _11978_ (.RESET_B(net122),
    .D(_00409_),
    .Q(\mac_inst.accumulator[22] ),
    .CLK(clknet_leaf_50_clk));
 sg13g2_dfrbpq_1 _11979_ (.RESET_B(net187),
    .D(net652),
    .Q(\mac_inst.accumulator[23] ),
    .CLK(clknet_leaf_47_clk));
 sg13g2_tiehi _11570__28 (.L_HI(net28));
 sg13g2_tiehi _11571__29 (.L_HI(net29));
 sg13g2_tiehi _11572__30 (.L_HI(net30));
 sg13g2_tiehi _11966__31 (.L_HI(net31));
 sg13g2_tiehi _11864__32 (.L_HI(net32));
 sg13g2_tiehi _11922__33 (.L_HI(net33));
 sg13g2_tiehi _11863__34 (.L_HI(net34));
 sg13g2_tiehi _11951__35 (.L_HI(net35));
 sg13g2_tiehi _11862__36 (.L_HI(net36));
 sg13g2_tiehi _11921__37 (.L_HI(net37));
 sg13g2_tiehi _11861__38 (.L_HI(net38));
 sg13g2_tiehi _11973__39 (.L_HI(net39));
 sg13g2_tiehi _11860__40 (.L_HI(net40));
 sg13g2_tiehi _11920__41 (.L_HI(net41));
 sg13g2_tiehi _11859__42 (.L_HI(net42));
 sg13g2_tiehi _11573__43 (.L_HI(net43));
 sg13g2_tiehi _11950__44 (.L_HI(net44));
 sg13g2_tiehi _11858__45 (.L_HI(net45));
 sg13g2_tiehi _11919__46 (.L_HI(net46));
 sg13g2_tiehi _11857__47 (.L_HI(net47));
 sg13g2_tiehi _11965__48 (.L_HI(net48));
 sg13g2_tiehi _11856__49 (.L_HI(net49));
 sg13g2_tiehi _11918__50 (.L_HI(net50));
 sg13g2_tiehi _11855__51 (.L_HI(net51));
 sg13g2_tiehi _11949__52 (.L_HI(net52));
 sg13g2_tiehi _11854__53 (.L_HI(net53));
 sg13g2_tiehi _11917__54 (.L_HI(net54));
 sg13g2_tiehi _11853__55 (.L_HI(net55));
 sg13g2_tiehi _11852__56 (.L_HI(net56));
 sg13g2_tiehi _11916__57 (.L_HI(net57));
 sg13g2_tiehi _11851__58 (.L_HI(net58));
 sg13g2_tiehi _11948__59 (.L_HI(net59));
 sg13g2_tiehi _11850__60 (.L_HI(net60));
 sg13g2_tiehi _11915__61 (.L_HI(net61));
 sg13g2_tiehi _11849__62 (.L_HI(net62));
 sg13g2_tiehi _11964__63 (.L_HI(net63));
 sg13g2_tiehi _11848__64 (.L_HI(net64));
 sg13g2_tiehi _11914__65 (.L_HI(net65));
 sg13g2_tiehi _11847__66 (.L_HI(net66));
 sg13g2_tiehi _11947__67 (.L_HI(net67));
 sg13g2_tiehi _11846__68 (.L_HI(net68));
 sg13g2_tiehi _11913__69 (.L_HI(net69));
 sg13g2_tiehi _11845__70 (.L_HI(net70));
 sg13g2_tiehi _11972__71 (.L_HI(net71));
 sg13g2_tiehi _11844__72 (.L_HI(net72));
 sg13g2_tiehi _11912__73 (.L_HI(net73));
 sg13g2_tiehi _11843__74 (.L_HI(net74));
 sg13g2_tiehi _11946__75 (.L_HI(net75));
 sg13g2_tiehi _11842__76 (.L_HI(net76));
 sg13g2_tiehi _11911__77 (.L_HI(net77));
 sg13g2_tiehi _11841__78 (.L_HI(net78));
 sg13g2_tiehi _11963__79 (.L_HI(net79));
 sg13g2_tiehi _11840__80 (.L_HI(net80));
 sg13g2_tiehi _11910__81 (.L_HI(net81));
 sg13g2_tiehi _11839__82 (.L_HI(net82));
 sg13g2_tiehi _11945__83 (.L_HI(net83));
 sg13g2_tiehi _11838__84 (.L_HI(net84));
 sg13g2_tiehi _11909__85 (.L_HI(net85));
 sg13g2_tiehi _11837__86 (.L_HI(net86));
 sg13g2_tiehi _11976__87 (.L_HI(net87));
 sg13g2_tiehi _11836__88 (.L_HI(net88));
 sg13g2_tiehi _11908__89 (.L_HI(net89));
 sg13g2_tiehi _11835__90 (.L_HI(net90));
 sg13g2_tiehi _11944__91 (.L_HI(net91));
 sg13g2_tiehi _11655__92 (.L_HI(net92));
 sg13g2_tiehi _11656__93 (.L_HI(net93));
 sg13g2_tiehi _11657__94 (.L_HI(net94));
 sg13g2_tiehi _11658__95 (.L_HI(net95));
 sg13g2_tiehi _11834__96 (.L_HI(net96));
 sg13g2_tiehi _11907__97 (.L_HI(net97));
 sg13g2_tiehi _11833__98 (.L_HI(net98));
 sg13g2_tiehi _11962__99 (.L_HI(net99));
 sg13g2_tiehi _11832__100 (.L_HI(net100));
 sg13g2_tiehi _11906__101 (.L_HI(net101));
 sg13g2_tiehi _11831__102 (.L_HI(net102));
 sg13g2_tiehi _11943__103 (.L_HI(net103));
 sg13g2_tiehi _11830__104 (.L_HI(net104));
 sg13g2_tiehi _11905__105 (.L_HI(net105));
 sg13g2_tiehi _11971__106 (.L_HI(net106));
 sg13g2_tiehi _11826__107 (.L_HI(net107));
 sg13g2_tiehi _11904__108 (.L_HI(net108));
 sg13g2_tiehi _11825__109 (.L_HI(net109));
 sg13g2_tiehi _11942__110 (.L_HI(net110));
 sg13g2_tiehi _11824__111 (.L_HI(net111));
 sg13g2_tiehi _11903__112 (.L_HI(net112));
 sg13g2_tiehi _11823__113 (.L_HI(net113));
 sg13g2_tiehi _11961__114 (.L_HI(net114));
 sg13g2_tiehi _11822__115 (.L_HI(net115));
 sg13g2_tiehi _11902__116 (.L_HI(net116));
 sg13g2_tiehi _11821__117 (.L_HI(net117));
 sg13g2_tiehi _11941__118 (.L_HI(net118));
 sg13g2_tiehi _11820__119 (.L_HI(net119));
 sg13g2_tiehi _11901__120 (.L_HI(net120));
 sg13g2_tiehi _11819__121 (.L_HI(net121));
 sg13g2_tiehi _11978__122 (.L_HI(net122));
 sg13g2_tiehi _11818__123 (.L_HI(net123));
 sg13g2_tiehi _11900__124 (.L_HI(net124));
 sg13g2_tiehi _11817__125 (.L_HI(net125));
 sg13g2_tiehi _11940__126 (.L_HI(net126));
 sg13g2_tiehi _11816__127 (.L_HI(net127));
 sg13g2_tiehi _11899__128 (.L_HI(net128));
 sg13g2_tiehi _11815__129 (.L_HI(net129));
 sg13g2_tiehi _11960__130 (.L_HI(net130));
 sg13g2_tiehi _11814__131 (.L_HI(net131));
 sg13g2_tiehi _11898__132 (.L_HI(net132));
 sg13g2_tiehi _11813__133 (.L_HI(net133));
 sg13g2_tiehi _11939__134 (.L_HI(net134));
 sg13g2_tiehi _11812__135 (.L_HI(net135));
 sg13g2_tiehi _11897__136 (.L_HI(net136));
 sg13g2_tiehi _11811__137 (.L_HI(net137));
 sg13g2_tiehi _11970__138 (.L_HI(net138));
 sg13g2_tiehi _11810__139 (.L_HI(net139));
 sg13g2_tiehi _11896__140 (.L_HI(net140));
 sg13g2_tiehi _11809__141 (.L_HI(net141));
 sg13g2_tiehi _11938__142 (.L_HI(net142));
 sg13g2_tiehi _11808__143 (.L_HI(net143));
 sg13g2_tiehi _11895__144 (.L_HI(net144));
 sg13g2_tiehi _11807__145 (.L_HI(net145));
 sg13g2_tiehi _11959__146 (.L_HI(net146));
 sg13g2_tiehi _11806__147 (.L_HI(net147));
 sg13g2_tiehi _11894__148 (.L_HI(net148));
 sg13g2_tiehi _11805__149 (.L_HI(net149));
 sg13g2_tiehi _11937__150 (.L_HI(net150));
 sg13g2_tiehi _11804__151 (.L_HI(net151));
 sg13g2_tiehi _11893__152 (.L_HI(net152));
 sg13g2_tiehi _11803__153 (.L_HI(net153));
 sg13g2_tiehi _11975__154 (.L_HI(net154));
 sg13g2_tiehi _11802__155 (.L_HI(net155));
 sg13g2_tiehi _11892__156 (.L_HI(net156));
 sg13g2_tiehi _11801__157 (.L_HI(net157));
 sg13g2_tiehi _11936__158 (.L_HI(net158));
 sg13g2_tiehi _11800__159 (.L_HI(net159));
 sg13g2_tiehi _11891__160 (.L_HI(net160));
 sg13g2_tiehi _11799__161 (.L_HI(net161));
 sg13g2_tiehi _11958__162 (.L_HI(net162));
 sg13g2_tiehi _11798__163 (.L_HI(net163));
 sg13g2_tiehi _11659__164 (.L_HI(net164));
 sg13g2_tiehi _11890__165 (.L_HI(net165));
 sg13g2_tiehi _11797__166 (.L_HI(net166));
 sg13g2_tiehi _11935__167 (.L_HI(net167));
 sg13g2_tiehi _11796__168 (.L_HI(net168));
 sg13g2_tiehi _11889__169 (.L_HI(net169));
 sg13g2_tiehi _11795__170 (.L_HI(net170));
 sg13g2_tiehi _11969__171 (.L_HI(net171));
 sg13g2_tiehi _11794__172 (.L_HI(net172));
 sg13g2_tiehi _11888__173 (.L_HI(net173));
 sg13g2_tiehi _11793__174 (.L_HI(net174));
 sg13g2_tiehi _11934__175 (.L_HI(net175));
 sg13g2_tiehi _11792__176 (.L_HI(net176));
 sg13g2_tiehi _11887__177 (.L_HI(net177));
 sg13g2_tiehi _11791__178 (.L_HI(net178));
 sg13g2_tiehi _11957__179 (.L_HI(net179));
 sg13g2_tiehi _11790__180 (.L_HI(net180));
 sg13g2_tiehi _11886__181 (.L_HI(net181));
 sg13g2_tiehi _11789__182 (.L_HI(net182));
 sg13g2_tiehi _11933__183 (.L_HI(net183));
 sg13g2_tiehi _11788__184 (.L_HI(net184));
 sg13g2_tiehi _11885__185 (.L_HI(net185));
 sg13g2_tiehi _11787__186 (.L_HI(net186));
 sg13g2_tiehi _11979__187 (.L_HI(net187));
 sg13g2_tiehi _11786__188 (.L_HI(net188));
 sg13g2_tiehi _11884__189 (.L_HI(net189));
 sg13g2_tiehi _11785__190 (.L_HI(net190));
 sg13g2_tiehi _11932__191 (.L_HI(net191));
 sg13g2_tiehi _11784__192 (.L_HI(net192));
 sg13g2_tiehi _11883__193 (.L_HI(net193));
 sg13g2_tiehi _11783__194 (.L_HI(net194));
 sg13g2_tiehi _11956__195 (.L_HI(net195));
 sg13g2_tiehi _11782__196 (.L_HI(net196));
 sg13g2_tiehi _11882__197 (.L_HI(net197));
 sg13g2_tiehi _11781__198 (.L_HI(net198));
 sg13g2_tiehi _11931__199 (.L_HI(net199));
 sg13g2_tiehi _11780__200 (.L_HI(net200));
 sg13g2_tiehi _11881__201 (.L_HI(net201));
 sg13g2_tiehi _11779__202 (.L_HI(net202));
 sg13g2_tiehi _11968__203 (.L_HI(net203));
 sg13g2_tiehi _11778__204 (.L_HI(net204));
 sg13g2_tiehi _11880__205 (.L_HI(net205));
 sg13g2_tiehi _11777__206 (.L_HI(net206));
 sg13g2_tiehi _11930__207 (.L_HI(net207));
 sg13g2_tiehi _11776__208 (.L_HI(net208));
 sg13g2_tiehi _11879__209 (.L_HI(net209));
 sg13g2_tiehi _11775__210 (.L_HI(net210));
 sg13g2_tiehi _11955__211 (.L_HI(net211));
 sg13g2_tiehi _11774__212 (.L_HI(net212));
 sg13g2_tiehi _11878__213 (.L_HI(net213));
 sg13g2_tiehi _11773__214 (.L_HI(net214));
 sg13g2_tiehi _11929__215 (.L_HI(net215));
 sg13g2_tiehi _11772__216 (.L_HI(net216));
 sg13g2_tiehi _11877__217 (.L_HI(net217));
 sg13g2_tiehi _11771__218 (.L_HI(net218));
 sg13g2_tiehi _11974__219 (.L_HI(net219));
 sg13g2_tiehi _11770__220 (.L_HI(net220));
 sg13g2_tiehi _11876__221 (.L_HI(net221));
 sg13g2_tiehi _11769__222 (.L_HI(net222));
 sg13g2_tiehi _11928__223 (.L_HI(net223));
 sg13g2_tiehi _11768__224 (.L_HI(net224));
 sg13g2_tiehi _11875__225 (.L_HI(net225));
 sg13g2_tiehi _11767__226 (.L_HI(net226));
 sg13g2_tiehi _11954__227 (.L_HI(net227));
 sg13g2_tiehi _11766__228 (.L_HI(net228));
 sg13g2_tiehi _11874__229 (.L_HI(net229));
 sg13g2_tiehi _11765__230 (.L_HI(net230));
 sg13g2_tiehi _11927__231 (.L_HI(net231));
 sg13g2_tiehi _11764__232 (.L_HI(net232));
 sg13g2_tiehi _11873__233 (.L_HI(net233));
 sg13g2_tiehi _11763__234 (.L_HI(net234));
 sg13g2_tiehi _11967__235 (.L_HI(net235));
 sg13g2_tiehi _11762__236 (.L_HI(net236));
 sg13g2_tiehi _11872__237 (.L_HI(net237));
 sg13g2_tiehi _11761__238 (.L_HI(net238));
 sg13g2_tiehi _11926__239 (.L_HI(net239));
 sg13g2_tiehi _11760__240 (.L_HI(net240));
 sg13g2_tiehi _11871__241 (.L_HI(net241));
 sg13g2_tiehi _11759__242 (.L_HI(net242));
 sg13g2_tiehi _11953__243 (.L_HI(net243));
 sg13g2_tiehi _11758__244 (.L_HI(net244));
 sg13g2_tiehi _11870__245 (.L_HI(net245));
 sg13g2_tiehi _11757__246 (.L_HI(net246));
 sg13g2_tiehi _11925__247 (.L_HI(net247));
 sg13g2_tiehi _11756__248 (.L_HI(net248));
 sg13g2_tiehi _11869__249 (.L_HI(net249));
 sg13g2_tiehi _11755__250 (.L_HI(net250));
 sg13g2_tiehi _11977__251 (.L_HI(net251));
 sg13g2_tiehi _11754__252 (.L_HI(net252));
 sg13g2_tiehi _11868__253 (.L_HI(net253));
 sg13g2_tiehi _11753__254 (.L_HI(net254));
 sg13g2_tiehi _11924__255 (.L_HI(net255));
 sg13g2_tiehi _11752__256 (.L_HI(net256));
 sg13g2_tiehi _11867__257 (.L_HI(net257));
 sg13g2_tiehi _11751__258 (.L_HI(net258));
 sg13g2_tiehi _11952__259 (.L_HI(net259));
 sg13g2_tiehi _11750__260 (.L_HI(net260));
 sg13g2_tiehi _11866__261 (.L_HI(net261));
 sg13g2_tiehi _11749__262 (.L_HI(net262));
 sg13g2_tiehi _11923__263 (.L_HI(net263));
 sg13g2_tiehi _11748__264 (.L_HI(net264));
 sg13g2_tiehi _11865__265 (.L_HI(net265));
 sg13g2_tiehi _11747__266 (.L_HI(net266));
 sg13g2_tiehi _11666__267 (.L_HI(net267));
 sg13g2_tiehi _11665__268 (.L_HI(net268));
 sg13g2_tiehi _11664__269 (.L_HI(net269));
 sg13g2_tiehi _11663__270 (.L_HI(net270));
 sg13g2_tiehi _11662__271 (.L_HI(net271));
 sg13g2_tiehi _11661__272 (.L_HI(net272));
 sg13g2_tiehi _11660__273 (.L_HI(net273));
 sg13g2_buf_8 clkbuf_leaf_0_clk (.A(clknet_4_2_0_clk),
    .X(clknet_leaf_0_clk));
 sg13g2_tielo tt_um_herald_12 (.L_LO(net12));
 sg13g2_tielo tt_um_herald_13 (.L_LO(net13));
 sg13g2_tielo tt_um_herald_14 (.L_LO(net14));
 sg13g2_tielo tt_um_herald_15 (.L_LO(net15));
 sg13g2_tielo tt_um_herald_16 (.L_LO(net16));
 sg13g2_tielo tt_um_herald_17 (.L_LO(net17));
 sg13g2_tielo tt_um_herald_18 (.L_LO(net18));
 sg13g2_tielo tt_um_herald_19 (.L_LO(net19));
 sg13g2_tielo tt_um_herald_20 (.L_LO(net20));
 sg13g2_tielo tt_um_herald_21 (.L_LO(net21));
 sg13g2_tielo tt_um_herald_22 (.L_LO(net22));
 sg13g2_tielo tt_um_herald_23 (.L_LO(net23));
 sg13g2_tielo tt_um_herald_24 (.L_LO(net24));
 sg13g2_tielo tt_um_herald_25 (.L_LO(net25));
 sg13g2_tielo tt_um_herald_26 (.L_LO(net26));
 sg13g2_tiehi _11574__27 (.L_HI(net27));
 PRAWNS_ART prawns_art_inst ();
 sg13g2_buf_8 fanout1200 (.A(_05280_),
    .X(net1200));
 sg13g2_buf_2 fanout1201 (.A(_05224_),
    .X(net1201));
 sg13g2_buf_8 fanout1202 (.A(_01058_),
    .X(net1202));
 sg13g2_buf_8 fanout1203 (.A(net1204),
    .X(net1203));
 sg13g2_buf_8 fanout1204 (.A(_00773_),
    .X(net1204));
 sg13g2_buf_8 fanout1205 (.A(net1206),
    .X(net1205));
 sg13g2_buf_8 fanout1206 (.A(_00773_),
    .X(net1206));
 sg13g2_buf_8 fanout1207 (.A(net1208),
    .X(net1207));
 sg13g2_buf_1 fanout1208 (.A(net1209),
    .X(net1208));
 sg13g2_buf_8 fanout1209 (.A(_00773_),
    .X(net1209));
 sg13g2_buf_8 fanout1210 (.A(net1211),
    .X(net1210));
 sg13g2_buf_8 fanout1211 (.A(net1215),
    .X(net1211));
 sg13g2_buf_8 fanout1212 (.A(net1213),
    .X(net1212));
 sg13g2_buf_8 fanout1213 (.A(net1215),
    .X(net1213));
 sg13g2_buf_8 fanout1214 (.A(net1215),
    .X(net1214));
 sg13g2_buf_8 fanout1215 (.A(net1226),
    .X(net1215));
 sg13g2_buf_8 fanout1216 (.A(net1217),
    .X(net1216));
 sg13g2_buf_8 fanout1217 (.A(net1218),
    .X(net1217));
 sg13g2_buf_8 fanout1218 (.A(net1226),
    .X(net1218));
 sg13g2_buf_8 fanout1219 (.A(net1223),
    .X(net1219));
 sg13g2_buf_1 fanout1220 (.A(net1223),
    .X(net1220));
 sg13g2_buf_8 fanout1221 (.A(net1223),
    .X(net1221));
 sg13g2_buf_1 fanout1222 (.A(net1223),
    .X(net1222));
 sg13g2_buf_2 fanout1223 (.A(net1226),
    .X(net1223));
 sg13g2_buf_8 fanout1224 (.A(net1225),
    .X(net1224));
 sg13g2_buf_8 fanout1225 (.A(net1226),
    .X(net1225));
 sg13g2_buf_8 fanout1226 (.A(_00559_),
    .X(net1226));
 sg13g2_buf_8 fanout1227 (.A(net1230),
    .X(net1227));
 sg13g2_buf_8 fanout1228 (.A(net1230),
    .X(net1228));
 sg13g2_buf_2 fanout1229 (.A(net1230),
    .X(net1229));
 sg13g2_buf_8 fanout1230 (.A(_00775_),
    .X(net1230));
 sg13g2_buf_8 fanout1231 (.A(_00757_),
    .X(net1231));
 sg13g2_buf_8 fanout1232 (.A(_00757_),
    .X(net1232));
 sg13g2_buf_8 fanout1233 (.A(_00934_),
    .X(net1233));
 sg13g2_buf_2 fanout1234 (.A(_00934_),
    .X(net1234));
 sg13g2_buf_8 fanout1235 (.A(_00933_),
    .X(net1235));
 sg13g2_buf_8 fanout1236 (.A(net1237),
    .X(net1236));
 sg13g2_buf_8 fanout1237 (.A(net1240),
    .X(net1237));
 sg13g2_buf_8 fanout1238 (.A(net1239),
    .X(net1238));
 sg13g2_buf_8 fanout1239 (.A(net1240),
    .X(net1239));
 sg13g2_buf_8 fanout1240 (.A(_00926_),
    .X(net1240));
 sg13g2_buf_8 fanout1241 (.A(net1242),
    .X(net1241));
 sg13g2_buf_8 fanout1242 (.A(net1243),
    .X(net1242));
 sg13g2_buf_2 fanout1243 (.A(_00925_),
    .X(net1243));
 sg13g2_buf_8 fanout1244 (.A(net1246),
    .X(net1244));
 sg13g2_buf_1 fanout1245 (.A(net1246),
    .X(net1245));
 sg13g2_buf_2 fanout1246 (.A(_00925_),
    .X(net1246));
 sg13g2_buf_8 fanout1247 (.A(net1248),
    .X(net1247));
 sg13g2_buf_8 fanout1248 (.A(_00763_),
    .X(net1248));
 sg13g2_buf_8 fanout1249 (.A(net1250),
    .X(net1249));
 sg13g2_buf_8 fanout1250 (.A(_00532_),
    .X(net1250));
 sg13g2_buf_8 fanout1251 (.A(net1252),
    .X(net1251));
 sg13g2_buf_8 fanout1252 (.A(_00454_),
    .X(net1252));
 sg13g2_buf_8 fanout1253 (.A(net1254),
    .X(net1253));
 sg13g2_buf_8 fanout1254 (.A(net1256),
    .X(net1254));
 sg13g2_buf_2 fanout1255 (.A(net1256),
    .X(net1255));
 sg13g2_buf_8 fanout1256 (.A(_00412_),
    .X(net1256));
 sg13g2_buf_8 fanout1257 (.A(net1258),
    .X(net1257));
 sg13g2_buf_8 fanout1258 (.A(net1266),
    .X(net1258));
 sg13g2_buf_8 fanout1259 (.A(net1266),
    .X(net1259));
 sg13g2_buf_1 fanout1260 (.A(net1266),
    .X(net1260));
 sg13g2_buf_8 fanout1261 (.A(net1265),
    .X(net1261));
 sg13g2_buf_8 fanout1262 (.A(net1264),
    .X(net1262));
 sg13g2_buf_1 fanout1263 (.A(net1264),
    .X(net1263));
 sg13g2_buf_8 fanout1264 (.A(net1265),
    .X(net1264));
 sg13g2_buf_8 fanout1265 (.A(net1266),
    .X(net1265));
 sg13g2_buf_8 fanout1266 (.A(_00411_),
    .X(net1266));
 sg13g2_buf_8 fanout1267 (.A(net1268),
    .X(net1267));
 sg13g2_buf_2 fanout1268 (.A(net1271),
    .X(net1268));
 sg13g2_buf_8 fanout1269 (.A(net1271),
    .X(net1269));
 sg13g2_buf_1 fanout1270 (.A(net1271),
    .X(net1270));
 sg13g2_buf_8 fanout1271 (.A(_05636_),
    .X(net1271));
 sg13g2_buf_8 fanout1272 (.A(net1276),
    .X(net1272));
 sg13g2_buf_8 fanout1273 (.A(net1274),
    .X(net1273));
 sg13g2_buf_2 fanout1274 (.A(net1275),
    .X(net1274));
 sg13g2_buf_1 fanout1275 (.A(net1276),
    .X(net1275));
 sg13g2_buf_8 fanout1276 (.A(_05633_),
    .X(net1276));
 sg13g2_buf_8 fanout1277 (.A(_00551_),
    .X(net1277));
 sg13g2_buf_8 fanout1278 (.A(_00546_),
    .X(net1278));
 sg13g2_buf_2 fanout1279 (.A(_00546_),
    .X(net1279));
 sg13g2_buf_8 fanout1280 (.A(_00484_),
    .X(net1280));
 sg13g2_buf_1 fanout1281 (.A(_00484_),
    .X(net1281));
 sg13g2_buf_8 fanout1282 (.A(_00484_),
    .X(net1282));
 sg13g2_buf_8 fanout1283 (.A(net1284),
    .X(net1283));
 sg13g2_buf_8 fanout1284 (.A(_00482_),
    .X(net1284));
 sg13g2_buf_8 fanout1285 (.A(net1286),
    .X(net1285));
 sg13g2_buf_8 fanout1286 (.A(net1292),
    .X(net1286));
 sg13g2_buf_8 fanout1287 (.A(net1292),
    .X(net1287));
 sg13g2_buf_2 fanout1288 (.A(net1292),
    .X(net1288));
 sg13g2_buf_8 fanout1289 (.A(net1291),
    .X(net1289));
 sg13g2_buf_1 fanout1290 (.A(net1291),
    .X(net1290));
 sg13g2_buf_8 fanout1291 (.A(net1292),
    .X(net1291));
 sg13g2_buf_8 fanout1292 (.A(_00481_),
    .X(net1292));
 sg13g2_buf_8 fanout1293 (.A(net1295),
    .X(net1293));
 sg13g2_buf_1 fanout1294 (.A(net1295),
    .X(net1294));
 sg13g2_buf_8 fanout1295 (.A(net1296),
    .X(net1295));
 sg13g2_buf_8 fanout1296 (.A(net1305),
    .X(net1296));
 sg13g2_buf_8 fanout1297 (.A(net1298),
    .X(net1297));
 sg13g2_buf_8 fanout1298 (.A(net1304),
    .X(net1298));
 sg13g2_buf_8 fanout1299 (.A(net1304),
    .X(net1299));
 sg13g2_buf_8 fanout1300 (.A(net1302),
    .X(net1300));
 sg13g2_buf_1 fanout1301 (.A(net1302),
    .X(net1301));
 sg13g2_buf_8 fanout1302 (.A(net1303),
    .X(net1302));
 sg13g2_buf_8 fanout1303 (.A(net1304),
    .X(net1303));
 sg13g2_buf_8 fanout1304 (.A(net1305),
    .X(net1304));
 sg13g2_buf_8 fanout1305 (.A(_00480_),
    .X(net1305));
 sg13g2_buf_8 fanout1306 (.A(_00424_),
    .X(net1306));
 sg13g2_buf_8 fanout1307 (.A(_00419_),
    .X(net1307));
 sg13g2_buf_8 fanout1308 (.A(net1312),
    .X(net1308));
 sg13g2_buf_8 fanout1309 (.A(net1310),
    .X(net1309));
 sg13g2_buf_1 fanout1310 (.A(net1311),
    .X(net1310));
 sg13g2_buf_1 fanout1311 (.A(net1312),
    .X(net1311));
 sg13g2_buf_2 fanout1312 (.A(net1313),
    .X(net1312));
 sg13g2_buf_8 fanout1313 (.A(_05639_),
    .X(net1313));
 sg13g2_buf_8 fanout1314 (.A(net1315),
    .X(net1314));
 sg13g2_buf_2 fanout1315 (.A(net1318),
    .X(net1315));
 sg13g2_buf_8 fanout1316 (.A(net1318),
    .X(net1316));
 sg13g2_buf_1 fanout1317 (.A(net1318),
    .X(net1317));
 sg13g2_buf_8 fanout1318 (.A(_05606_),
    .X(net1318));
 sg13g2_buf_8 fanout1319 (.A(_05364_),
    .X(net1319));
 sg13g2_buf_8 fanout1320 (.A(_00531_),
    .X(net1320));
 sg13g2_buf_8 fanout1321 (.A(_00476_),
    .X(net1321));
 sg13g2_buf_8 fanout1322 (.A(_00476_),
    .X(net1322));
 sg13g2_buf_8 fanout1323 (.A(net1324),
    .X(net1323));
 sg13g2_buf_8 fanout1324 (.A(_00464_),
    .X(net1324));
 sg13g2_buf_8 fanout1325 (.A(_00421_),
    .X(net1325));
 sg13g2_buf_8 fanout1326 (.A(_05627_),
    .X(net1326));
 sg13g2_buf_1 fanout1327 (.A(_05627_),
    .X(net1327));
 sg13g2_buf_8 fanout1328 (.A(_05363_),
    .X(net1328));
 sg13g2_buf_8 fanout1329 (.A(_05363_),
    .X(net1329));
 sg13g2_buf_8 fanout1330 (.A(net1331),
    .X(net1330));
 sg13g2_buf_8 fanout1331 (.A(net1335),
    .X(net1331));
 sg13g2_buf_1 fanout1332 (.A(net1335),
    .X(net1332));
 sg13g2_buf_8 fanout1333 (.A(net1334),
    .X(net1333));
 sg13g2_buf_8 fanout1334 (.A(net1335),
    .X(net1334));
 sg13g2_buf_8 fanout1335 (.A(_05158_),
    .X(net1335));
 sg13g2_buf_8 fanout1336 (.A(net1337),
    .X(net1336));
 sg13g2_buf_8 fanout1337 (.A(_05158_),
    .X(net1337));
 sg13g2_buf_8 fanout1338 (.A(net1339),
    .X(net1338));
 sg13g2_buf_8 fanout1339 (.A(net1340),
    .X(net1339));
 sg13g2_buf_8 fanout1340 (.A(_05158_),
    .X(net1340));
 sg13g2_buf_8 fanout1341 (.A(_01582_),
    .X(net1341));
 sg13g2_buf_8 fanout1342 (.A(_01142_),
    .X(net1342));
 sg13g2_buf_8 fanout1343 (.A(net1345),
    .X(net1343));
 sg13g2_buf_1 fanout1344 (.A(net1345),
    .X(net1344));
 sg13g2_buf_8 fanout1345 (.A(_00907_),
    .X(net1345));
 sg13g2_buf_8 fanout1346 (.A(_00906_),
    .X(net1346));
 sg13g2_buf_8 fanout1347 (.A(_00545_),
    .X(net1347));
 sg13g2_buf_8 fanout1348 (.A(_00478_),
    .X(net1348));
 sg13g2_buf_8 fanout1349 (.A(_00478_),
    .X(net1349));
 sg13g2_buf_8 fanout1350 (.A(net1351),
    .X(net1350));
 sg13g2_buf_8 fanout1351 (.A(net1358),
    .X(net1351));
 sg13g2_buf_8 fanout1352 (.A(net1358),
    .X(net1352));
 sg13g2_buf_8 fanout1353 (.A(net1357),
    .X(net1353));
 sg13g2_buf_8 fanout1354 (.A(net1355),
    .X(net1354));
 sg13g2_buf_2 fanout1355 (.A(net1356),
    .X(net1355));
 sg13g2_buf_8 fanout1356 (.A(net1357),
    .X(net1356));
 sg13g2_buf_2 fanout1357 (.A(net1358),
    .X(net1357));
 sg13g2_buf_2 fanout1358 (.A(_00474_),
    .X(net1358));
 sg13g2_buf_8 fanout1359 (.A(_00462_),
    .X(net1359));
 sg13g2_buf_8 fanout1360 (.A(net1363),
    .X(net1360));
 sg13g2_buf_8 fanout1361 (.A(net1363),
    .X(net1361));
 sg13g2_buf_1 fanout1362 (.A(net1363),
    .X(net1362));
 sg13g2_buf_8 fanout1363 (.A(_00460_),
    .X(net1363));
 sg13g2_buf_8 fanout1364 (.A(net1365),
    .X(net1364));
 sg13g2_buf_8 fanout1365 (.A(net1369),
    .X(net1365));
 sg13g2_buf_8 fanout1366 (.A(net1367),
    .X(net1366));
 sg13g2_buf_2 fanout1367 (.A(net1369),
    .X(net1367));
 sg13g2_buf_2 fanout1368 (.A(net1369),
    .X(net1368));
 sg13g2_buf_8 fanout1369 (.A(_00460_),
    .X(net1369));
 sg13g2_buf_8 fanout1370 (.A(_00459_),
    .X(net1370));
 sg13g2_buf_8 fanout1371 (.A(net1372),
    .X(net1371));
 sg13g2_buf_8 fanout1372 (.A(_00459_),
    .X(net1372));
 sg13g2_buf_8 fanout1373 (.A(net1374),
    .X(net1373));
 sg13g2_buf_8 fanout1374 (.A(net1381),
    .X(net1374));
 sg13g2_buf_8 fanout1375 (.A(net1381),
    .X(net1375));
 sg13g2_buf_8 fanout1376 (.A(net1380),
    .X(net1376));
 sg13g2_buf_8 fanout1377 (.A(net1378),
    .X(net1377));
 sg13g2_buf_2 fanout1378 (.A(net1379),
    .X(net1378));
 sg13g2_buf_8 fanout1379 (.A(net1380),
    .X(net1379));
 sg13g2_buf_2 fanout1380 (.A(net1381),
    .X(net1380));
 sg13g2_buf_8 fanout1381 (.A(_00458_),
    .X(net1381));
 sg13g2_buf_8 fanout1382 (.A(_05623_),
    .X(net1382));
 sg13g2_buf_8 fanout1383 (.A(net1384),
    .X(net1383));
 sg13g2_buf_8 fanout1384 (.A(_05597_),
    .X(net1384));
 sg13g2_buf_8 fanout1385 (.A(net1386),
    .X(net1385));
 sg13g2_buf_8 fanout1386 (.A(_05591_),
    .X(net1386));
 sg13g2_buf_2 fanout1387 (.A(_05591_),
    .X(net1387));
 sg13g2_buf_8 fanout1388 (.A(net1389),
    .X(net1388));
 sg13g2_buf_8 fanout1389 (.A(_05590_),
    .X(net1389));
 sg13g2_buf_8 fanout1390 (.A(net1391),
    .X(net1390));
 sg13g2_buf_8 fanout1391 (.A(_05589_),
    .X(net1391));
 sg13g2_buf_8 fanout1392 (.A(net1393),
    .X(net1392));
 sg13g2_buf_8 fanout1393 (.A(_05589_),
    .X(net1393));
 sg13g2_buf_8 fanout1394 (.A(net1395),
    .X(net1394));
 sg13g2_buf_8 fanout1395 (.A(net1396),
    .X(net1395));
 sg13g2_buf_8 fanout1396 (.A(net1397),
    .X(net1396));
 sg13g2_buf_2 fanout1397 (.A(_05588_),
    .X(net1397));
 sg13g2_buf_8 fanout1398 (.A(net1402),
    .X(net1398));
 sg13g2_buf_1 fanout1399 (.A(net1402),
    .X(net1399));
 sg13g2_buf_8 fanout1400 (.A(net1402),
    .X(net1400));
 sg13g2_buf_1 fanout1401 (.A(net1402),
    .X(net1401));
 sg13g2_buf_8 fanout1402 (.A(_05539_),
    .X(net1402));
 sg13g2_buf_8 fanout1403 (.A(net1404),
    .X(net1403));
 sg13g2_buf_2 fanout1404 (.A(net1405),
    .X(net1404));
 sg13g2_buf_2 fanout1405 (.A(net801),
    .X(net1405));
 sg13g2_buf_8 fanout1406 (.A(net793),
    .X(net1406));
 sg13g2_buf_8 fanout1407 (.A(net1408),
    .X(net1407));
 sg13g2_buf_1 fanout1408 (.A(net1409),
    .X(net1408));
 sg13g2_buf_1 fanout1409 (.A(net1410),
    .X(net1409));
 sg13g2_buf_8 fanout1410 (.A(net797),
    .X(net1410));
 sg13g2_buf_8 fanout1411 (.A(net818),
    .X(net1411));
 sg13g2_buf_8 fanout1412 (.A(net833),
    .X(net1412));
 sg13g2_buf_8 fanout1413 (.A(\cordic_inst.cordic_state[52] ),
    .X(net1413));
 sg13g2_buf_8 fanout1414 (.A(\cordic_inst.cordic_state[50] ),
    .X(net1414));
 sg13g2_buf_8 fanout1415 (.A(\cordic_inst.cordic_state[48] ),
    .X(net1415));
 sg13g2_buf_8 fanout1416 (.A(net842),
    .X(net1416));
 sg13g2_buf_8 fanout1417 (.A(net817),
    .X(net1417));
 sg13g2_buf_8 fanout1418 (.A(\cordic_inst.cordic_state[45] ),
    .X(net1418));
 sg13g2_buf_8 fanout1419 (.A(net802),
    .X(net1419));
 sg13g2_buf_8 fanout1420 (.A(\cordic_inst.cordic_state[43] ),
    .X(net1420));
 sg13g2_buf_8 fanout1421 (.A(net798),
    .X(net1421));
 sg13g2_buf_8 fanout1422 (.A(\cordic_inst.cordic_state[41] ),
    .X(net1422));
 sg13g2_buf_8 fanout1423 (.A(net828),
    .X(net1423));
 sg13g2_buf_8 fanout1424 (.A(net825),
    .X(net1424));
 sg13g2_buf_8 fanout1425 (.A(\cordic_inst.cordic_state[38] ),
    .X(net1425));
 sg13g2_buf_8 fanout1426 (.A(\cordic_inst.cordic_state[37] ),
    .X(net1426));
 sg13g2_buf_8 fanout1427 (.A(net1434),
    .X(net1427));
 sg13g2_buf_1 fanout1428 (.A(net1434),
    .X(net1428));
 sg13g2_buf_8 fanout1429 (.A(net1430),
    .X(net1429));
 sg13g2_buf_8 fanout1430 (.A(net1434),
    .X(net1430));
 sg13g2_buf_8 fanout1431 (.A(net1432),
    .X(net1431));
 sg13g2_buf_1 fanout1432 (.A(net1434),
    .X(net1432));
 sg13g2_buf_8 fanout1433 (.A(net1434),
    .X(net1433));
 sg13g2_buf_8 fanout1434 (.A(\cordic_inst.cordic_state[7] ),
    .X(net1434));
 sg13g2_buf_8 fanout1435 (.A(net1436),
    .X(net1435));
 sg13g2_buf_8 fanout1436 (.A(net1437),
    .X(net1436));
 sg13g2_buf_8 fanout1437 (.A(net1438),
    .X(net1437));
 sg13g2_buf_8 fanout1438 (.A(net860),
    .X(net1438));
 sg13g2_buf_8 fanout1439 (.A(net1441),
    .X(net1439));
 sg13g2_buf_1 fanout1440 (.A(net1441),
    .X(net1440));
 sg13g2_buf_1 fanout1441 (.A(\cordic_inst.cordic_state[6] ),
    .X(net1441));
 sg13g2_buf_8 fanout1442 (.A(net1443),
    .X(net1442));
 sg13g2_buf_8 fanout1443 (.A(net1445),
    .X(net1443));
 sg13g2_buf_8 fanout1444 (.A(net1445),
    .X(net1444));
 sg13g2_buf_8 fanout1445 (.A(\cordic_inst.cordic_state[5] ),
    .X(net1445));
 sg13g2_buf_8 fanout1446 (.A(net1450),
    .X(net1446));
 sg13g2_buf_8 fanout1447 (.A(net1448),
    .X(net1447));
 sg13g2_buf_8 fanout1448 (.A(net1449),
    .X(net1448));
 sg13g2_buf_8 fanout1449 (.A(net1450),
    .X(net1449));
 sg13g2_buf_8 fanout1450 (.A(\cordic_inst.cordic_state[4] ),
    .X(net1450));
 sg13g2_buf_8 fanout1451 (.A(net1452),
    .X(net1451));
 sg13g2_buf_2 fanout1452 (.A(net1453),
    .X(net1452));
 sg13g2_buf_8 fanout1453 (.A(\cordic_inst.cordic_state[4] ),
    .X(net1453));
 sg13g2_buf_8 fanout1454 (.A(net1456),
    .X(net1454));
 sg13g2_buf_8 fanout1455 (.A(net1456),
    .X(net1455));
 sg13g2_buf_8 fanout1456 (.A(net1457),
    .X(net1456));
 sg13g2_buf_8 fanout1457 (.A(net1463),
    .X(net1457));
 sg13g2_buf_8 fanout1458 (.A(net1463),
    .X(net1458));
 sg13g2_buf_8 fanout1459 (.A(net1460),
    .X(net1459));
 sg13g2_buf_8 fanout1460 (.A(net1463),
    .X(net1460));
 sg13g2_buf_8 fanout1461 (.A(net1462),
    .X(net1461));
 sg13g2_buf_8 fanout1462 (.A(net1463),
    .X(net1462));
 sg13g2_buf_8 fanout1463 (.A(\cordic_inst.cordic_state[3] ),
    .X(net1463));
 sg13g2_buf_8 fanout1464 (.A(net668),
    .X(net1464));
 sg13g2_buf_8 fanout1465 (.A(net813),
    .X(net1465));
 sg13g2_buf_8 fanout1466 (.A(net1468),
    .X(net1466));
 sg13g2_buf_2 fanout1467 (.A(net1468),
    .X(net1467));
 sg13g2_buf_8 fanout1468 (.A(mac_en_msu),
    .X(net1468));
 sg13g2_buf_8 fanout1469 (.A(net1471),
    .X(net1469));
 sg13g2_buf_1 fanout1470 (.A(net1471),
    .X(net1470));
 sg13g2_buf_1 fanout1471 (.A(net1473),
    .X(net1471));
 sg13g2_buf_8 fanout1472 (.A(net1473),
    .X(net1472));
 sg13g2_buf_8 fanout1473 (.A(mac_en_multiply),
    .X(net1473));
 sg13g2_buf_8 fanout1474 (.A(net1479),
    .X(net1474));
 sg13g2_buf_8 fanout1475 (.A(net1478),
    .X(net1475));
 sg13g2_buf_8 fanout1476 (.A(net1478),
    .X(net1476));
 sg13g2_buf_1 fanout1477 (.A(net1478),
    .X(net1477));
 sg13g2_buf_8 fanout1478 (.A(net1479),
    .X(net1478));
 sg13g2_buf_8 fanout1479 (.A(cordic_en_atan2),
    .X(net1479));
 sg13g2_buf_8 fanout1480 (.A(net1481),
    .X(net1480));
 sg13g2_buf_8 fanout1481 (.A(cordic_en_sin_cos),
    .X(net1481));
 sg13g2_buf_8 fanout1482 (.A(net1483),
    .X(net1482));
 sg13g2_buf_2 fanout1483 (.A(net1484),
    .X(net1483));
 sg13g2_buf_1 fanout1484 (.A(cordic_en_sin_cos),
    .X(net1484));
 sg13g2_buf_8 fanout1485 (.A(net1489),
    .X(net1485));
 sg13g2_buf_1 fanout1486 (.A(net1489),
    .X(net1486));
 sg13g2_buf_8 fanout1487 (.A(net1488),
    .X(net1487));
 sg13g2_buf_8 fanout1488 (.A(net1489),
    .X(net1488));
 sg13g2_buf_8 fanout1489 (.A(net792),
    .X(net1489));
 sg13g2_buf_8 fanout1490 (.A(net1491),
    .X(net1490));
 sg13g2_buf_8 fanout1491 (.A(\cordic_inst.MUX_cordic_state$write_1__VAL_1[54] ),
    .X(net1491));
 sg13g2_buf_8 fanout1492 (.A(net837),
    .X(net1492));
 sg13g2_buf_8 fanout1493 (.A(net1495),
    .X(net1493));
 sg13g2_buf_1 fanout1494 (.A(net1495),
    .X(net1494));
 sg13g2_buf_8 fanout1495 (.A(\cordic_inst.MUX_cordic_state$write_1__VAL_1[53] ),
    .X(net1495));
 sg13g2_buf_8 fanout1496 (.A(net835),
    .X(net1496));
 sg13g2_buf_8 fanout1497 (.A(net1499),
    .X(net1497));
 sg13g2_buf_8 fanout1498 (.A(net1499),
    .X(net1498));
 sg13g2_buf_8 fanout1499 (.A(net845),
    .X(net1499));
 sg13g2_buf_8 fanout1500 (.A(net1501),
    .X(net1500));
 sg13g2_buf_8 fanout1501 (.A(net1502),
    .X(net1501));
 sg13g2_buf_8 fanout1502 (.A(net856),
    .X(net1502));
 sg13g2_buf_8 fanout1503 (.A(net1505),
    .X(net1503));
 sg13g2_buf_1 fanout1504 (.A(net1505),
    .X(net1504));
 sg13g2_buf_8 fanout1505 (.A(net1506),
    .X(net1505));
 sg13g2_buf_8 fanout1506 (.A(net848),
    .X(net1506));
 sg13g2_buf_8 fanout1507 (.A(net838),
    .X(net1507));
 sg13g2_buf_8 fanout1508 (.A(net1509),
    .X(net1508));
 sg13g2_buf_8 fanout1509 (.A(\cordic_inst.MUX_cordic_state$write_1__VAL_1[49] ),
    .X(net1509));
 sg13g2_buf_8 fanout1510 (.A(net1512),
    .X(net1510));
 sg13g2_buf_8 fanout1511 (.A(net1512),
    .X(net1511));
 sg13g2_buf_8 fanout1512 (.A(net1513),
    .X(net1512));
 sg13g2_buf_8 fanout1513 (.A(net821),
    .X(net1513));
 sg13g2_buf_8 fanout1514 (.A(net1515),
    .X(net1514));
 sg13g2_buf_8 fanout1515 (.A(net841),
    .X(net1515));
 sg13g2_buf_8 fanout1516 (.A(net1517),
    .X(net1516));
 sg13g2_buf_8 fanout1517 (.A(net1518),
    .X(net1517));
 sg13g2_buf_8 fanout1518 (.A(net861),
    .X(net1518));
 sg13g2_buf_8 fanout1519 (.A(net1524),
    .X(net1519));
 sg13g2_buf_1 fanout1520 (.A(net1524),
    .X(net1520));
 sg13g2_buf_8 fanout1521 (.A(net1524),
    .X(net1521));
 sg13g2_buf_1 fanout1522 (.A(net1524),
    .X(net1522));
 sg13g2_buf_8 fanout1523 (.A(net1524),
    .X(net1523));
 sg13g2_buf_8 fanout1524 (.A(net1525),
    .X(net1524));
 sg13g2_buf_8 fanout1525 (.A(net800),
    .X(net1525));
 sg13g2_buf_8 fanout1526 (.A(net840),
    .X(net1526));
 sg13g2_buf_8 fanout1527 (.A(net1530),
    .X(net1527));
 sg13g2_buf_8 fanout1528 (.A(net1529),
    .X(net1528));
 sg13g2_buf_8 fanout1529 (.A(net1530),
    .X(net1529));
 sg13g2_buf_8 fanout1530 (.A(\cordic_inst.MUX_cordic_state$write_1__VAL_1[61] ),
    .X(net1530));
 sg13g2_buf_8 fanout1531 (.A(net1536),
    .X(net1531));
 sg13g2_buf_8 fanout1532 (.A(net1536),
    .X(net1532));
 sg13g2_buf_8 fanout1533 (.A(net1535),
    .X(net1533));
 sg13g2_buf_1 fanout1534 (.A(net1535),
    .X(net1534));
 sg13g2_buf_1 fanout1535 (.A(net1536),
    .X(net1535));
 sg13g2_buf_8 fanout1536 (.A(net853),
    .X(net1536));
 sg13g2_buf_8 fanout1537 (.A(net1542),
    .X(net1537));
 sg13g2_buf_8 fanout1538 (.A(net1539),
    .X(net1538));
 sg13g2_buf_8 fanout1539 (.A(net1540),
    .X(net1539));
 sg13g2_buf_2 fanout1540 (.A(net1541),
    .X(net1540));
 sg13g2_buf_8 fanout1541 (.A(net1542),
    .X(net1541));
 sg13g2_buf_8 fanout1542 (.A(net536),
    .X(net1542));
 sg13g2_buf_8 fanout1543 (.A(net1544),
    .X(net1543));
 sg13g2_buf_8 fanout1544 (.A(\cordic_inst.MUX_cordic_state$write_1__VAL_1[58] ),
    .X(net1544));
 sg13g2_buf_8 fanout1545 (.A(net1547),
    .X(net1545));
 sg13g2_buf_8 fanout1546 (.A(net1547),
    .X(net1546));
 sg13g2_buf_8 fanout1547 (.A(net1548),
    .X(net1547));
 sg13g2_buf_8 fanout1548 (.A(\cordic_inst.MUX_cordic_state$write_1__VAL_1[58] ),
    .X(net1548));
 sg13g2_buf_8 fanout1549 (.A(net1550),
    .X(net1549));
 sg13g2_buf_8 fanout1550 (.A(net811),
    .X(net1550));
 sg13g2_buf_8 fanout1551 (.A(net1552),
    .X(net1551));
 sg13g2_buf_2 fanout1552 (.A(net1553),
    .X(net1552));
 sg13g2_buf_8 fanout1553 (.A(net1554),
    .X(net1553));
 sg13g2_buf_8 fanout1554 (.A(\cordic_inst.MUX_cordic_state$write_1__VAL_1[57] ),
    .X(net1554));
 sg13g2_buf_8 fanout1555 (.A(net1556),
    .X(net1555));
 sg13g2_buf_8 fanout1556 (.A(net1558),
    .X(net1556));
 sg13g2_buf_8 fanout1557 (.A(net1558),
    .X(net1557));
 sg13g2_buf_8 fanout1558 (.A(net1559),
    .X(net1558));
 sg13g2_buf_8 fanout1559 (.A(net463),
    .X(net1559));
 sg13g2_buf_8 fanout1560 (.A(net693),
    .X(net1560));
 sg13g2_buf_8 fanout1561 (.A(net804),
    .X(net1561));
 sg13g2_buf_8 fanout1562 (.A(net1565),
    .X(net1562));
 sg13g2_buf_8 fanout1563 (.A(net1564),
    .X(net1563));
 sg13g2_buf_8 fanout1564 (.A(net1565),
    .X(net1564));
 sg13g2_buf_8 fanout1565 (.A(net852),
    .X(net1565));
 sg13g2_buf_8 fanout1566 (.A(net1567),
    .X(net1566));
 sg13g2_buf_8 fanout1567 (.A(net1568),
    .X(net1567));
 sg13g2_buf_8 fanout1568 (.A(net1569),
    .X(net1568));
 sg13g2_buf_8 fanout1569 (.A(net815),
    .X(net1569));
 sg13g2_buf_8 fanout1570 (.A(net1571),
    .X(net1570));
 sg13g2_buf_8 fanout1571 (.A(net1573),
    .X(net1571));
 sg13g2_buf_8 fanout1572 (.A(net1573),
    .X(net1572));
 sg13g2_buf_8 fanout1573 (.A(net858),
    .X(net1573));
 sg13g2_buf_8 fanout1574 (.A(net1575),
    .X(net1574));
 sg13g2_buf_8 fanout1575 (.A(net1577),
    .X(net1575));
 sg13g2_buf_8 fanout1576 (.A(net1578),
    .X(net1576));
 sg13g2_buf_8 fanout1577 (.A(net1578),
    .X(net1577));
 sg13g2_buf_8 fanout1578 (.A(net854),
    .X(net1578));
 sg13g2_buf_8 fanout1579 (.A(net1582),
    .X(net1579));
 sg13g2_buf_8 fanout1580 (.A(net1581),
    .X(net1580));
 sg13g2_buf_8 fanout1581 (.A(net1582),
    .X(net1581));
 sg13g2_buf_8 fanout1582 (.A(net1583),
    .X(net1582));
 sg13g2_buf_8 fanout1583 (.A(net846),
    .X(net1583));
 sg13g2_buf_8 fanout1584 (.A(net1589),
    .X(net1584));
 sg13g2_buf_8 fanout1585 (.A(net1586),
    .X(net1585));
 sg13g2_buf_1 fanout1586 (.A(net1589),
    .X(net1586));
 sg13g2_buf_8 fanout1587 (.A(net1589),
    .X(net1587));
 sg13g2_buf_1 fanout1588 (.A(net1589),
    .X(net1588));
 sg13g2_buf_8 fanout1589 (.A(net1590),
    .X(net1589));
 sg13g2_buf_8 fanout1590 (.A(net849),
    .X(net1590));
 sg13g2_buf_8 fanout1591 (.A(net1596),
    .X(net1591));
 sg13g2_buf_8 fanout1592 (.A(net1593),
    .X(net1592));
 sg13g2_buf_1 fanout1593 (.A(net1596),
    .X(net1593));
 sg13g2_buf_8 fanout1594 (.A(net1596),
    .X(net1594));
 sg13g2_buf_1 fanout1595 (.A(net1596),
    .X(net1595));
 sg13g2_buf_8 fanout1596 (.A(net1597),
    .X(net1596));
 sg13g2_buf_8 fanout1597 (.A(net850),
    .X(net1597));
 sg13g2_buf_8 fanout1598 (.A(net1600),
    .X(net1598));
 sg13g2_buf_8 fanout1599 (.A(net1600),
    .X(net1599));
 sg13g2_buf_8 fanout1600 (.A(net1601),
    .X(net1600));
 sg13g2_buf_8 fanout1601 (.A(net1602),
    .X(net1601));
 sg13g2_buf_8 fanout1602 (.A(net851),
    .X(net1602));
 sg13g2_buf_8 fanout1603 (.A(net1605),
    .X(net1603));
 sg13g2_buf_8 fanout1604 (.A(net1605),
    .X(net1604));
 sg13g2_buf_8 fanout1605 (.A(net1606),
    .X(net1605));
 sg13g2_buf_8 fanout1606 (.A(net822),
    .X(net1606));
 sg13g2_buf_8 fanout1607 (.A(net1608),
    .X(net1607));
 sg13g2_buf_8 fanout1608 (.A(net1611),
    .X(net1608));
 sg13g2_buf_8 fanout1609 (.A(net1610),
    .X(net1609));
 sg13g2_buf_8 fanout1610 (.A(net1611),
    .X(net1610));
 sg13g2_buf_8 fanout1611 (.A(net809),
    .X(net1611));
 sg13g2_buf_8 fanout1612 (.A(net1614),
    .X(net1612));
 sg13g2_buf_8 fanout1613 (.A(net1614),
    .X(net1613));
 sg13g2_buf_8 fanout1614 (.A(net1615),
    .X(net1614));
 sg13g2_buf_8 fanout1615 (.A(net808),
    .X(net1615));
 sg13g2_buf_8 fanout1616 (.A(net1622),
    .X(net1616));
 sg13g2_buf_1 fanout1617 (.A(net1622),
    .X(net1617));
 sg13g2_buf_8 fanout1618 (.A(net1619),
    .X(net1618));
 sg13g2_buf_8 fanout1619 (.A(net1622),
    .X(net1619));
 sg13g2_buf_8 fanout1620 (.A(net1621),
    .X(net1620));
 sg13g2_buf_2 fanout1621 (.A(net1622),
    .X(net1621));
 sg13g2_buf_8 fanout1622 (.A(net857),
    .X(net1622));
 sg13g2_buf_8 fanout1623 (.A(net1624),
    .X(net1623));
 sg13g2_buf_8 fanout1624 (.A(\cordic_inst.MUX_cordic_state$write_1__VAL_1[35] ),
    .X(net1624));
 sg13g2_buf_8 fanout1625 (.A(net1626),
    .X(net1625));
 sg13g2_buf_8 fanout1626 (.A(\cordic_inst.MUX_cordic_state$write_1__VAL_1[35] ),
    .X(net1626));
 sg13g2_buf_8 fanout1627 (.A(net839),
    .X(net1627));
 sg13g2_buf_8 fanout1628 (.A(net1629),
    .X(net1628));
 sg13g2_buf_8 fanout1629 (.A(net1632),
    .X(net1629));
 sg13g2_buf_8 fanout1630 (.A(net1632),
    .X(net1630));
 sg13g2_buf_8 fanout1631 (.A(net1632),
    .X(net1631));
 sg13g2_buf_8 fanout1632 (.A(net843),
    .X(net1632));
 sg13g2_buf_2 fanout1633 (.A(net1635),
    .X(net1633));
 sg13g2_buf_8 fanout1634 (.A(net1635),
    .X(net1634));
 sg13g2_buf_8 fanout1635 (.A(\cordic_inst.MUX_cordic_state$write_1__VAL_1[33] ),
    .X(net1635));
 sg13g2_buf_2 fanout1636 (.A(net1637),
    .X(net1636));
 sg13g2_buf_1 fanout1637 (.A(net1639),
    .X(net1637));
 sg13g2_buf_2 fanout1638 (.A(net1639),
    .X(net1638));
 sg13g2_buf_8 fanout1639 (.A(\cordic_inst.MUX_cordic_state$write_1__VAL_1[33] ),
    .X(net1639));
 sg13g2_buf_2 fanout1640 (.A(net1641),
    .X(net1640));
 sg13g2_buf_1 fanout1641 (.A(net1642),
    .X(net1641));
 sg13g2_buf_2 fanout1642 (.A(net1643),
    .X(net1642));
 sg13g2_buf_2 fanout1643 (.A(\cordic_inst.MUX_cordic_state$write_1__VAL_1[33] ),
    .X(net1643));
 sg13g2_buf_2 fanout1644 (.A(net1645),
    .X(net1644));
 sg13g2_buf_8 fanout1645 (.A(net1654),
    .X(net1645));
 sg13g2_buf_2 fanout1646 (.A(net1647),
    .X(net1646));
 sg13g2_buf_1 fanout1647 (.A(net1649),
    .X(net1647));
 sg13g2_buf_2 fanout1648 (.A(net1649),
    .X(net1648));
 sg13g2_buf_1 fanout1649 (.A(net1654),
    .X(net1649));
 sg13g2_buf_2 fanout1650 (.A(net1651),
    .X(net1650));
 sg13g2_buf_1 fanout1651 (.A(net1652),
    .X(net1651));
 sg13g2_buf_2 fanout1652 (.A(net1654),
    .X(net1652));
 sg13g2_buf_8 fanout1653 (.A(net1654),
    .X(net1653));
 sg13g2_buf_8 fanout1654 (.A(net859),
    .X(net1654));
 sg13g2_buf_8 fanout1655 (.A(net1656),
    .X(net1655));
 sg13g2_buf_8 fanout1656 (.A(net1657),
    .X(net1656));
 sg13g2_buf_8 fanout1657 (.A(net469),
    .X(net1657));
 sg13g2_buf_8 fanout1658 (.A(net1661),
    .X(net1658));
 sg13g2_buf_1 fanout1659 (.A(net1661),
    .X(net1659));
 sg13g2_buf_8 fanout1660 (.A(net1661),
    .X(net1660));
 sg13g2_buf_8 fanout1661 (.A(net847),
    .X(net1661));
 sg13g2_buf_8 fanout1662 (.A(net1665),
    .X(net1662));
 sg13g2_buf_8 fanout1663 (.A(net1665),
    .X(net1663));
 sg13g2_buf_1 fanout1664 (.A(net1665),
    .X(net1664));
 sg13g2_buf_8 fanout1665 (.A(net482),
    .X(net1665));
 sg13g2_buf_8 fanout1666 (.A(net834),
    .X(net1666));
 sg13g2_buf_1 fanout1667 (.A(\cordic_inst.MUX_cordic_state$write_1__VAL_1[76] ),
    .X(net1667));
 sg13g2_buf_2 fanout1668 (.A(net1669),
    .X(net1668));
 sg13g2_buf_8 fanout1669 (.A(\cordic_inst.MUX_cordic_state$write_1__VAL_1[76] ),
    .X(net1669));
 sg13g2_buf_8 fanout1670 (.A(net831),
    .X(net1670));
 sg13g2_buf_8 fanout1671 (.A(net1673),
    .X(net1671));
 sg13g2_buf_1 fanout1672 (.A(net1673),
    .X(net1672));
 sg13g2_buf_8 fanout1673 (.A(\cordic_inst.MUX_cordic_state$write_1__VAL_1[75] ),
    .X(net1673));
 sg13g2_buf_8 fanout1674 (.A(net1678),
    .X(net1674));
 sg13g2_buf_8 fanout1675 (.A(net1677),
    .X(net1675));
 sg13g2_buf_1 fanout1676 (.A(net1677),
    .X(net1676));
 sg13g2_buf_8 fanout1677 (.A(net1678),
    .X(net1677));
 sg13g2_buf_8 fanout1678 (.A(net844),
    .X(net1678));
 sg13g2_buf_8 fanout1679 (.A(net1683),
    .X(net1679));
 sg13g2_buf_8 fanout1680 (.A(net1681),
    .X(net1680));
 sg13g2_buf_8 fanout1681 (.A(net1682),
    .X(net1681));
 sg13g2_buf_2 fanout1682 (.A(net1683),
    .X(net1682));
 sg13g2_buf_2 fanout1683 (.A(net855),
    .X(net1683));
 sg13g2_buf_8 fanout1684 (.A(net1685),
    .X(net1684));
 sg13g2_buf_8 fanout1685 (.A(net1688),
    .X(net1685));
 sg13g2_buf_8 fanout1686 (.A(net1688),
    .X(net1686));
 sg13g2_buf_8 fanout1687 (.A(net1688),
    .X(net1687));
 sg13g2_buf_8 fanout1688 (.A(\cordic_inst.MUX_cordic_state$write_1__VAL_1[72] ),
    .X(net1688));
 sg13g2_buf_8 fanout1689 (.A(net1690),
    .X(net1689));
 sg13g2_buf_1 fanout1690 (.A(net1691),
    .X(net1690));
 sg13g2_buf_8 fanout1691 (.A(net1692),
    .X(net1691));
 sg13g2_buf_8 fanout1692 (.A(\cordic_inst.MUX_cordic_state$write_1__VAL_1[71] ),
    .X(net1692));
 sg13g2_buf_8 fanout1693 (.A(net401),
    .X(net1693));
 sg13g2_buf_8 fanout1694 (.A(net1695),
    .X(net1694));
 sg13g2_buf_1 fanout1695 (.A(net1697),
    .X(net1695));
 sg13g2_buf_8 fanout1696 (.A(net1697),
    .X(net1696));
 sg13g2_buf_8 fanout1697 (.A(\cordic_inst.MUX_cordic_state$write_1__VAL_1[70] ),
    .X(net1697));
 sg13g2_buf_8 fanout1698 (.A(net832),
    .X(net1698));
 sg13g2_buf_8 fanout1699 (.A(net1700),
    .X(net1699));
 sg13g2_buf_8 fanout1700 (.A(net1703),
    .X(net1700));
 sg13g2_buf_8 fanout1701 (.A(net1703),
    .X(net1701));
 sg13g2_buf_8 fanout1702 (.A(net1703),
    .X(net1702));
 sg13g2_buf_8 fanout1703 (.A(net812),
    .X(net1703));
 sg13g2_buf_8 fanout1704 (.A(net1705),
    .X(net1704));
 sg13g2_buf_8 fanout1705 (.A(net1708),
    .X(net1705));
 sg13g2_buf_2 fanout1706 (.A(net1707),
    .X(net1706));
 sg13g2_buf_8 fanout1707 (.A(net1708),
    .X(net1707));
 sg13g2_buf_8 fanout1708 (.A(net1709),
    .X(net1708));
 sg13g2_buf_8 fanout1709 (.A(net795),
    .X(net1709));
 sg13g2_buf_8 fanout1710 (.A(net1711),
    .X(net1710));
 sg13g2_buf_8 fanout1711 (.A(net1714),
    .X(net1711));
 sg13g2_buf_2 fanout1712 (.A(net1713),
    .X(net1712));
 sg13g2_buf_8 fanout1713 (.A(net1714),
    .X(net1713));
 sg13g2_buf_8 fanout1714 (.A(net816),
    .X(net1714));
 sg13g2_buf_8 fanout1715 (.A(net1716),
    .X(net1715));
 sg13g2_buf_8 fanout1716 (.A(net1719),
    .X(net1716));
 sg13g2_buf_8 fanout1717 (.A(net1718),
    .X(net1717));
 sg13g2_buf_8 fanout1718 (.A(net1719),
    .X(net1718));
 sg13g2_buf_8 fanout1719 (.A(net1720),
    .X(net1719));
 sg13g2_buf_8 fanout1720 (.A(net807),
    .X(net1720));
 sg13g2_buf_8 fanout1721 (.A(net1722),
    .X(net1721));
 sg13g2_buf_8 fanout1722 (.A(net1726),
    .X(net1722));
 sg13g2_buf_8 fanout1723 (.A(net1725),
    .X(net1723));
 sg13g2_buf_1 fanout1724 (.A(net1725),
    .X(net1724));
 sg13g2_buf_8 fanout1725 (.A(net1726),
    .X(net1725));
 sg13g2_buf_8 fanout1726 (.A(net1727),
    .X(net1726));
 sg13g2_buf_8 fanout1727 (.A(net428),
    .X(net1727));
 sg13g2_buf_8 fanout1728 (.A(net1729),
    .X(net1728));
 sg13g2_buf_8 fanout1729 (.A(net1733),
    .X(net1729));
 sg13g2_buf_8 fanout1730 (.A(net1731),
    .X(net1730));
 sg13g2_buf_8 fanout1731 (.A(net1732),
    .X(net1731));
 sg13g2_buf_8 fanout1732 (.A(net1733),
    .X(net1732));
 sg13g2_buf_8 fanout1733 (.A(net823),
    .X(net1733));
 sg13g2_buf_8 fanout1734 (.A(net1735),
    .X(net1734));
 sg13g2_buf_8 fanout1735 (.A(net1745),
    .X(net1735));
 sg13g2_buf_8 fanout1736 (.A(net1745),
    .X(net1736));
 sg13g2_buf_8 fanout1737 (.A(net1745),
    .X(net1737));
 sg13g2_buf_8 fanout1738 (.A(net1739),
    .X(net1738));
 sg13g2_buf_8 fanout1739 (.A(net1742),
    .X(net1739));
 sg13g2_buf_8 fanout1740 (.A(net1741),
    .X(net1740));
 sg13g2_buf_8 fanout1741 (.A(net1742),
    .X(net1741));
 sg13g2_buf_8 fanout1742 (.A(net1745),
    .X(net1742));
 sg13g2_buf_8 fanout1743 (.A(net1744),
    .X(net1743));
 sg13g2_buf_8 fanout1744 (.A(net1745),
    .X(net1744));
 sg13g2_buf_8 fanout1745 (.A(net1750),
    .X(net1745));
 sg13g2_buf_8 fanout1746 (.A(net1747),
    .X(net1746));
 sg13g2_buf_8 fanout1747 (.A(net1750),
    .X(net1747));
 sg13g2_buf_8 fanout1748 (.A(net1750),
    .X(net1748));
 sg13g2_buf_1 fanout1749 (.A(net1750),
    .X(net1749));
 sg13g2_buf_8 fanout1750 (.A(_05593_),
    .X(net1750));
 sg13g2_buf_8 fanout1751 (.A(net1753),
    .X(net1751));
 sg13g2_buf_1 fanout1752 (.A(net1753),
    .X(net1752));
 sg13g2_buf_8 fanout1753 (.A(net1764),
    .X(net1753));
 sg13g2_buf_8 fanout1754 (.A(net1756),
    .X(net1754));
 sg13g2_buf_8 fanout1755 (.A(net1756),
    .X(net1755));
 sg13g2_buf_8 fanout1756 (.A(net1764),
    .X(net1756));
 sg13g2_buf_8 fanout1757 (.A(net1760),
    .X(net1757));
 sg13g2_buf_1 fanout1758 (.A(net1760),
    .X(net1758));
 sg13g2_buf_8 fanout1759 (.A(net1760),
    .X(net1759));
 sg13g2_buf_8 fanout1760 (.A(net1764),
    .X(net1760));
 sg13g2_buf_8 fanout1761 (.A(net1762),
    .X(net1761));
 sg13g2_buf_8 fanout1762 (.A(net1763),
    .X(net1762));
 sg13g2_buf_8 fanout1763 (.A(net1764),
    .X(net1763));
 sg13g2_buf_8 fanout1764 (.A(rst_n),
    .X(net1764));
 sg13g2_buf_8 fanout1765 (.A(net1794),
    .X(net1765));
 sg13g2_buf_8 fanout1766 (.A(net1794),
    .X(net1766));
 sg13g2_buf_8 fanout1767 (.A(net1771),
    .X(net1767));
 sg13g2_buf_1 fanout1768 (.A(net1771),
    .X(net1768));
 sg13g2_buf_8 fanout1769 (.A(net1770),
    .X(net1769));
 sg13g2_buf_8 fanout1770 (.A(net1771),
    .X(net1770));
 sg13g2_buf_8 fanout1771 (.A(net1777),
    .X(net1771));
 sg13g2_buf_8 fanout1772 (.A(net1773),
    .X(net1772));
 sg13g2_buf_8 fanout1773 (.A(net1777),
    .X(net1773));
 sg13g2_buf_8 fanout1774 (.A(net1775),
    .X(net1774));
 sg13g2_buf_8 fanout1775 (.A(net1776),
    .X(net1775));
 sg13g2_buf_8 fanout1776 (.A(net1777),
    .X(net1776));
 sg13g2_buf_8 fanout1777 (.A(net1794),
    .X(net1777));
 sg13g2_buf_8 fanout1778 (.A(net1779),
    .X(net1778));
 sg13g2_buf_8 fanout1779 (.A(net1780),
    .X(net1779));
 sg13g2_buf_8 fanout1780 (.A(net1793),
    .X(net1780));
 sg13g2_buf_8 fanout1781 (.A(net1782),
    .X(net1781));
 sg13g2_buf_8 fanout1782 (.A(net1783),
    .X(net1782));
 sg13g2_buf_8 fanout1783 (.A(net1793),
    .X(net1783));
 sg13g2_buf_8 fanout1784 (.A(net1789),
    .X(net1784));
 sg13g2_buf_1 fanout1785 (.A(net1786),
    .X(net1785));
 sg13g2_buf_8 fanout1786 (.A(net1789),
    .X(net1786));
 sg13g2_buf_8 fanout1787 (.A(net1789),
    .X(net1787));
 sg13g2_buf_2 fanout1788 (.A(net1789),
    .X(net1788));
 sg13g2_buf_8 fanout1789 (.A(net1793),
    .X(net1789));
 sg13g2_buf_8 fanout1790 (.A(net1791),
    .X(net1790));
 sg13g2_buf_8 fanout1791 (.A(net1792),
    .X(net1791));
 sg13g2_buf_8 fanout1792 (.A(net1793),
    .X(net1792));
 sg13g2_buf_8 fanout1793 (.A(net1794),
    .X(net1793));
 sg13g2_buf_8 fanout1794 (.A(rst_n),
    .X(net1794));
 sg13g2_buf_2 input1 (.A(ui_in[0]),
    .X(net1));
 sg13g2_buf_2 input2 (.A(ui_in[1]),
    .X(net2));
 sg13g2_buf_2 input3 (.A(ui_in[2]),
    .X(net3));
 sg13g2_buf_2 input4 (.A(ui_in[3]),
    .X(net4));
 sg13g2_buf_2 input5 (.A(ui_in[4]),
    .X(net5));
 sg13g2_buf_2 input6 (.A(ui_in[5]),
    .X(net6));
 sg13g2_buf_2 input7 (.A(ui_in[6]),
    .X(net7));
 sg13g2_buf_2 input8 (.A(ui_in[7]),
    .X(net8));
 sg13g2_buf_1 input9 (.A(uio_in[0]),
    .X(net9));
 sg13g2_buf_1 input10 (.A(uio_in[1]),
    .X(net10));
 sg13g2_tielo tt_um_herald_11 (.L_LO(net11));
 sg13g2_buf_8 clkbuf_leaf_1_clk (.A(clknet_4_2_0_clk),
    .X(clknet_leaf_1_clk));
 sg13g2_buf_8 clkbuf_leaf_2_clk (.A(clknet_4_2_0_clk),
    .X(clknet_leaf_2_clk));
 sg13g2_buf_8 clkbuf_leaf_3_clk (.A(clknet_4_2_0_clk),
    .X(clknet_leaf_3_clk));
 sg13g2_buf_8 clkbuf_leaf_4_clk (.A(clknet_4_3_0_clk),
    .X(clknet_leaf_4_clk));
 sg13g2_buf_8 clkbuf_leaf_7_clk (.A(clknet_4_8_0_clk),
    .X(clknet_leaf_7_clk));
 sg13g2_buf_8 clkbuf_leaf_8_clk (.A(clknet_4_8_0_clk),
    .X(clknet_leaf_8_clk));
 sg13g2_buf_8 clkbuf_leaf_9_clk (.A(clknet_4_8_0_clk),
    .X(clknet_leaf_9_clk));
 sg13g2_buf_8 clkbuf_leaf_10_clk (.A(clknet_4_10_0_clk),
    .X(clknet_leaf_10_clk));
 sg13g2_buf_8 clkbuf_leaf_11_clk (.A(clknet_4_10_0_clk),
    .X(clknet_leaf_11_clk));
 sg13g2_buf_8 clkbuf_leaf_12_clk (.A(clknet_4_10_0_clk),
    .X(clknet_leaf_12_clk));
 sg13g2_buf_8 clkbuf_leaf_13_clk (.A(clknet_4_11_0_clk),
    .X(clknet_leaf_13_clk));
 sg13g2_buf_8 clkbuf_leaf_14_clk (.A(clknet_4_10_0_clk),
    .X(clknet_leaf_14_clk));
 sg13g2_buf_8 clkbuf_leaf_15_clk (.A(clknet_4_9_0_clk),
    .X(clknet_leaf_15_clk));
 sg13g2_buf_8 clkbuf_leaf_16_clk (.A(clknet_4_11_0_clk),
    .X(clknet_leaf_16_clk));
 sg13g2_buf_8 clkbuf_leaf_17_clk (.A(clknet_4_11_0_clk),
    .X(clknet_leaf_17_clk));
 sg13g2_buf_8 clkbuf_leaf_18_clk (.A(clknet_4_11_0_clk),
    .X(clknet_leaf_18_clk));
 sg13g2_buf_8 clkbuf_leaf_19_clk (.A(clknet_4_9_0_clk),
    .X(clknet_leaf_19_clk));
 sg13g2_buf_8 clkbuf_leaf_20_clk (.A(clknet_4_9_0_clk),
    .X(clknet_leaf_20_clk));
 sg13g2_buf_8 clkbuf_leaf_21_clk (.A(clknet_4_8_0_clk),
    .X(clknet_leaf_21_clk));
 sg13g2_buf_8 clkbuf_leaf_22_clk (.A(clknet_4_3_0_clk),
    .X(clknet_leaf_22_clk));
 sg13g2_buf_8 clkbuf_leaf_23_clk (.A(clknet_4_6_0_clk),
    .X(clknet_leaf_23_clk));
 sg13g2_buf_8 clkbuf_leaf_24_clk (.A(clknet_4_12_0_clk),
    .X(clknet_leaf_24_clk));
 sg13g2_buf_8 clkbuf_leaf_25_clk (.A(clknet_4_12_0_clk),
    .X(clknet_leaf_25_clk));
 sg13g2_buf_8 clkbuf_leaf_26_clk (.A(clknet_4_9_0_clk),
    .X(clknet_leaf_26_clk));
 sg13g2_buf_8 clkbuf_leaf_27_clk (.A(clknet_4_14_0_clk),
    .X(clknet_leaf_27_clk));
 sg13g2_buf_8 clkbuf_leaf_28_clk (.A(clknet_4_14_0_clk),
    .X(clknet_leaf_28_clk));
 sg13g2_buf_8 clkbuf_leaf_29_clk (.A(clknet_4_14_0_clk),
    .X(clknet_leaf_29_clk));
 sg13g2_buf_8 clkbuf_leaf_30_clk (.A(clknet_4_14_0_clk),
    .X(clknet_leaf_30_clk));
 sg13g2_buf_8 clkbuf_leaf_31_clk (.A(clknet_4_15_0_clk),
    .X(clknet_leaf_31_clk));
 sg13g2_buf_8 clkbuf_leaf_32_clk (.A(clknet_4_15_0_clk),
    .X(clknet_leaf_32_clk));
 sg13g2_buf_8 clkbuf_leaf_33_clk (.A(clknet_4_15_0_clk),
    .X(clknet_leaf_33_clk));
 sg13g2_buf_8 clkbuf_leaf_34_clk (.A(clknet_4_13_0_clk),
    .X(clknet_leaf_34_clk));
 sg13g2_buf_8 clkbuf_leaf_35_clk (.A(clknet_4_15_0_clk),
    .X(clknet_leaf_35_clk));
 sg13g2_buf_8 clkbuf_leaf_36_clk (.A(clknet_4_12_0_clk),
    .X(clknet_leaf_36_clk));
 sg13g2_buf_8 clkbuf_leaf_37_clk (.A(clknet_4_13_0_clk),
    .X(clknet_leaf_37_clk));
 sg13g2_buf_8 clkbuf_leaf_38_clk (.A(clknet_4_13_0_clk),
    .X(clknet_leaf_38_clk));
 sg13g2_buf_8 clkbuf_leaf_39_clk (.A(clknet_4_13_0_clk),
    .X(clknet_leaf_39_clk));
 sg13g2_buf_8 clkbuf_leaf_40_clk (.A(clknet_4_12_0_clk),
    .X(clknet_leaf_40_clk));
 sg13g2_buf_8 clkbuf_leaf_41_clk (.A(clknet_4_12_0_clk),
    .X(clknet_leaf_41_clk));
 sg13g2_buf_8 clkbuf_leaf_42_clk (.A(clknet_4_7_0_clk),
    .X(clknet_leaf_42_clk));
 sg13g2_buf_8 clkbuf_leaf_43_clk (.A(clknet_4_6_0_clk),
    .X(clknet_leaf_43_clk));
 sg13g2_buf_8 clkbuf_leaf_44_clk (.A(clknet_4_7_0_clk),
    .X(clknet_leaf_44_clk));
 sg13g2_buf_8 clkbuf_leaf_45_clk (.A(clknet_4_7_0_clk),
    .X(clknet_leaf_45_clk));
 sg13g2_buf_8 clkbuf_leaf_46_clk (.A(clknet_4_7_0_clk),
    .X(clknet_leaf_46_clk));
 sg13g2_buf_8 clkbuf_leaf_47_clk (.A(clknet_4_5_0_clk),
    .X(clknet_leaf_47_clk));
 sg13g2_buf_8 clkbuf_leaf_48_clk (.A(clknet_4_5_0_clk),
    .X(clknet_leaf_48_clk));
 sg13g2_buf_8 clkbuf_leaf_49_clk (.A(clknet_4_5_0_clk),
    .X(clknet_leaf_49_clk));
 sg13g2_buf_8 clkbuf_leaf_50_clk (.A(clknet_4_5_0_clk),
    .X(clknet_leaf_50_clk));
 sg13g2_buf_8 clkbuf_leaf_51_clk (.A(clknet_4_4_0_clk),
    .X(clknet_leaf_51_clk));
 sg13g2_buf_8 clkbuf_leaf_52_clk (.A(clknet_4_4_0_clk),
    .X(clknet_leaf_52_clk));
 sg13g2_buf_8 clkbuf_leaf_53_clk (.A(clknet_4_4_0_clk),
    .X(clknet_leaf_53_clk));
 sg13g2_buf_8 clkbuf_leaf_54_clk (.A(clknet_4_4_0_clk),
    .X(clknet_leaf_54_clk));
 sg13g2_buf_8 clkbuf_leaf_55_clk (.A(clknet_4_4_0_clk),
    .X(clknet_leaf_55_clk));
 sg13g2_buf_8 clkbuf_leaf_56_clk (.A(clknet_4_6_0_clk),
    .X(clknet_leaf_56_clk));
 sg13g2_buf_8 clkbuf_leaf_57_clk (.A(clknet_4_6_0_clk),
    .X(clknet_leaf_57_clk));
 sg13g2_buf_8 clkbuf_leaf_58_clk (.A(clknet_4_1_0_clk),
    .X(clknet_leaf_58_clk));
 sg13g2_buf_8 clkbuf_leaf_59_clk (.A(clknet_4_3_0_clk),
    .X(clknet_leaf_59_clk));
 sg13g2_buf_8 clkbuf_leaf_60_clk (.A(clknet_4_1_0_clk),
    .X(clknet_leaf_60_clk));
 sg13g2_buf_8 clkbuf_leaf_61_clk (.A(clknet_4_1_0_clk),
    .X(clknet_leaf_61_clk));
 sg13g2_buf_8 clkbuf_leaf_62_clk (.A(clknet_4_0_0_clk),
    .X(clknet_leaf_62_clk));
 sg13g2_buf_8 clkbuf_leaf_63_clk (.A(clknet_4_0_0_clk),
    .X(clknet_leaf_63_clk));
 sg13g2_buf_8 clkbuf_leaf_64_clk (.A(clknet_4_0_0_clk),
    .X(clknet_leaf_64_clk));
 sg13g2_buf_8 clkbuf_leaf_65_clk (.A(clknet_4_1_0_clk),
    .X(clknet_leaf_65_clk));
 sg13g2_buf_8 clkbuf_leaf_67_clk (.A(clknet_4_0_0_clk),
    .X(clknet_leaf_67_clk));
 sg13g2_buf_8 clkbuf_leaf_68_clk (.A(clknet_4_2_0_clk),
    .X(clknet_leaf_68_clk));
 sg13g2_buf_8 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_buf_8 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sg13g2_buf_8 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sg13g2_buf_8 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sg13g2_buf_8 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sg13g2_buf_8 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sg13g2_buf_8 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sg13g2_buf_8 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sg13g2_buf_8 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sg13g2_buf_8 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sg13g2_buf_8 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sg13g2_buf_8 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sg13g2_buf_8 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sg13g2_buf_8 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sg13g2_buf_8 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sg13g2_buf_8 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sg13g2_buf_8 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sg13g2_inv_2 clkload0 (.A(clknet_4_0_0_clk));
 sg13g2_buf_8 clkload1 (.A(clknet_4_1_0_clk));
 sg13g2_inv_4 clkload2 (.A(clknet_4_3_0_clk));
 sg13g2_buf_8 clkload3 (.A(clknet_4_5_0_clk));
 sg13g2_buf_8 clkload4 (.A(clknet_4_6_0_clk));
 sg13g2_buf_8 clkload5 (.A(clknet_4_7_0_clk));
 sg13g2_inv_2 clkload6 (.A(clknet_4_8_0_clk));
 sg13g2_buf_8 clkload7 (.A(clknet_4_9_0_clk));
 sg13g2_buf_8 clkload8 (.A(clknet_4_10_0_clk));
 sg13g2_buf_8 clkload9 (.A(clknet_4_11_0_clk));
 sg13g2_buf_8 clkload10 (.A(clknet_4_13_0_clk));
 sg13g2_buf_8 clkload11 (.A(clknet_4_14_0_clk));
 sg13g2_buf_8 clkload12 (.A(clknet_4_15_0_clk));
 sg13g2_inv_2 clkload13 (.A(clknet_leaf_64_clk));
 sg13g2_buf_1 clkload14 (.A(clknet_leaf_67_clk));
 sg13g2_buf_8 clkload15 (.A(clknet_leaf_58_clk));
 sg13g2_inv_4 clkload16 (.A(clknet_leaf_60_clk));
 sg13g2_inv_8 clkload17 (.A(clknet_leaf_65_clk));
 sg13g2_inv_8 clkload18 (.A(clknet_leaf_2_clk));
 sg13g2_inv_2 clkload19 (.A(clknet_leaf_3_clk));
 sg13g2_buf_8 clkload20 (.A(clknet_leaf_68_clk));
 sg13g2_inv_2 clkload21 (.A(clknet_leaf_4_clk));
 sg13g2_buf_8 clkload22 (.A(clknet_leaf_59_clk));
 sg13g2_inv_4 clkload23 (.A(clknet_leaf_51_clk));
 sg13g2_inv_1 clkload24 (.A(clknet_leaf_53_clk));
 sg13g2_buf_8 clkload25 (.A(clknet_leaf_47_clk));
 sg13g2_inv_1 clkload26 (.A(clknet_leaf_49_clk));
 sg13g2_inv_2 clkload27 (.A(clknet_leaf_50_clk));
 sg13g2_inv_2 clkload28 (.A(clknet_leaf_23_clk));
 sg13g2_inv_1 clkload29 (.A(clknet_leaf_57_clk));
 sg13g2_buf_1 clkload30 (.A(clknet_leaf_42_clk));
 sg13g2_inv_1 clkload31 (.A(clknet_leaf_45_clk));
 sg13g2_inv_2 clkload32 (.A(clknet_leaf_46_clk));
 sg13g2_inv_4 clkload33 (.A(clknet_leaf_7_clk));
 sg13g2_inv_2 clkload34 (.A(clknet_leaf_21_clk));
 sg13g2_inv_2 clkload35 (.A(clknet_leaf_15_clk));
 sg13g2_buf_8 clkload36 (.A(clknet_leaf_14_clk));
 sg13g2_inv_2 clkload37 (.A(clknet_leaf_13_clk));
 sg13g2_inv_4 clkload38 (.A(clknet_leaf_16_clk));
 sg13g2_inv_2 clkload39 (.A(clknet_leaf_17_clk));
 sg13g2_inv_1 clkload40 (.A(clknet_leaf_25_clk));
 sg13g2_inv_2 clkload41 (.A(clknet_leaf_36_clk));
 sg13g2_inv_2 clkload42 (.A(clknet_leaf_39_clk));
 sg13g2_inv_2 clkload43 (.A(clknet_leaf_29_clk));
 sg13g2_inv_2 clkload44 (.A(clknet_leaf_30_clk));
 sg13g2_buf_8 clkload45 (.A(clknet_leaf_31_clk));
 sg13g2_inv_1 clkload46 (.A(clknet_leaf_33_clk));
 sg13g2_inv_1 clkload47 (.A(clknet_leaf_35_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(mac_en_get_msu),
    .X(net274));
 sg13g2_dlygate4sd3_1 hold2 (.A(_00385_),
    .X(net275));
 sg13g2_dlygate4sd3_1 hold3 (.A(mac_en_get_mac),
    .X(net276));
 sg13g2_dlygate4sd3_1 hold4 (.A(_00386_),
    .X(net277));
 sg13g2_dlygate4sd3_1 hold5 (.A(mac_en_get_multiply),
    .X(net278));
 sg13g2_dlygate4sd3_1 hold6 (.A(_00384_),
    .X(net279));
 sg13g2_dlygate4sd3_1 hold7 (.A(\result_reg[6] ),
    .X(net280));
 sg13g2_dlygate4sd3_1 hold8 (.A(_00159_),
    .X(net281));
 sg13g2_dlygate4sd3_1 hold9 (.A(\result_reg[29] ),
    .X(net282));
 sg13g2_dlygate4sd3_1 hold10 (.A(_00068_),
    .X(net283));
 sg13g2_dlygate4sd3_1 hold11 (.A(\result_reg[67] ),
    .X(net284));
 sg13g2_dlygate4sd3_1 hold12 (.A(_00106_),
    .X(net285));
 sg13g2_dlygate4sd3_1 hold13 (.A(\result_reg[13] ),
    .X(net286));
 sg13g2_dlygate4sd3_1 hold14 (.A(_00166_),
    .X(net287));
 sg13g2_dlygate4sd3_1 hold15 (.A(\result_reg[53] ),
    .X(net288));
 sg13g2_dlygate4sd3_1 hold16 (.A(_00092_),
    .X(net289));
 sg13g2_dlygate4sd3_1 hold17 (.A(\result_reg[50] ),
    .X(net290));
 sg13g2_dlygate4sd3_1 hold18 (.A(_00089_),
    .X(net291));
 sg13g2_dlygate4sd3_1 hold19 (.A(\result_reg[26] ),
    .X(net292));
 sg13g2_dlygate4sd3_1 hold20 (.A(_00065_),
    .X(net293));
 sg13g2_dlygate4sd3_1 hold21 (.A(\result_reg[10] ),
    .X(net294));
 sg13g2_dlygate4sd3_1 hold22 (.A(_00163_),
    .X(net295));
 sg13g2_dlygate4sd3_1 hold23 (.A(\result_reg[11] ),
    .X(net296));
 sg13g2_dlygate4sd3_1 hold24 (.A(_00164_),
    .X(net297));
 sg13g2_dlygate4sd3_1 hold25 (.A(\result_reg[18] ),
    .X(net298));
 sg13g2_dlygate4sd3_1 hold26 (.A(_00171_),
    .X(net299));
 sg13g2_dlygate4sd3_1 hold27 (.A(\result_reg[27] ),
    .X(net300));
 sg13g2_dlygate4sd3_1 hold28 (.A(_00066_),
    .X(net301));
 sg13g2_dlygate4sd3_1 hold29 (.A(\result_reg[28] ),
    .X(net302));
 sg13g2_dlygate4sd3_1 hold30 (.A(_00067_),
    .X(net303));
 sg13g2_dlygate4sd3_1 hold31 (.A(\result_reg[4] ),
    .X(net304));
 sg13g2_dlygate4sd3_1 hold32 (.A(_00157_),
    .X(net305));
 sg13g2_dlygate4sd3_1 hold33 (.A(\result_reg[7] ),
    .X(net306));
 sg13g2_dlygate4sd3_1 hold34 (.A(_00160_),
    .X(net307));
 sg13g2_dlygate4sd3_1 hold35 (.A(\result_reg[60] ),
    .X(net308));
 sg13g2_dlygate4sd3_1 hold36 (.A(_00099_),
    .X(net309));
 sg13g2_dlygate4sd3_1 hold37 (.A(\result_reg[21] ),
    .X(net310));
 sg13g2_dlygate4sd3_1 hold38 (.A(_00174_),
    .X(net311));
 sg13g2_dlygate4sd3_1 hold39 (.A(\result_reg[3] ),
    .X(net312));
 sg13g2_dlygate4sd3_1 hold40 (.A(_00156_),
    .X(net313));
 sg13g2_dlygate4sd3_1 hold41 (.A(\result_reg[20] ),
    .X(net314));
 sg13g2_dlygate4sd3_1 hold42 (.A(_00173_),
    .X(net315));
 sg13g2_dlygate4sd3_1 hold43 (.A(\result_reg[41] ),
    .X(net316));
 sg13g2_dlygate4sd3_1 hold44 (.A(_00080_),
    .X(net317));
 sg13g2_dlygate4sd3_1 hold45 (.A(\result_reg[5] ),
    .X(net318));
 sg13g2_dlygate4sd3_1 hold46 (.A(_00158_),
    .X(net319));
 sg13g2_dlygate4sd3_1 hold47 (.A(\result_reg[42] ),
    .X(net320));
 sg13g2_dlygate4sd3_1 hold48 (.A(_00081_),
    .X(net321));
 sg13g2_dlygate4sd3_1 hold49 (.A(\result_reg[55] ),
    .X(net322));
 sg13g2_dlygate4sd3_1 hold50 (.A(_00094_),
    .X(net323));
 sg13g2_dlygate4sd3_1 hold51 (.A(\result_reg[30] ),
    .X(net324));
 sg13g2_dlygate4sd3_1 hold52 (.A(_00069_),
    .X(net325));
 sg13g2_dlygate4sd3_1 hold53 (.A(\result_reg[68] ),
    .X(net326));
 sg13g2_dlygate4sd3_1 hold54 (.A(_00107_),
    .X(net327));
 sg13g2_dlygate4sd3_1 hold55 (.A(\result_reg[0] ),
    .X(net328));
 sg13g2_dlygate4sd3_1 hold56 (.A(_00153_),
    .X(net329));
 sg13g2_dlygate4sd3_1 hold57 (.A(\result_reg[54] ),
    .X(net330));
 sg13g2_dlygate4sd3_1 hold58 (.A(_00093_),
    .X(net331));
 sg13g2_dlygate4sd3_1 hold59 (.A(\result_reg[46] ),
    .X(net332));
 sg13g2_dlygate4sd3_1 hold60 (.A(_00085_),
    .X(net333));
 sg13g2_dlygate4sd3_1 hold61 (.A(\result_reg[1] ),
    .X(net334));
 sg13g2_dlygate4sd3_1 hold62 (.A(_00154_),
    .X(net335));
 sg13g2_dlygate4sd3_1 hold63 (.A(\result_reg[22] ),
    .X(net336));
 sg13g2_dlygate4sd3_1 hold64 (.A(_00175_),
    .X(net337));
 sg13g2_dlygate4sd3_1 hold65 (.A(\result_reg[19] ),
    .X(net338));
 sg13g2_dlygate4sd3_1 hold66 (.A(_00172_),
    .X(net339));
 sg13g2_dlygate4sd3_1 hold67 (.A(\result_reg[25] ),
    .X(net340));
 sg13g2_dlygate4sd3_1 hold68 (.A(_00064_),
    .X(net341));
 sg13g2_dlygate4sd3_1 hold69 (.A(\result_reg[8] ),
    .X(net342));
 sg13g2_dlygate4sd3_1 hold70 (.A(_00161_),
    .X(net343));
 sg13g2_dlygate4sd3_1 hold71 (.A(\result_reg[43] ),
    .X(net344));
 sg13g2_dlygate4sd3_1 hold72 (.A(_00082_),
    .X(net345));
 sg13g2_dlygate4sd3_1 hold73 (.A(\result_reg[61] ),
    .X(net346));
 sg13g2_dlygate4sd3_1 hold74 (.A(_00100_),
    .X(net347));
 sg13g2_dlygate4sd3_1 hold75 (.A(\result_reg[59] ),
    .X(net348));
 sg13g2_dlygate4sd3_1 hold76 (.A(_00098_),
    .X(net349));
 sg13g2_dlygate4sd3_1 hold77 (.A(\result_reg[24] ),
    .X(net350));
 sg13g2_dlygate4sd3_1 hold78 (.A(_00063_),
    .X(net351));
 sg13g2_dlygate4sd3_1 hold79 (.A(\result_reg[23] ),
    .X(net352));
 sg13g2_dlygate4sd3_1 hold80 (.A(_00176_),
    .X(net353));
 sg13g2_dlygate4sd3_1 hold81 (.A(\mac_inst.get_multiply[6] ),
    .X(net354));
 sg13g2_dlygate4sd3_1 hold82 (.A(\mac_inst.get_multiply[0] ),
    .X(net355));
 sg13g2_dlygate4sd3_1 hold83 (.A(\result_reg[9] ),
    .X(net356));
 sg13g2_dlygate4sd3_1 hold84 (.A(_00162_),
    .X(net357));
 sg13g2_dlygate4sd3_1 hold85 (.A(\cordic_inst.get_normalize[62] ),
    .X(net358));
 sg13g2_dlygate4sd3_1 hold86 (.A(_02008_),
    .X(net359));
 sg13g2_dlygate4sd3_1 hold87 (.A(\result_reg[47] ),
    .X(net360));
 sg13g2_dlygate4sd3_1 hold88 (.A(_00086_),
    .X(net361));
 sg13g2_dlygate4sd3_1 hold89 (.A(\mac_inst.get_multiply[17] ),
    .X(net362));
 sg13g2_dlygate4sd3_1 hold90 (.A(\cordic_inst.get_normalize[63] ),
    .X(net363));
 sg13g2_dlygate4sd3_1 hold91 (.A(_00102_),
    .X(net364));
 sg13g2_dlygate4sd3_1 hold92 (.A(\mac_inst.get_msu[1] ),
    .X(net365));
 sg13g2_dlygate4sd3_1 hold93 (.A(_05168_),
    .X(net366));
 sg13g2_dlygate4sd3_1 hold94 (.A(_00337_),
    .X(net367));
 sg13g2_dlygate4sd3_1 hold95 (.A(\mac_inst.get_multiply[10] ),
    .X(net368));
 sg13g2_dlygate4sd3_1 hold96 (.A(\mac_inst.get_mac[3] ),
    .X(net369));
 sg13g2_dlygate4sd3_1 hold97 (.A(\mac_inst.get_multiply[2] ),
    .X(net370));
 sg13g2_dlygate4sd3_1 hold98 (.A(\mac_inst.get_msu[6] ),
    .X(net371));
 sg13g2_dlygate4sd3_1 hold99 (.A(_05207_),
    .X(net372));
 sg13g2_dlygate4sd3_1 hold100 (.A(_00342_),
    .X(net373));
 sg13g2_dlygate4sd3_1 hold101 (.A(\mac_inst.get_multiply[13] ),
    .X(net374));
 sg13g2_dlygate4sd3_1 hold102 (.A(\cordic_inst.get_normalize[27] ),
    .X(net375));
 sg13g2_dlygate4sd3_1 hold103 (.A(_02021_),
    .X(net376));
 sg13g2_dlygate4sd3_1 hold104 (.A(\mac_inst.get_msu[7] ),
    .X(net377));
 sg13g2_dlygate4sd3_1 hold105 (.A(\mac_inst.get_mac[5] ),
    .X(net378));
 sg13g2_dlygate4sd3_1 hold106 (.A(\cordic_inst.get_normalize[71] ),
    .X(net379));
 sg13g2_dlygate4sd3_1 hold107 (.A(_00110_),
    .X(net380));
 sg13g2_dlygate4sd3_1 hold108 (.A(\result_reg[44] ),
    .X(net381));
 sg13g2_dlygate4sd3_1 hold109 (.A(_00083_),
    .X(net382));
 sg13g2_dlygate4sd3_1 hold110 (.A(\cordic_inst.get_normalize[57] ),
    .X(net383));
 sg13g2_dlygate4sd3_1 hold111 (.A(_00096_),
    .X(net384));
 sg13g2_dlygate4sd3_1 hold112 (.A(\result_reg[2] ),
    .X(net385));
 sg13g2_dlygate4sd3_1 hold113 (.A(_00155_),
    .X(net386));
 sg13g2_dlygate4sd3_1 hold114 (.A(\result_reg[17] ),
    .X(net387));
 sg13g2_dlygate4sd3_1 hold115 (.A(_00170_),
    .X(net388));
 sg13g2_dlygate4sd3_1 hold116 (.A(\result_reg[39] ),
    .X(net389));
 sg13g2_dlygate4sd3_1 hold117 (.A(_00078_),
    .X(net390));
 sg13g2_dlygate4sd3_1 hold118 (.A(\cordic_inst.get_normalize[38] ),
    .X(net391));
 sg13g2_dlygate4sd3_1 hold119 (.A(_02032_),
    .X(net392));
 sg13g2_dlygate4sd3_1 hold120 (.A(\result_reg[64] ),
    .X(net393));
 sg13g2_dlygate4sd3_1 hold121 (.A(_00103_),
    .X(net394));
 sg13g2_dlygate4sd3_1 hold122 (.A(\result_reg[49] ),
    .X(net395));
 sg13g2_dlygate4sd3_1 hold123 (.A(_00088_),
    .X(net396));
 sg13g2_dlygate4sd3_1 hold124 (.A(\cordic_inst.get_normalize[50] ),
    .X(net397));
 sg13g2_dlygate4sd3_1 hold125 (.A(_01996_),
    .X(net398));
 sg13g2_dlygate4sd3_1 hold126 (.A(\cordic_inst.get_normalize[66] ),
    .X(net399));
 sg13g2_dlygate4sd3_1 hold127 (.A(_02012_),
    .X(net400));
 sg13g2_dlygate4sd3_1 hold128 (.A(\cordic_inst.MUX_cordic_state$write_1__VAL_1[71] ),
    .X(net401));
 sg13g2_dlygate4sd3_1 hold129 (.A(\result_reg[35] ),
    .X(net402));
 sg13g2_dlygate4sd3_1 hold130 (.A(_00074_),
    .X(net403));
 sg13g2_dlygate4sd3_1 hold131 (.A(\mac_inst.get_multiply[14] ),
    .X(net404));
 sg13g2_dlygate4sd3_1 hold132 (.A(\mac_inst.get_msu[11] ),
    .X(net405));
 sg13g2_dlygate4sd3_1 hold133 (.A(\mac_inst.get_msu[23] ),
    .X(net406));
 sg13g2_dlygate4sd3_1 hold134 (.A(_05362_),
    .X(net407));
 sg13g2_dlygate4sd3_1 hold135 (.A(\mac_inst.get_msu[2] ),
    .X(net408));
 sg13g2_dlygate4sd3_1 hold136 (.A(_05176_),
    .X(net409));
 sg13g2_dlygate4sd3_1 hold137 (.A(\result_reg[31] ),
    .X(net410));
 sg13g2_dlygate4sd3_1 hold138 (.A(_00070_),
    .X(net411));
 sg13g2_dlygate4sd3_1 hold139 (.A(\cordic_inst.get_normalize[29] ),
    .X(net412));
 sg13g2_dlygate4sd3_1 hold140 (.A(_02023_),
    .X(net413));
 sg13g2_dlygate4sd3_1 hold141 (.A(\cordic_inst.get_normalize[32] ),
    .X(net414));
 sg13g2_dlygate4sd3_1 hold142 (.A(_02026_),
    .X(net415));
 sg13g2_dlygate4sd3_1 hold143 (.A(\cordic_inst.get_normalize[60] ),
    .X(net416));
 sg13g2_dlygate4sd3_1 hold144 (.A(_02006_),
    .X(net417));
 sg13g2_dlygate4sd3_1 hold145 (.A(\cordic_inst.get_normalize[48] ),
    .X(net418));
 sg13g2_dlygate4sd3_1 hold146 (.A(_00087_),
    .X(net419));
 sg13g2_dlygate4sd3_1 hold147 (.A(\mac_inst.get_msu[4] ),
    .X(net420));
 sg13g2_dlygate4sd3_1 hold148 (.A(_05191_),
    .X(net421));
 sg13g2_dlygate4sd3_1 hold149 (.A(\cordic_inst.get_normalize[46] ),
    .X(net422));
 sg13g2_dlygate4sd3_1 hold150 (.A(_02040_),
    .X(net423));
 sg13g2_dlygate4sd3_1 hold151 (.A(\mac_inst.get_multiply[15] ),
    .X(net424));
 sg13g2_dlygate4sd3_1 hold152 (.A(\cordic_inst.get_normalize[61] ),
    .X(net425));
 sg13g2_dlygate4sd3_1 hold153 (.A(_02007_),
    .X(net426));
 sg13g2_dlygate4sd3_1 hold154 (.A(\mac_inst.get_multiply[21] ),
    .X(net427));
 sg13g2_dlygate4sd3_1 hold155 (.A(\cordic_inst.MUX_cordic_state$write_1__VAL_1[65] ),
    .X(net428));
 sg13g2_dlygate4sd3_1 hold156 (.A(\cordic_inst.get_normalize[64] ),
    .X(net429));
 sg13g2_dlygate4sd3_1 hold157 (.A(_02010_),
    .X(net430));
 sg13g2_dlygate4sd3_1 hold158 (.A(\result_reg[37] ),
    .X(net431));
 sg13g2_dlygate4sd3_1 hold159 (.A(_00076_),
    .X(net432));
 sg13g2_dlygate4sd3_1 hold160 (.A(\mac_inst.get_msu[12] ),
    .X(net433));
 sg13g2_dlygate4sd3_1 hold161 (.A(\cordic_inst.get_normalize[52] ),
    .X(net434));
 sg13g2_dlygate4sd3_1 hold162 (.A(_01998_),
    .X(net435));
 sg13g2_dlygate4sd3_1 hold163 (.A(\cordic_inst.get_normalize[25] ),
    .X(net436));
 sg13g2_dlygate4sd3_1 hold164 (.A(_02019_),
    .X(net437));
 sg13g2_dlygate4sd3_1 hold165 (.A(\cordic_inst.get_normalize[53] ),
    .X(net438));
 sg13g2_dlygate4sd3_1 hold166 (.A(_01999_),
    .X(net439));
 sg13g2_dlygate4sd3_1 hold167 (.A(\result_reg[65] ),
    .X(net440));
 sg13g2_dlygate4sd3_1 hold168 (.A(_00104_),
    .X(net441));
 sg13g2_dlygate4sd3_1 hold169 (.A(\cordic_inst.get_normalize[68] ),
    .X(net442));
 sg13g2_dlygate4sd3_1 hold170 (.A(_02014_),
    .X(net443));
 sg13g2_dlygate4sd3_1 hold171 (.A(\cordic_inst.get_normalize[24] ),
    .X(net444));
 sg13g2_dlygate4sd3_1 hold172 (.A(_02018_),
    .X(net445));
 sg13g2_dlygate4sd3_1 hold173 (.A(\cordic_inst.get_normalize[59] ),
    .X(net446));
 sg13g2_dlygate4sd3_1 hold174 (.A(_02005_),
    .X(net447));
 sg13g2_dlygate4sd3_1 hold175 (.A(\mac_inst.get_msu[22] ),
    .X(net448));
 sg13g2_dlygate4sd3_1 hold176 (.A(\cordic_inst.get_normalize[34] ),
    .X(net449));
 sg13g2_dlygate4sd3_1 hold177 (.A(_02028_),
    .X(net450));
 sg13g2_dlygate4sd3_1 hold178 (.A(\result_reg[38] ),
    .X(net451));
 sg13g2_dlygate4sd3_1 hold179 (.A(_00077_),
    .X(net452));
 sg13g2_dlygate4sd3_1 hold180 (.A(\cordic_inst.get_normalize[56] ),
    .X(net453));
 sg13g2_dlygate4sd3_1 hold181 (.A(_02002_),
    .X(net454));
 sg13g2_dlygate4sd3_1 hold182 (.A(\cordic_inst.get_normalize[37] ),
    .X(net455));
 sg13g2_dlygate4sd3_1 hold183 (.A(_02031_),
    .X(net456));
 sg13g2_dlygate4sd3_1 hold184 (.A(\cordic_inst.get_normalize[42] ),
    .X(net457));
 sg13g2_dlygate4sd3_1 hold185 (.A(_02036_),
    .X(net458));
 sg13g2_dlygate4sd3_1 hold186 (.A(\cordic_inst.get_normalize[58] ),
    .X(net459));
 sg13g2_dlygate4sd3_1 hold187 (.A(_02004_),
    .X(net460));
 sg13g2_dlygate4sd3_1 hold188 (.A(\mac_inst.get_msu[13] ),
    .X(net461));
 sg13g2_dlygate4sd3_1 hold189 (.A(_00349_),
    .X(net462));
 sg13g2_dlygate4sd3_1 hold190 (.A(\cordic_inst.MUX_cordic_state$write_1__VAL_1[56] ),
    .X(net463));
 sg13g2_dlygate4sd3_1 hold191 (.A(\cordic_inst.get_normalize[36] ),
    .X(net464));
 sg13g2_dlygate4sd3_1 hold192 (.A(_02030_),
    .X(net465));
 sg13g2_dlygate4sd3_1 hold193 (.A(\cordic_inst.get_normalize[51] ),
    .X(net466));
 sg13g2_dlygate4sd3_1 hold194 (.A(_00090_),
    .X(net467));
 sg13g2_dlygate4sd3_1 hold195 (.A(\mac_inst.get_multiply[19] ),
    .X(net468));
 sg13g2_dlygate4sd3_1 hold196 (.A(\cordic_inst.MUX_cordic_state$write_1__VAL_1[79] ),
    .X(net469));
 sg13g2_dlygate4sd3_1 hold197 (.A(\cordic_inst.get_normalize[45] ),
    .X(net470));
 sg13g2_dlygate4sd3_1 hold198 (.A(_02039_),
    .X(net471));
 sg13g2_dlygate4sd3_1 hold199 (.A(\cordic_inst.get_normalize[49] ),
    .X(net472));
 sg13g2_dlygate4sd3_1 hold200 (.A(_01995_),
    .X(net473));
 sg13g2_dlygate4sd3_1 hold201 (.A(\cordic_inst.get_normalize[69] ),
    .X(net474));
 sg13g2_dlygate4sd3_1 hold202 (.A(_00108_),
    .X(net475));
 sg13g2_dlygate4sd3_1 hold203 (.A(\mac_inst.get_msu[0] ),
    .X(net476));
 sg13g2_dlygate4sd3_1 hold204 (.A(_05160_),
    .X(net477));
 sg13g2_dlygate4sd3_1 hold205 (.A(\result_reg[33] ),
    .X(net478));
 sg13g2_dlygate4sd3_1 hold206 (.A(_00072_),
    .X(net479));
 sg13g2_dlygate4sd3_1 hold207 (.A(\result_reg[45] ),
    .X(net480));
 sg13g2_dlygate4sd3_1 hold208 (.A(_00084_),
    .X(net481));
 sg13g2_dlygate4sd3_1 hold209 (.A(\cordic_inst.MUX_cordic_state$write_1__VAL_1[77] ),
    .X(net482));
 sg13g2_dlygate4sd3_1 hold210 (.A(\cordic_inst.operation_pending ),
    .X(net483));
 sg13g2_dlygate4sd3_1 hold211 (.A(_01990_),
    .X(net484));
 sg13g2_dlygate4sd3_1 hold212 (.A(_00262_),
    .X(net485));
 sg13g2_dlygate4sd3_1 hold213 (.A(\result_reg[66] ),
    .X(net486));
 sg13g2_dlygate4sd3_1 hold214 (.A(\mac_inst.get_msu[5] ),
    .X(net487));
 sg13g2_dlygate4sd3_1 hold215 (.A(_05199_),
    .X(net488));
 sg13g2_dlygate4sd3_1 hold216 (.A(\cordic_inst.get_normalize[39] ),
    .X(net489));
 sg13g2_dlygate4sd3_1 hold217 (.A(_02033_),
    .X(net490));
 sg13g2_dlygate4sd3_1 hold218 (.A(\result_reg[56] ),
    .X(net491));
 sg13g2_dlygate4sd3_1 hold219 (.A(\cordic_inst.get_normalize[54] ),
    .X(net492));
 sg13g2_dlygate4sd3_1 hold220 (.A(_02000_),
    .X(net493));
 sg13g2_dlygate4sd3_1 hold221 (.A(\cordic_inst.get_normalize[30] ),
    .X(net494));
 sg13g2_dlygate4sd3_1 hold222 (.A(_02024_),
    .X(net495));
 sg13g2_dlygate4sd3_1 hold223 (.A(\mac_inst.get_msu[17] ),
    .X(net496));
 sg13g2_dlygate4sd3_1 hold224 (.A(_00353_),
    .X(net497));
 sg13g2_dlygate4sd3_1 hold225 (.A(\result_reg[52] ),
    .X(net498));
 sg13g2_dlygate4sd3_1 hold226 (.A(\cordic_inst.operation_started ),
    .X(net499));
 sg13g2_dlygate4sd3_1 hold227 (.A(_01987_),
    .X(net500));
 sg13g2_dlygate4sd3_1 hold228 (.A(\mac_inst.get_multiply[20] ),
    .X(net501));
 sg13g2_dlygate4sd3_1 hold229 (.A(\cordic_inst.get_normalize[35] ),
    .X(net502));
 sg13g2_dlygate4sd3_1 hold230 (.A(_02029_),
    .X(net503));
 sg13g2_dlygate4sd3_1 hold231 (.A(\result_reg[36] ),
    .X(net504));
 sg13g2_dlygate4sd3_1 hold232 (.A(_00075_),
    .X(net505));
 sg13g2_dlygate4sd3_1 hold233 (.A(\mac_inst.get_msu[18] ),
    .X(net506));
 sg13g2_dlygate4sd3_1 hold234 (.A(\cordic_inst.get_normalize[70] ),
    .X(net507));
 sg13g2_dlygate4sd3_1 hold235 (.A(_02016_),
    .X(net508));
 sg13g2_dlygate4sd3_1 hold236 (.A(\result_reg[58] ),
    .X(net509));
 sg13g2_dlygate4sd3_1 hold237 (.A(\mac_inst.get_msu[21] ),
    .X(net510));
 sg13g2_dlygate4sd3_1 hold238 (.A(\cordic_inst.get_normalize[33] ),
    .X(net511));
 sg13g2_dlygate4sd3_1 hold239 (.A(_02027_),
    .X(net512));
 sg13g2_dlygate4sd3_1 hold240 (.A(\cordic_inst.get_normalize[40] ),
    .X(net513));
 sg13g2_dlygate4sd3_1 hold241 (.A(_02034_),
    .X(net514));
 sg13g2_dlygate4sd3_1 hold242 (.A(\mac_inst.get_mac[4] ),
    .X(net515));
 sg13g2_dlygate4sd3_1 hold243 (.A(\cordic_inst.get_normalize[31] ),
    .X(net516));
 sg13g2_dlygate4sd3_1 hold244 (.A(_02025_),
    .X(net517));
 sg13g2_dlygate4sd3_1 hold245 (.A(\cordic_inst.get_normalize[43] ),
    .X(net518));
 sg13g2_dlygate4sd3_1 hold246 (.A(_02037_),
    .X(net519));
 sg13g2_dlygate4sd3_1 hold247 (.A(\cordic_inst.get_normalize[65] ),
    .X(net520));
 sg13g2_dlygate4sd3_1 hold248 (.A(_02011_),
    .X(net521));
 sg13g2_dlygate4sd3_1 hold249 (.A(\mac_inst.get_msu[3] ),
    .X(net522));
 sg13g2_dlygate4sd3_1 hold250 (.A(\cordic_inst.current_op[3] ),
    .X(net523));
 sg13g2_dlygate4sd3_1 hold251 (.A(\result_reg[32] ),
    .X(net524));
 sg13g2_dlygate4sd3_1 hold252 (.A(_00071_),
    .X(net525));
 sg13g2_dlygate4sd3_1 hold253 (.A(\result_reg[70] ),
    .X(net526));
 sg13g2_dlygate4sd3_1 hold254 (.A(\mac_inst.get_multiply[22] ),
    .X(net527));
 sg13g2_dlygate4sd3_1 hold255 (.A(\cordic_inst.get_normalize[47] ),
    .X(net528));
 sg13g2_dlygate4sd3_1 hold256 (.A(_02041_),
    .X(net529));
 sg13g2_dlygate4sd3_1 hold257 (.A(\result_reg[40] ),
    .X(net530));
 sg13g2_dlygate4sd3_1 hold258 (.A(_00079_),
    .X(net531));
 sg13g2_dlygate4sd3_1 hold259 (.A(\result_reg[34] ),
    .X(net532));
 sg13g2_dlygate4sd3_1 hold260 (.A(_00073_),
    .X(net533));
 sg13g2_dlygate4sd3_1 hold261 (.A(\mac_inst.get_msu[14] ),
    .X(net534));
 sg13g2_dlygate4sd3_1 hold262 (.A(_00350_),
    .X(net535));
 sg13g2_dlygate4sd3_1 hold263 (.A(\cordic_inst.MUX_cordic_state$write_1__VAL_1[59] ),
    .X(net536));
 sg13g2_dlygate4sd3_1 hold264 (.A(\mac_inst.get_mac[6] ),
    .X(net537));
 sg13g2_dlygate4sd3_1 hold265 (.A(\mac_inst.get_mac[1] ),
    .X(net538));
 sg13g2_dlygate4sd3_1 hold266 (.A(_05368_),
    .X(net539));
 sg13g2_dlygate4sd3_1 hold267 (.A(\result_reg[62] ),
    .X(net540));
 sg13g2_dlygate4sd3_1 hold268 (.A(\cordic_inst.get_normalize[67] ),
    .X(net541));
 sg13g2_dlygate4sd3_1 hold269 (.A(_02013_),
    .X(net542));
 sg13g2_dlygate4sd3_1 hold270 (.A(\mac_inst.get_mac[2] ),
    .X(net543));
 sg13g2_dlygate4sd3_1 hold271 (.A(_05372_),
    .X(net544));
 sg13g2_dlygate4sd3_1 hold272 (.A(\cordic_inst.current_op[2] ),
    .X(net545));
 sg13g2_dlygate4sd3_1 hold273 (.A(\cordic_inst.get_normalize[41] ),
    .X(net546));
 sg13g2_dlygate4sd3_1 hold274 (.A(_02035_),
    .X(net547));
 sg13g2_dlygate4sd3_1 hold275 (.A(\mac_inst.get_msu[19] ),
    .X(net548));
 sg13g2_dlygate4sd3_1 hold276 (.A(_00355_),
    .X(net549));
 sg13g2_dlygate4sd3_1 hold277 (.A(\mac_inst.get_mac[7] ),
    .X(net550));
 sg13g2_dlygate4sd3_1 hold278 (.A(\mac_inst.get_mac[22] ),
    .X(net551));
 sg13g2_dlygate4sd3_1 hold279 (.A(\mac_inst.accumulator[12] ),
    .X(net552));
 sg13g2_dlygate4sd3_1 hold280 (.A(\mac_inst.get_msu[20] ),
    .X(net553));
 sg13g2_dlygate4sd3_1 hold281 (.A(\mac_inst.accumulator[9] ),
    .X(net554));
 sg13g2_dlygate4sd3_1 hold282 (.A(\cordic_inst.get_normalize[44] ),
    .X(net555));
 sg13g2_dlygate4sd3_1 hold283 (.A(_02038_),
    .X(net556));
 sg13g2_dlygate4sd3_1 hold284 (.A(\mac_inst.get_msu[10] ),
    .X(net557));
 sg13g2_dlygate4sd3_1 hold285 (.A(\mac_inst.get_mac[18] ),
    .X(net558));
 sg13g2_dlygate4sd3_1 hold286 (.A(_05460_),
    .X(net559));
 sg13g2_dlygate4sd3_1 hold287 (.A(\mac_inst.get_mac[8] ),
    .X(net560));
 sg13g2_dlygate4sd3_1 hold288 (.A(\mac_inst.get_mac[9] ),
    .X(net561));
 sg13g2_dlygate4sd3_1 hold289 (.A(_00369_),
    .X(net562));
 sg13g2_dlygate4sd3_1 hold290 (.A(\mac_inst.get_mac[12] ),
    .X(net563));
 sg13g2_dlygate4sd3_1 hold291 (.A(\cordic_inst.current_op[1] ),
    .X(net564));
 sg13g2_dlygate4sd3_1 hold292 (.A(_00475_),
    .X(net565));
 sg13g2_dlygate4sd3_1 hold293 (.A(\result_reg[14] ),
    .X(net566));
 sg13g2_dlygate4sd3_1 hold294 (.A(_00167_),
    .X(net567));
 sg13g2_dlygate4sd3_1 hold295 (.A(\cmd_reg[7] ),
    .X(net568));
 sg13g2_dlygate4sd3_1 hold296 (.A(_00136_),
    .X(net569));
 sg13g2_dlygate4sd3_1 hold297 (.A(\mac_inst.get_mac[14] ),
    .X(net570));
 sg13g2_dlygate4sd3_1 hold298 (.A(\result_reg[15] ),
    .X(net571));
 sg13g2_dlygate4sd3_1 hold299 (.A(_00168_),
    .X(net572));
 sg13g2_dlygate4sd3_1 hold300 (.A(\mac_inst.get_msu[15] ),
    .X(net573));
 sg13g2_dlygate4sd3_1 hold301 (.A(_00028_),
    .X(net574));
 sg13g2_dlygate4sd3_1 hold302 (.A(_00027_),
    .X(net575));
 sg13g2_dlygate4sd3_1 hold303 (.A(\result_reg[12] ),
    .X(net576));
 sg13g2_dlygate4sd3_1 hold304 (.A(_00165_),
    .X(net577));
 sg13g2_dlygate4sd3_1 hold305 (.A(\cordic_inst.get_normalize[55] ),
    .X(net578));
 sg13g2_dlygate4sd3_1 hold306 (.A(_02001_),
    .X(net579));
 sg13g2_dlygate4sd3_1 hold307 (.A(\mac_inst.get_multiply[7] ),
    .X(net580));
 sg13g2_dlygate4sd3_1 hold308 (.A(\mac_inst.get_mac[16] ),
    .X(net581));
 sg13g2_dlygate4sd3_1 hold309 (.A(\cmd_reg[6] ),
    .X(net582));
 sg13g2_dlygate4sd3_1 hold310 (.A(_00135_),
    .X(net583));
 sg13g2_dlygate4sd3_1 hold311 (.A(\cordic_atan2_result[10] ),
    .X(net584));
 sg13g2_dlygate4sd3_1 hold312 (.A(_00199_),
    .X(net585));
 sg13g2_dlygate4sd3_1 hold313 (.A(\mac_inst.get_msu[9] ),
    .X(net586));
 sg13g2_dlygate4sd3_1 hold314 (.A(_00345_),
    .X(net587));
 sg13g2_dlygate4sd3_1 hold315 (.A(\mac_inst.get_mac[10] ),
    .X(net588));
 sg13g2_dlygate4sd3_1 hold316 (.A(\mac_inst.get_mac[15] ),
    .X(net589));
 sg13g2_dlygate4sd3_1 hold317 (.A(_05440_),
    .X(net590));
 sg13g2_dlygate4sd3_1 hold318 (.A(_00375_),
    .X(net591));
 sg13g2_dlygate4sd3_1 hold319 (.A(\mac_inst.get_msu[16] ),
    .X(net592));
 sg13g2_dlygate4sd3_1 hold320 (.A(\mac_inst.get_mac[20] ),
    .X(net593));
 sg13g2_dlygate4sd3_1 hold321 (.A(\mac_inst.get_multiply[3] ),
    .X(net594));
 sg13g2_dlygate4sd3_1 hold322 (.A(\mac_inst.get_msu[8] ),
    .X(net595));
 sg13g2_dlygate4sd3_1 hold323 (.A(_00344_),
    .X(net596));
 sg13g2_dlygate4sd3_1 hold324 (.A(\mac_inst.get_multiply[5] ),
    .X(net597));
 sg13g2_dlygate4sd3_1 hold325 (.A(\mac_inst.get_mac[0] ),
    .X(net598));
 sg13g2_dlygate4sd3_1 hold326 (.A(_05365_),
    .X(net599));
 sg13g2_dlygate4sd3_1 hold327 (.A(\mac_inst.get_mac[17] ),
    .X(net600));
 sg13g2_dlygate4sd3_1 hold328 (.A(_00377_),
    .X(net601));
 sg13g2_dlygate4sd3_1 hold329 (.A(\mac_inst.get_mac[13] ),
    .X(net602));
 sg13g2_dlygate4sd3_1 hold330 (.A(\mac_inst.get_multiply[4] ),
    .X(net603));
 sg13g2_dlygate4sd3_1 hold331 (.A(_00316_),
    .X(net604));
 sg13g2_dlygate4sd3_1 hold332 (.A(\result_reg[16] ),
    .X(net605));
 sg13g2_dlygate4sd3_1 hold333 (.A(_00169_),
    .X(net606));
 sg13g2_dlygate4sd3_1 hold334 (.A(\mac_inst.get_mac[11] ),
    .X(net607));
 sg13g2_dlygate4sd3_1 hold335 (.A(_00371_),
    .X(net608));
 sg13g2_dlygate4sd3_1 hold336 (.A(\cordic_inst.get_normalize[26] ),
    .X(net609));
 sg13g2_dlygate4sd3_1 hold337 (.A(\mac_inst.accumulator[17] ),
    .X(net610));
 sg13g2_dlygate4sd3_1 hold338 (.A(_05523_),
    .X(net611));
 sg13g2_dlygate4sd3_1 hold339 (.A(\cordic_inst.get_normalize[28] ),
    .X(net612));
 sg13g2_dlygate4sd3_1 hold340 (.A(_02022_),
    .X(net613));
 sg13g2_dlygate4sd3_1 hold341 (.A(\mac_inst.get_multiply[9] ),
    .X(net614));
 sg13g2_dlygate4sd3_1 hold342 (.A(\mac_inst.get_multiply[1] ),
    .X(net615));
 sg13g2_dlygate4sd3_1 hold343 (.A(_02528_),
    .X(net616));
 sg13g2_dlygate4sd3_1 hold344 (.A(_00313_),
    .X(net617));
 sg13g2_dlygate4sd3_1 hold345 (.A(\mac_inst.get_multiply[11] ),
    .X(net618));
 sg13g2_dlygate4sd3_1 hold346 (.A(\cmd_reg[5] ),
    .X(net619));
 sg13g2_dlygate4sd3_1 hold347 (.A(_00134_),
    .X(net620));
 sg13g2_dlygate4sd3_1 hold348 (.A(\mac_inst.get_multiply[16] ),
    .X(net621));
 sg13g2_dlygate4sd3_1 hold349 (.A(_04332_),
    .X(net622));
 sg13g2_dlygate4sd3_1 hold350 (.A(_00328_),
    .X(net623));
 sg13g2_dlygate4sd3_1 hold351 (.A(\mac_inst.get_multiply[12] ),
    .X(net624));
 sg13g2_dlygate4sd3_1 hold352 (.A(\cmd_reg[4] ),
    .X(net625));
 sg13g2_dlygate4sd3_1 hold353 (.A(_00133_),
    .X(net626));
 sg13g2_dlygate4sd3_1 hold354 (.A(\cordic_inst.cordic_state[52] ),
    .X(net627));
 sg13g2_dlygate4sd3_1 hold355 (.A(\mac_inst.get_multiply[18] ),
    .X(net628));
 sg13g2_dlygate4sd3_1 hold356 (.A(_04582_),
    .X(net629));
 sg13g2_dlygate4sd3_1 hold357 (.A(_00330_),
    .X(net630));
 sg13g2_dlygate4sd3_1 hold358 (.A(uo_out[0]),
    .X(net631));
 sg13g2_dlygate4sd3_1 hold359 (.A(_00692_),
    .X(net632));
 sg13g2_dlygate4sd3_1 hold360 (.A(cordic_en_get_sqrt),
    .X(net633));
 sg13g2_dlygate4sd3_1 hold361 (.A(_01991_),
    .X(net634));
 sg13g2_dlygate4sd3_1 hold362 (.A(_01993_),
    .X(net635));
 sg13g2_dlygate4sd3_1 hold363 (.A(uo_out[5]),
    .X(net636));
 sg13g2_dlygate4sd3_1 hold364 (.A(_00732_),
    .X(net637));
 sg13g2_dlygate4sd3_1 hold365 (.A(\mac_inst.get_multiply[8] ),
    .X(net638));
 sg13g2_dlygate4sd3_1 hold366 (.A(\mac_inst.get_mac[21] ),
    .X(net639));
 sg13g2_dlygate4sd3_1 hold367 (.A(_00381_),
    .X(net640));
 sg13g2_dlygate4sd3_1 hold368 (.A(uo_out[6]),
    .X(net641));
 sg13g2_dlygate4sd3_1 hold369 (.A(_00740_),
    .X(net642));
 sg13g2_dlygate4sd3_1 hold370 (.A(\mac_inst.get_mac[19] ),
    .X(net643));
 sg13g2_dlygate4sd3_1 hold371 (.A(uo_out[1]),
    .X(net644));
 sg13g2_dlygate4sd3_1 hold372 (.A(_00700_),
    .X(net645));
 sg13g2_dlygate4sd3_1 hold373 (.A(\cordic_atan2_result[18] ),
    .X(net646));
 sg13g2_dlygate4sd3_1 hold374 (.A(uo_out[2]),
    .X(net647));
 sg13g2_dlygate4sd3_1 hold375 (.A(_00708_),
    .X(net648));
 sg13g2_dlygate4sd3_1 hold376 (.A(uo_out[3]),
    .X(net649));
 sg13g2_dlygate4sd3_1 hold377 (.A(_00716_),
    .X(net650));
 sg13g2_dlygate4sd3_1 hold378 (.A(\mac_inst.accumulator[23] ),
    .X(net651));
 sg13g2_dlygate4sd3_1 hold379 (.A(_00410_),
    .X(net652));
 sg13g2_dlygate4sd3_1 hold380 (.A(\cordic_atan2_result[14] ),
    .X(net653));
 sg13g2_dlygate4sd3_1 hold381 (.A(_01065_),
    .X(net654));
 sg13g2_dlygate4sd3_1 hold382 (.A(uo_out[4]),
    .X(net655));
 sg13g2_dlygate4sd3_1 hold383 (.A(_00724_),
    .X(net656));
 sg13g2_dlygate4sd3_1 hold384 (.A(\cordic_atan2_result[4] ),
    .X(net657));
 sg13g2_dlygate4sd3_1 hold385 (.A(\mac_inst.get_multiply[23] ),
    .X(net658));
 sg13g2_dlygate4sd3_1 hold386 (.A(_05155_),
    .X(net659));
 sg13g2_dlygate4sd3_1 hold387 (.A(_00335_),
    .X(net660));
 sg13g2_dlygate4sd3_1 hold388 (.A(\cordic_inst.current_op[0] ),
    .X(net661));
 sg13g2_dlygate4sd3_1 hold389 (.A(_00473_),
    .X(net662));
 sg13g2_dlygate4sd3_1 hold390 (.A(\exec_phase[1] ),
    .X(net663));
 sg13g2_dlygate4sd3_1 hold391 (.A(_00468_),
    .X(net664));
 sg13g2_dlygate4sd3_1 hold392 (.A(_00026_),
    .X(net665));
 sg13g2_dlygate4sd3_1 hold393 (.A(\mac_inst.get_mac[23] ),
    .X(net666));
 sg13g2_dlygate4sd3_1 hold394 (.A(_00383_),
    .X(net667));
 sg13g2_dlygate4sd3_1 hold395 (.A(\byte_counter[2] ),
    .X(net668));
 sg13g2_dlygate4sd3_1 hold396 (.A(_00179_),
    .X(net669));
 sg13g2_dlygate4sd3_1 hold397 (.A(\cordic_atan2_result[6] ),
    .X(net670));
 sg13g2_dlygate4sd3_1 hold398 (.A(_00983_),
    .X(net671));
 sg13g2_dlygate4sd3_1 hold399 (.A(\cordic_atan2_result[0] ),
    .X(net672));
 sg13g2_dlygate4sd3_1 hold400 (.A(_00189_),
    .X(net673));
 sg13g2_dlygate4sd3_1 hold401 (.A(\cordic_atan2_result[13] ),
    .X(net674));
 sg13g2_dlygate4sd3_1 hold402 (.A(_01056_),
    .X(net675));
 sg13g2_dlygate4sd3_1 hold403 (.A(\cordic_atan2_result[17] ),
    .X(net676));
 sg13g2_dlygate4sd3_1 hold404 (.A(\cordic_inst.cordic_state[48] ),
    .X(net677));
 sg13g2_dlygate4sd3_1 hold405 (.A(\cordic_inst.cordic_state[59] ),
    .X(net678));
 sg13g2_dlygate4sd3_1 hold406 (.A(\cordic_atan2_result[22] ),
    .X(net679));
 sg13g2_dlygate4sd3_1 hold407 (.A(\cordic_inst.cordic_state[62] ),
    .X(net680));
 sg13g2_dlygate4sd3_1 hold408 (.A(\cordic_atan2_result[16] ),
    .X(net681));
 sg13g2_dlygate4sd3_1 hold409 (.A(\cordic_atan2_result[5] ),
    .X(net682));
 sg13g2_dlygate4sd3_1 hold410 (.A(_00973_),
    .X(net683));
 sg13g2_dlygate4sd3_1 hold411 (.A(\mac_inst.accumulator[21] ),
    .X(net684));
 sg13g2_dlygate4sd3_1 hold412 (.A(\cordic_inst.IF_IF_cordic_state_BITS_2_TO_1_EQ_1_THEN_NOT_c_ETC___d36[1] ),
    .X(net685));
 sg13g2_dlygate4sd3_1 hold413 (.A(\cordic_atan2_result[11] ),
    .X(net686));
 sg13g2_dlygate4sd3_1 hold414 (.A(_01034_),
    .X(net687));
 sg13g2_dlygate4sd3_1 hold415 (.A(\cordic_inst.cordic_state[41] ),
    .X(net688));
 sg13g2_dlygate4sd3_1 hold416 (.A(\cordic_inst.cordic_state[35] ),
    .X(net689));
 sg13g2_dlygate4sd3_1 hold417 (.A(\cordic_atan2_result[7] ),
    .X(net690));
 sg13g2_dlygate4sd3_1 hold418 (.A(\cmd_reg[3] ),
    .X(net691));
 sg13g2_dlygate4sd3_1 hold419 (.A(_00132_),
    .X(net692));
 sg13g2_dlygate4sd3_1 hold420 (.A(\cmd_reg[1] ),
    .X(net693));
 sg13g2_dlygate4sd3_1 hold421 (.A(_00130_),
    .X(net694));
 sg13g2_dlygate4sd3_1 hold422 (.A(\cordic_atan2_result[2] ),
    .X(net695));
 sg13g2_dlygate4sd3_1 hold423 (.A(_00945_),
    .X(net696));
 sg13g2_dlygate4sd3_1 hold424 (.A(\cordic_atan2_result[12] ),
    .X(net697));
 sg13g2_dlygate4sd3_1 hold425 (.A(_01043_),
    .X(net698));
 sg13g2_dlygate4sd3_1 hold426 (.A(\cordic_inst.cordic_state[34] ),
    .X(net699));
 sg13g2_dlygate4sd3_1 hold427 (.A(_00215_),
    .X(net700));
 sg13g2_dlygate4sd3_1 hold428 (.A(\cordic_inst.cordic_state[38] ),
    .X(net701));
 sg13g2_dlygate4sd3_1 hold429 (.A(_00219_),
    .X(net702));
 sg13g2_dlygate4sd3_1 hold430 (.A(\cordic_atan2_result[15] ),
    .X(net703));
 sg13g2_dlygate4sd3_1 hold431 (.A(\mac_inst.accumulator[22] ),
    .X(net704));
 sg13g2_dlygate4sd3_1 hold432 (.A(\cordic_inst.cordic_state[50] ),
    .X(net705));
 sg13g2_dlygate4sd3_1 hold433 (.A(_00231_),
    .X(net706));
 sg13g2_dlygate4sd3_1 hold434 (.A(\cordic_atan2_result[8] ),
    .X(net707));
 sg13g2_dlygate4sd3_1 hold435 (.A(_01003_),
    .X(net708));
 sg13g2_dlygate4sd3_1 hold436 (.A(\cordic_atan2_result[3] ),
    .X(net709));
 sg13g2_dlygate4sd3_1 hold437 (.A(_00954_),
    .X(net710));
 sg13g2_dlygate4sd3_1 hold438 (.A(\cordic_atan2_result[19] ),
    .X(net711));
 sg13g2_dlygate4sd3_1 hold439 (.A(\mac_inst.accumulator[16] ),
    .X(net712));
 sg13g2_dlygate4sd3_1 hold440 (.A(\mac_inst.accumulator[19] ),
    .X(net713));
 sg13g2_dlygate4sd3_1 hold441 (.A(_00406_),
    .X(net714));
 sg13g2_dlygate4sd3_1 hold442 (.A(\cmd_reg[0] ),
    .X(net715));
 sg13g2_dlygate4sd3_1 hold443 (.A(\cordic_inst.cordic_state[0] ),
    .X(net716));
 sg13g2_dlygate4sd3_1 hold444 (.A(_00183_),
    .X(net717));
 sg13g2_dlygate4sd3_1 hold445 (.A(\cmd_reg[2] ),
    .X(net718));
 sg13g2_dlygate4sd3_1 hold446 (.A(_00131_),
    .X(net719));
 sg13g2_dlygate4sd3_1 hold447 (.A(\mac_inst.accumulator[13] ),
    .X(net720));
 sg13g2_dlygate4sd3_1 hold448 (.A(\mac_inst.accumulator[5] ),
    .X(net721));
 sg13g2_dlygate4sd3_1 hold449 (.A(\cordic_inst.cordic_state[57] ),
    .X(net722));
 sg13g2_dlygate4sd3_1 hold450 (.A(_00238_),
    .X(net723));
 sg13g2_dlygate4sd3_1 hold451 (.A(\state[0] ),
    .X(net724));
 sg13g2_dlygate4sd3_1 hold452 (.A(_00126_),
    .X(net725));
 sg13g2_dlygate4sd3_1 hold453 (.A(\mac_inst.accumulator[2] ),
    .X(net726));
 sg13g2_dlygate4sd3_1 hold454 (.A(_05498_),
    .X(net727));
 sg13g2_dlygate4sd3_1 hold455 (.A(\cordic_atan2_result[9] ),
    .X(net728));
 sg13g2_dlygate4sd3_1 hold456 (.A(\cordic_inst.cordic_state[74] ),
    .X(net729));
 sg13g2_dlygate4sd3_1 hold457 (.A(_01922_),
    .X(net730));
 sg13g2_dlygate4sd3_1 hold458 (.A(\cordic_atan2_result[20] ),
    .X(net731));
 sg13g2_dlygate4sd3_1 hold459 (.A(\cordic_inst.cordic_state[43] ),
    .X(net732));
 sg13g2_dlygate4sd3_1 hold460 (.A(\mac_inst.accumulator[0] ),
    .X(net733));
 sg13g2_dlygate4sd3_1 hold461 (.A(_00387_),
    .X(net734));
 sg13g2_dlygate4sd3_1 hold462 (.A(\mac_inst.accumulator[1] ),
    .X(net735));
 sg13g2_dlygate4sd3_1 hold463 (.A(_05497_),
    .X(net736));
 sg13g2_dlygate4sd3_1 hold464 (.A(cordic_busy),
    .X(net737));
 sg13g2_dlygate4sd3_1 hold465 (.A(\cordic_atan2_result[23] ),
    .X(net738));
 sg13g2_dlygate4sd3_1 hold466 (.A(\cordic_inst.cordic_state[66] ),
    .X(net739));
 sg13g2_dlygate4sd3_1 hold467 (.A(_01802_),
    .X(net740));
 sg13g2_dlygate4sd3_1 hold468 (.A(\cordic_inst.cordic_state[72] ),
    .X(net741));
 sg13g2_dlygate4sd3_1 hold469 (.A(\cordic_inst.cordic_state[36] ),
    .X(net742));
 sg13g2_dlygate4sd3_1 hold470 (.A(\cordic_inst.cordic_state[45] ),
    .X(net743));
 sg13g2_dlygate4sd3_1 hold471 (.A(\cordic_inst.cordic_state[77] ),
    .X(net744));
 sg13g2_dlygate4sd3_1 hold472 (.A(_01964_),
    .X(net745));
 sg13g2_dlygate4sd3_1 hold473 (.A(\mac_inst.accumulator[11] ),
    .X(net746));
 sg13g2_dlygate4sd3_1 hold474 (.A(\mac_inst.accumulator[15] ),
    .X(net747));
 sg13g2_dlygate4sd3_1 hold475 (.A(_00402_),
    .X(net748));
 sg13g2_dlygate4sd3_1 hold476 (.A(\cordic_inst.cordic_state[61] ),
    .X(net749));
 sg13g2_dlygate4sd3_1 hold477 (.A(_00242_),
    .X(net750));
 sg13g2_dlygate4sd3_1 hold478 (.A(\cordic_inst.cordic_state[68] ),
    .X(net751));
 sg13g2_dlygate4sd3_1 hold479 (.A(\cordic_inst.cordic_state[70] ),
    .X(net752));
 sg13g2_dlygate4sd3_1 hold480 (.A(_00251_),
    .X(net753));
 sg13g2_dlygate4sd3_1 hold481 (.A(uo_out[7]),
    .X(net754));
 sg13g2_dlygate4sd3_1 hold482 (.A(_00748_),
    .X(net755));
 sg13g2_dlygate4sd3_1 hold483 (.A(_00125_),
    .X(net756));
 sg13g2_dlygate4sd3_1 hold484 (.A(\cordic_inst.cordic_state[37] ),
    .X(net757));
 sg13g2_dlygate4sd3_1 hold485 (.A(\cordic_inst.cordic_state[51] ),
    .X(net758));
 sg13g2_dlygate4sd3_1 hold486 (.A(_01513_),
    .X(net759));
 sg13g2_dlygate4sd3_1 hold487 (.A(\cordic_inst.cordic_state[71] ),
    .X(net760));
 sg13g2_dlygate4sd3_1 hold488 (.A(\state[0] ),
    .X(net761));
 sg13g2_dlygate4sd3_1 hold489 (.A(\cordic_inst.cordic_state[63] ),
    .X(net762));
 sg13g2_dlygate4sd3_1 hold490 (.A(_00244_),
    .X(net763));
 sg13g2_dlygate4sd3_1 hold491 (.A(\cordic_inst.cordic_state[56] ),
    .X(net764));
 sg13g2_dlygate4sd3_1 hold492 (.A(_00237_),
    .X(net765));
 sg13g2_dlygate4sd3_1 hold493 (.A(\cordic_atan2_result[21] ),
    .X(net766));
 sg13g2_dlygate4sd3_1 hold494 (.A(\cordic_inst.cordic_state[33] ),
    .X(net767));
 sg13g2_dlygate4sd3_1 hold495 (.A(\cordic_inst.cordic_state[65] ),
    .X(net768));
 sg13g2_dlygate4sd3_1 hold496 (.A(\cordic_inst.cordic_state[64] ),
    .X(net769));
 sg13g2_dlygate4sd3_1 hold497 (.A(_00245_),
    .X(net770));
 sg13g2_dlygate4sd3_1 hold498 (.A(\cordic_inst.cordic_state[49] ),
    .X(net771));
 sg13g2_dlygate4sd3_1 hold499 (.A(\byte_counter[3] ),
    .X(net772));
 sg13g2_dlygate4sd3_1 hold500 (.A(_00180_),
    .X(net773));
 sg13g2_dlygate4sd3_1 hold501 (.A(\byte_counter[1] ),
    .X(net774));
 sg13g2_dlygate4sd3_1 hold502 (.A(_00178_),
    .X(net775));
 sg13g2_dlygate4sd3_1 hold503 (.A(\cordic_atan2_result[1] ),
    .X(net776));
 sg13g2_dlygate4sd3_1 hold504 (.A(\cordic_inst.cordic_state[73] ),
    .X(net777));
 sg13g2_dlygate4sd3_1 hold505 (.A(_00254_),
    .X(net778));
 sg13g2_dlygate4sd3_1 hold506 (.A(\cordic_inst.cordic_state[58] ),
    .X(net779));
 sg13g2_dlygate4sd3_1 hold507 (.A(_00239_),
    .X(net780));
 sg13g2_dlygate4sd3_1 hold508 (.A(\cordic_inst.cordic_state[60] ),
    .X(net781));
 sg13g2_dlygate4sd3_1 hold509 (.A(\cordic_inst.cordic_state[78] ),
    .X(net782));
 sg13g2_dlygate4sd3_1 hold510 (.A(_00259_),
    .X(net783));
 sg13g2_dlygate4sd3_1 hold511 (.A(\cordic_inst.cordic_state[75] ),
    .X(net784));
 sg13g2_dlygate4sd3_1 hold512 (.A(_00256_),
    .X(net785));
 sg13g2_dlygate4sd3_1 hold513 (.A(\cordic_inst.cordic_state[32] ),
    .X(net786));
 sg13g2_dlygate4sd3_1 hold514 (.A(_00213_),
    .X(net787));
 sg13g2_dlygate4sd3_1 hold515 (.A(\mac_inst.accumulator[18] ),
    .X(net788));
 sg13g2_dlygate4sd3_1 hold516 (.A(\cmd_reg[6] ),
    .X(net789));
 sg13g2_dlygate4sd3_1 hold517 (.A(\exec_phase[2] ),
    .X(net790));
 sg13g2_dlygate4sd3_1 hold518 (.A(\cordic_inst.cordic_state[69] ),
    .X(net791));
 sg13g2_dlygate4sd3_1 hold519 (.A(\cordic_inst.MUX_cordic_state$write_1__VAL_1[55] ),
    .X(net792));
 sg13g2_dlygate4sd3_1 hold520 (.A(\cordic_inst.cordic_state[76] ),
    .X(net793));
 sg13g2_dlygate4sd3_1 hold521 (.A(_00257_),
    .X(net794));
 sg13g2_dlygate4sd3_1 hold522 (.A(\cordic_inst.MUX_cordic_state$write_1__VAL_1[68] ),
    .X(net795));
 sg13g2_dlygate4sd3_1 hold523 (.A(\mac_inst.accumulator[4] ),
    .X(net796));
 sg13g2_dlygate4sd3_1 hold524 (.A(\cordic_inst.cordic_state[55] ),
    .X(net797));
 sg13g2_dlygate4sd3_1 hold525 (.A(\cordic_inst.cordic_state[42] ),
    .X(net798));
 sg13g2_dlygate4sd3_1 hold526 (.A(_01379_),
    .X(net799));
 sg13g2_dlygate4sd3_1 hold527 (.A(\cordic_inst.MUX_cordic_state$write_1__VAL_1[62] ),
    .X(net800));
 sg13g2_dlygate4sd3_1 hold528 (.A(\cordic_inst.cordic_state[79] ),
    .X(net801));
 sg13g2_dlygate4sd3_1 hold529 (.A(\cordic_inst.cordic_state[44] ),
    .X(net802));
 sg13g2_dlygate4sd3_1 hold530 (.A(_01414_),
    .X(net803));
 sg13g2_dlygate4sd3_1 hold531 (.A(\state[2] ),
    .X(net804));
 sg13g2_dlygate4sd3_1 hold532 (.A(\mac_inst.accumulator[8] ),
    .X(net805));
 sg13g2_dlygate4sd3_1 hold533 (.A(wr_prev),
    .X(net806));
 sg13g2_dlygate4sd3_1 hold534 (.A(\cordic_inst.MUX_cordic_state$write_1__VAL_1[66] ),
    .X(net807));
 sg13g2_dlygate4sd3_1 hold535 (.A(\cordic_inst.MUX_cordic_state$write_1__VAL_1[37] ),
    .X(net808));
 sg13g2_dlygate4sd3_1 hold536 (.A(\cordic_inst.MUX_cordic_state$write_1__VAL_1[38] ),
    .X(net809));
 sg13g2_dlygate4sd3_1 hold537 (.A(\state[1] ),
    .X(net810));
 sg13g2_dlygate4sd3_1 hold538 (.A(\cordic_inst.MUX_cordic_state$write_1__VAL_1[57] ),
    .X(net811));
 sg13g2_dlygate4sd3_1 hold539 (.A(\cordic_inst.MUX_cordic_state$write_1__VAL_1[69] ),
    .X(net812));
 sg13g2_dlygate4sd3_1 hold540 (.A(\byte_counter[0] ),
    .X(net813));
 sg13g2_dlygate4sd3_1 hold541 (.A(\mac_inst.accumulator[10] ),
    .X(net814));
 sg13g2_dlygate4sd3_1 hold542 (.A(\cordic_inst.MUX_cordic_state$write_1__VAL_1[46] ),
    .X(net815));
 sg13g2_dlygate4sd3_1 hold543 (.A(\cordic_inst.MUX_cordic_state$write_1__VAL_1[67] ),
    .X(net816));
 sg13g2_dlygate4sd3_1 hold544 (.A(\cordic_inst.cordic_state[46] ),
    .X(net817));
 sg13g2_dlygate4sd3_1 hold545 (.A(\cordic_inst.cordic_state[54] ),
    .X(net818));
 sg13g2_dlygate4sd3_1 hold546 (.A(\mac_inst.accumulator[20] ),
    .X(net819));
 sg13g2_dlygate4sd3_1 hold547 (.A(\cordic_inst.cordic_state[67] ),
    .X(net820));
 sg13g2_dlygate4sd3_1 hold548 (.A(\cordic_inst.MUX_cordic_state$write_1__VAL_1[48] ),
    .X(net821));
 sg13g2_dlygate4sd3_1 hold549 (.A(\cordic_inst.MUX_cordic_state$write_1__VAL_1[39] ),
    .X(net822));
 sg13g2_dlygate4sd3_1 hold550 (.A(\cordic_inst.MUX_cordic_state$write_1__VAL_1[64] ),
    .X(net823));
 sg13g2_dlygate4sd3_1 hold551 (.A(\cmd_reg[5] ),
    .X(net824));
 sg13g2_dlygate4sd3_1 hold552 (.A(\cordic_inst.cordic_state[39] ),
    .X(net825));
 sg13g2_dlygate4sd3_1 hold553 (.A(\mac_inst.accumulator[7] ),
    .X(net826));
 sg13g2_dlygate4sd3_1 hold554 (.A(\mac_inst.accumulator[14] ),
    .X(net827));
 sg13g2_dlygate4sd3_1 hold555 (.A(\cordic_inst.cordic_state[40] ),
    .X(net828));
 sg13g2_dlygate4sd3_1 hold556 (.A(_00221_),
    .X(net829));
 sg13g2_dlygate4sd3_1 hold557 (.A(\mac_inst.accumulator[3] ),
    .X(net830));
 sg13g2_dlygate4sd3_1 hold558 (.A(\cordic_inst.MUX_cordic_state$write_1__VAL_1[75] ),
    .X(net831));
 sg13g2_dlygate4sd3_1 hold559 (.A(\cordic_inst.MUX_cordic_state$write_1__VAL_1[70] ),
    .X(net832));
 sg13g2_dlygate4sd3_1 hold560 (.A(\cordic_inst.cordic_state[53] ),
    .X(net833));
 sg13g2_dlygate4sd3_1 hold561 (.A(\cordic_inst.MUX_cordic_state$write_1__VAL_1[76] ),
    .X(net834));
 sg13g2_dlygate4sd3_1 hold562 (.A(\cordic_inst.MUX_cordic_state$write_1__VAL_1[53] ),
    .X(net835));
 sg13g2_dlygate4sd3_1 hold563 (.A(\mac_inst.accumulator[6] ),
    .X(net836));
 sg13g2_dlygate4sd3_1 hold564 (.A(\cordic_inst.MUX_cordic_state$write_1__VAL_1[54] ),
    .X(net837));
 sg13g2_dlygate4sd3_1 hold565 (.A(\cordic_inst.MUX_cordic_state$write_1__VAL_1[49] ),
    .X(net838));
 sg13g2_dlygate4sd3_1 hold566 (.A(\cordic_inst.MUX_cordic_state$write_1__VAL_1[35] ),
    .X(net839));
 sg13g2_dlygate4sd3_1 hold567 (.A(\cordic_inst.MUX_cordic_state$write_1__VAL_1[61] ),
    .X(net840));
 sg13g2_dlygate4sd3_1 hold568 (.A(\cordic_inst.MUX_cordic_state$write_1__VAL_1[63] ),
    .X(net841));
 sg13g2_dlygate4sd3_1 hold569 (.A(\cordic_inst.cordic_state[47] ),
    .X(net842));
 sg13g2_dlygate4sd3_1 hold570 (.A(\cordic_inst.MUX_cordic_state$write_1__VAL_1[34] ),
    .X(net843));
 sg13g2_dlygate4sd3_1 hold571 (.A(\cordic_inst.MUX_cordic_state$write_1__VAL_1[74] ),
    .X(net844));
 sg13g2_dlygate4sd3_1 hold572 (.A(\cordic_inst.MUX_cordic_state$write_1__VAL_1[52] ),
    .X(net845));
 sg13g2_dlygate4sd3_1 hold573 (.A(\cordic_inst.MUX_cordic_state$write_1__VAL_1[43] ),
    .X(net846));
 sg13g2_dlygate4sd3_1 hold574 (.A(\cordic_inst.MUX_cordic_state$write_1__VAL_1[78] ),
    .X(net847));
 sg13g2_dlygate4sd3_1 hold575 (.A(\cordic_inst.MUX_cordic_state$write_1__VAL_1[50] ),
    .X(net848));
 sg13g2_dlygate4sd3_1 hold576 (.A(\cordic_inst.MUX_cordic_state$write_1__VAL_1[42] ),
    .X(net849));
 sg13g2_dlygate4sd3_1 hold577 (.A(\cordic_inst.MUX_cordic_state$write_1__VAL_1[41] ),
    .X(net850));
 sg13g2_dlygate4sd3_1 hold578 (.A(\cordic_inst.MUX_cordic_state$write_1__VAL_1[40] ),
    .X(net851));
 sg13g2_dlygate4sd3_1 hold579 (.A(\cordic_inst.MUX_cordic_state$write_1__VAL_1[47] ),
    .X(net852));
 sg13g2_dlygate4sd3_1 hold580 (.A(\cordic_inst.MUX_cordic_state$write_1__VAL_1[60] ),
    .X(net853));
 sg13g2_dlygate4sd3_1 hold581 (.A(\cordic_inst.MUX_cordic_state$write_1__VAL_1[44] ),
    .X(net854));
 sg13g2_dlygate4sd3_1 hold582 (.A(\cordic_inst.MUX_cordic_state$write_1__VAL_1[73] ),
    .X(net855));
 sg13g2_dlygate4sd3_1 hold583 (.A(\cordic_inst.MUX_cordic_state$write_1__VAL_1[51] ),
    .X(net856));
 sg13g2_dlygate4sd3_1 hold584 (.A(\cordic_inst.MUX_cordic_state$write_1__VAL_1[36] ),
    .X(net857));
 sg13g2_dlygate4sd3_1 hold585 (.A(\cordic_inst.MUX_cordic_state$write_1__VAL_1[45] ),
    .X(net858));
 sg13g2_dlygate4sd3_1 hold586 (.A(\cordic_inst.MUX_cordic_state$write_1__VAL_1[32] ),
    .X(net859));
 sg13g2_dlygate4sd3_1 hold587 (.A(\cordic_inst.cordic_state[6] ),
    .X(net860));
 sg13g2_dlygate4sd3_1 hold588 (.A(\cordic_inst.MUX_cordic_state$write_1__VAL_1[63] ),
    .X(net861));
 sg13g2_antennanp ANTENNA_1 (.A(_01990_));
 sg13g2_antennanp ANTENNA_2 (.A(_01990_));
 sg13g2_antennanp ANTENNA_3 (.A(_05493_));
 sg13g2_antennanp ANTENNA_4 (.A(_05612_));
 sg13g2_antennanp ANTENNA_5 (.A(_05660_));
 sg13g2_antennanp ANTENNA_6 (.A(\mac_inst.RDY_get_multiply ));
 sg13g2_antennanp ANTENNA_7 (.A(uio_in[0]));
 sg13g2_antennanp ANTENNA_8 (.A(uio_in[1]));
 sg13g2_antennanp ANTENNA_9 (.A(net1211));
 sg13g2_antennanp ANTENNA_10 (.A(net1211));
 sg13g2_antennanp ANTENNA_11 (.A(net1211));
 sg13g2_antennanp ANTENNA_12 (.A(net1211));
 sg13g2_antennanp ANTENNA_13 (.A(net1212));
 sg13g2_antennanp ANTENNA_14 (.A(net1212));
 sg13g2_antennanp ANTENNA_15 (.A(net1212));
 sg13g2_antennanp ANTENNA_16 (.A(net1212));
 sg13g2_antennanp ANTENNA_17 (.A(net1254));
 sg13g2_antennanp ANTENNA_18 (.A(net1254));
 sg13g2_antennanp ANTENNA_19 (.A(net1313));
 sg13g2_antennanp ANTENNA_20 (.A(net1313));
 sg13g2_antennanp ANTENNA_21 (.A(net274));
 sg13g2_antennanp ANTENNA_22 (.A(net278));
 sg13g2_antennanp ANTENNA_23 (.A(net483));
 sg13g2_antennanp ANTENNA_24 (.A(net662));
 sg13g2_antennanp ANTENNA_25 (.A(_00015_));
 sg13g2_antennanp ANTENNA_26 (.A(_00477_));
 sg13g2_antennanp ANTENNA_27 (.A(cordic_busy));
 sg13g2_antennanp ANTENNA_28 (.A(net635));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_fill_2 FILLER_0_126 ();
 sg13g2_fill_1 FILLER_0_128 ();
 sg13g2_fill_1 FILLER_0_188 ();
 sg13g2_fill_1 FILLER_0_217 ();
 sg13g2_fill_2 FILLER_0_317 ();
 sg13g2_fill_1 FILLER_0_319 ();
 sg13g2_fill_2 FILLER_0_338 ();
 sg13g2_fill_1 FILLER_0_340 ();
 sg13g2_fill_1 FILLER_0_351 ();
 sg13g2_fill_2 FILLER_0_370 ();
 sg13g2_fill_1 FILLER_0_407 ();
 sg13g2_fill_1 FILLER_0_412 ();
 sg13g2_decap_8 FILLER_0_445 ();
 sg13g2_decap_8 FILLER_0_452 ();
 sg13g2_decap_8 FILLER_0_459 ();
 sg13g2_fill_1 FILLER_0_466 ();
 sg13g2_decap_8 FILLER_0_471 ();
 sg13g2_decap_8 FILLER_0_478 ();
 sg13g2_decap_8 FILLER_0_485 ();
 sg13g2_decap_8 FILLER_0_492 ();
 sg13g2_decap_8 FILLER_0_499 ();
 sg13g2_decap_8 FILLER_0_506 ();
 sg13g2_decap_8 FILLER_0_513 ();
 sg13g2_decap_8 FILLER_0_520 ();
 sg13g2_decap_8 FILLER_0_527 ();
 sg13g2_decap_8 FILLER_0_534 ();
 sg13g2_decap_8 FILLER_0_541 ();
 sg13g2_decap_8 FILLER_0_548 ();
 sg13g2_decap_8 FILLER_0_555 ();
 sg13g2_decap_8 FILLER_0_562 ();
 sg13g2_decap_8 FILLER_0_569 ();
 sg13g2_decap_8 FILLER_0_576 ();
 sg13g2_decap_8 FILLER_0_583 ();
 sg13g2_decap_8 FILLER_0_590 ();
 sg13g2_decap_8 FILLER_0_597 ();
 sg13g2_decap_8 FILLER_0_604 ();
 sg13g2_decap_8 FILLER_0_611 ();
 sg13g2_decap_8 FILLER_0_618 ();
 sg13g2_decap_8 FILLER_0_625 ();
 sg13g2_decap_8 FILLER_0_632 ();
 sg13g2_decap_8 FILLER_0_639 ();
 sg13g2_decap_8 FILLER_0_646 ();
 sg13g2_decap_8 FILLER_0_653 ();
 sg13g2_decap_8 FILLER_0_660 ();
 sg13g2_decap_8 FILLER_0_667 ();
 sg13g2_decap_8 FILLER_0_674 ();
 sg13g2_decap_8 FILLER_0_681 ();
 sg13g2_decap_8 FILLER_0_688 ();
 sg13g2_decap_8 FILLER_0_695 ();
 sg13g2_decap_8 FILLER_0_702 ();
 sg13g2_decap_8 FILLER_0_709 ();
 sg13g2_decap_8 FILLER_0_716 ();
 sg13g2_decap_8 FILLER_0_723 ();
 sg13g2_decap_8 FILLER_0_730 ();
 sg13g2_decap_8 FILLER_0_737 ();
 sg13g2_decap_8 FILLER_0_744 ();
 sg13g2_decap_8 FILLER_0_751 ();
 sg13g2_decap_8 FILLER_0_758 ();
 sg13g2_decap_8 FILLER_0_765 ();
 sg13g2_decap_8 FILLER_0_772 ();
 sg13g2_decap_8 FILLER_0_779 ();
 sg13g2_decap_8 FILLER_0_786 ();
 sg13g2_decap_8 FILLER_0_793 ();
 sg13g2_decap_8 FILLER_0_800 ();
 sg13g2_decap_8 FILLER_0_807 ();
 sg13g2_decap_8 FILLER_0_814 ();
 sg13g2_decap_8 FILLER_0_821 ();
 sg13g2_decap_8 FILLER_0_828 ();
 sg13g2_decap_8 FILLER_0_835 ();
 sg13g2_decap_8 FILLER_0_842 ();
 sg13g2_decap_8 FILLER_0_849 ();
 sg13g2_decap_4 FILLER_0_856 ();
 sg13g2_fill_2 FILLER_0_860 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_fill_2 FILLER_1_112 ();
 sg13g2_fill_2 FILLER_1_166 ();
 sg13g2_fill_2 FILLER_1_208 ();
 sg13g2_fill_1 FILLER_1_210 ();
 sg13g2_fill_2 FILLER_1_239 ();
 sg13g2_fill_2 FILLER_1_254 ();
 sg13g2_fill_2 FILLER_1_386 ();
 sg13g2_fill_2 FILLER_1_397 ();
 sg13g2_fill_2 FILLER_1_456 ();
 sg13g2_decap_8 FILLER_1_475 ();
 sg13g2_decap_8 FILLER_1_482 ();
 sg13g2_decap_8 FILLER_1_489 ();
 sg13g2_decap_8 FILLER_1_496 ();
 sg13g2_decap_4 FILLER_1_503 ();
 sg13g2_fill_2 FILLER_1_507 ();
 sg13g2_decap_8 FILLER_1_513 ();
 sg13g2_decap_8 FILLER_1_520 ();
 sg13g2_decap_8 FILLER_1_527 ();
 sg13g2_decap_8 FILLER_1_534 ();
 sg13g2_decap_8 FILLER_1_541 ();
 sg13g2_decap_8 FILLER_1_548 ();
 sg13g2_decap_8 FILLER_1_555 ();
 sg13g2_decap_8 FILLER_1_562 ();
 sg13g2_decap_8 FILLER_1_569 ();
 sg13g2_decap_8 FILLER_1_576 ();
 sg13g2_decap_8 FILLER_1_583 ();
 sg13g2_decap_8 FILLER_1_590 ();
 sg13g2_decap_8 FILLER_1_597 ();
 sg13g2_decap_8 FILLER_1_604 ();
 sg13g2_decap_8 FILLER_1_611 ();
 sg13g2_decap_8 FILLER_1_618 ();
 sg13g2_decap_8 FILLER_1_625 ();
 sg13g2_decap_8 FILLER_1_632 ();
 sg13g2_decap_8 FILLER_1_639 ();
 sg13g2_decap_8 FILLER_1_646 ();
 sg13g2_decap_8 FILLER_1_653 ();
 sg13g2_decap_8 FILLER_1_660 ();
 sg13g2_decap_8 FILLER_1_667 ();
 sg13g2_decap_8 FILLER_1_674 ();
 sg13g2_decap_8 FILLER_1_681 ();
 sg13g2_decap_8 FILLER_1_688 ();
 sg13g2_decap_8 FILLER_1_695 ();
 sg13g2_decap_8 FILLER_1_702 ();
 sg13g2_decap_8 FILLER_1_709 ();
 sg13g2_decap_8 FILLER_1_716 ();
 sg13g2_decap_8 FILLER_1_723 ();
 sg13g2_decap_8 FILLER_1_730 ();
 sg13g2_decap_8 FILLER_1_737 ();
 sg13g2_decap_8 FILLER_1_744 ();
 sg13g2_decap_8 FILLER_1_751 ();
 sg13g2_decap_8 FILLER_1_758 ();
 sg13g2_decap_8 FILLER_1_765 ();
 sg13g2_decap_8 FILLER_1_772 ();
 sg13g2_decap_8 FILLER_1_779 ();
 sg13g2_decap_8 FILLER_1_786 ();
 sg13g2_decap_8 FILLER_1_793 ();
 sg13g2_decap_8 FILLER_1_800 ();
 sg13g2_decap_8 FILLER_1_807 ();
 sg13g2_decap_8 FILLER_1_814 ();
 sg13g2_decap_8 FILLER_1_821 ();
 sg13g2_decap_8 FILLER_1_828 ();
 sg13g2_decap_8 FILLER_1_835 ();
 sg13g2_decap_8 FILLER_1_842 ();
 sg13g2_decap_8 FILLER_1_849 ();
 sg13g2_decap_4 FILLER_1_856 ();
 sg13g2_fill_2 FILLER_1_860 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_4 FILLER_2_105 ();
 sg13g2_fill_1 FILLER_2_109 ();
 sg13g2_fill_2 FILLER_2_153 ();
 sg13g2_fill_1 FILLER_2_164 ();
 sg13g2_fill_1 FILLER_2_213 ();
 sg13g2_fill_1 FILLER_2_298 ();
 sg13g2_fill_1 FILLER_2_304 ();
 sg13g2_fill_1 FILLER_2_355 ();
 sg13g2_fill_2 FILLER_2_406 ();
 sg13g2_fill_2 FILLER_2_486 ();
 sg13g2_fill_1 FILLER_2_488 ();
 sg13g2_fill_1 FILLER_2_509 ();
 sg13g2_fill_2 FILLER_2_514 ();
 sg13g2_fill_1 FILLER_2_516 ();
 sg13g2_decap_8 FILLER_2_526 ();
 sg13g2_decap_4 FILLER_2_533 ();
 sg13g2_fill_2 FILLER_2_537 ();
 sg13g2_decap_8 FILLER_2_543 ();
 sg13g2_decap_8 FILLER_2_550 ();
 sg13g2_decap_8 FILLER_2_557 ();
 sg13g2_decap_8 FILLER_2_564 ();
 sg13g2_decap_8 FILLER_2_571 ();
 sg13g2_decap_8 FILLER_2_578 ();
 sg13g2_decap_8 FILLER_2_585 ();
 sg13g2_decap_8 FILLER_2_592 ();
 sg13g2_decap_8 FILLER_2_599 ();
 sg13g2_decap_8 FILLER_2_606 ();
 sg13g2_decap_8 FILLER_2_613 ();
 sg13g2_decap_8 FILLER_2_620 ();
 sg13g2_decap_8 FILLER_2_627 ();
 sg13g2_decap_8 FILLER_2_634 ();
 sg13g2_decap_8 FILLER_2_641 ();
 sg13g2_decap_8 FILLER_2_648 ();
 sg13g2_decap_8 FILLER_2_655 ();
 sg13g2_decap_8 FILLER_2_662 ();
 sg13g2_decap_8 FILLER_2_669 ();
 sg13g2_decap_8 FILLER_2_676 ();
 sg13g2_decap_8 FILLER_2_683 ();
 sg13g2_decap_8 FILLER_2_690 ();
 sg13g2_decap_8 FILLER_2_697 ();
 sg13g2_decap_8 FILLER_2_704 ();
 sg13g2_decap_8 FILLER_2_711 ();
 sg13g2_decap_8 FILLER_2_718 ();
 sg13g2_decap_8 FILLER_2_725 ();
 sg13g2_decap_8 FILLER_2_732 ();
 sg13g2_decap_8 FILLER_2_739 ();
 sg13g2_decap_8 FILLER_2_746 ();
 sg13g2_decap_8 FILLER_2_753 ();
 sg13g2_decap_8 FILLER_2_760 ();
 sg13g2_decap_8 FILLER_2_767 ();
 sg13g2_decap_8 FILLER_2_774 ();
 sg13g2_decap_8 FILLER_2_781 ();
 sg13g2_decap_8 FILLER_2_788 ();
 sg13g2_decap_8 FILLER_2_795 ();
 sg13g2_decap_8 FILLER_2_802 ();
 sg13g2_decap_8 FILLER_2_809 ();
 sg13g2_decap_8 FILLER_2_816 ();
 sg13g2_decap_8 FILLER_2_823 ();
 sg13g2_decap_8 FILLER_2_830 ();
 sg13g2_decap_8 FILLER_2_837 ();
 sg13g2_decap_8 FILLER_2_844 ();
 sg13g2_decap_8 FILLER_2_851 ();
 sg13g2_decap_4 FILLER_2_858 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_4 FILLER_3_91 ();
 sg13g2_fill_2 FILLER_3_95 ();
 sg13g2_fill_2 FILLER_3_130 ();
 sg13g2_fill_1 FILLER_3_132 ();
 sg13g2_fill_2 FILLER_3_151 ();
 sg13g2_fill_1 FILLER_3_163 ();
 sg13g2_fill_2 FILLER_3_169 ();
 sg13g2_fill_1 FILLER_3_171 ();
 sg13g2_fill_1 FILLER_3_197 ();
 sg13g2_fill_1 FILLER_3_229 ();
 sg13g2_fill_1 FILLER_3_245 ();
 sg13g2_fill_2 FILLER_3_251 ();
 sg13g2_fill_1 FILLER_3_275 ();
 sg13g2_fill_2 FILLER_3_286 ();
 sg13g2_fill_2 FILLER_3_336 ();
 sg13g2_fill_2 FILLER_3_386 ();
 sg13g2_fill_1 FILLER_3_402 ();
 sg13g2_fill_1 FILLER_3_408 ();
 sg13g2_fill_2 FILLER_3_449 ();
 sg13g2_fill_2 FILLER_3_471 ();
 sg13g2_fill_1 FILLER_3_473 ();
 sg13g2_fill_2 FILLER_3_502 ();
 sg13g2_decap_8 FILLER_3_558 ();
 sg13g2_decap_8 FILLER_3_565 ();
 sg13g2_decap_8 FILLER_3_572 ();
 sg13g2_decap_8 FILLER_3_579 ();
 sg13g2_decap_8 FILLER_3_586 ();
 sg13g2_decap_8 FILLER_3_593 ();
 sg13g2_decap_8 FILLER_3_600 ();
 sg13g2_decap_8 FILLER_3_607 ();
 sg13g2_decap_8 FILLER_3_614 ();
 sg13g2_decap_8 FILLER_3_621 ();
 sg13g2_decap_8 FILLER_3_628 ();
 sg13g2_decap_8 FILLER_3_635 ();
 sg13g2_decap_8 FILLER_3_642 ();
 sg13g2_decap_8 FILLER_3_649 ();
 sg13g2_decap_8 FILLER_3_656 ();
 sg13g2_decap_8 FILLER_3_663 ();
 sg13g2_decap_8 FILLER_3_670 ();
 sg13g2_decap_8 FILLER_3_677 ();
 sg13g2_decap_8 FILLER_3_684 ();
 sg13g2_decap_8 FILLER_3_691 ();
 sg13g2_decap_8 FILLER_3_698 ();
 sg13g2_decap_8 FILLER_3_705 ();
 sg13g2_decap_8 FILLER_3_712 ();
 sg13g2_decap_8 FILLER_3_719 ();
 sg13g2_decap_8 FILLER_3_726 ();
 sg13g2_decap_8 FILLER_3_733 ();
 sg13g2_decap_8 FILLER_3_740 ();
 sg13g2_decap_8 FILLER_3_747 ();
 sg13g2_decap_8 FILLER_3_754 ();
 sg13g2_decap_8 FILLER_3_761 ();
 sg13g2_decap_8 FILLER_3_768 ();
 sg13g2_decap_8 FILLER_3_775 ();
 sg13g2_decap_8 FILLER_3_782 ();
 sg13g2_decap_8 FILLER_3_789 ();
 sg13g2_decap_8 FILLER_3_796 ();
 sg13g2_decap_8 FILLER_3_803 ();
 sg13g2_decap_8 FILLER_3_810 ();
 sg13g2_decap_8 FILLER_3_817 ();
 sg13g2_decap_8 FILLER_3_824 ();
 sg13g2_decap_8 FILLER_3_831 ();
 sg13g2_decap_8 FILLER_3_838 ();
 sg13g2_decap_8 FILLER_3_845 ();
 sg13g2_decap_8 FILLER_3_852 ();
 sg13g2_fill_2 FILLER_3_859 ();
 sg13g2_fill_1 FILLER_3_861 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_4 FILLER_4_98 ();
 sg13g2_fill_1 FILLER_4_158 ();
 sg13g2_fill_2 FILLER_4_179 ();
 sg13g2_fill_1 FILLER_4_259 ();
 sg13g2_fill_2 FILLER_4_285 ();
 sg13g2_fill_1 FILLER_4_292 ();
 sg13g2_fill_2 FILLER_4_321 ();
 sg13g2_fill_1 FILLER_4_397 ();
 sg13g2_fill_1 FILLER_4_441 ();
 sg13g2_fill_1 FILLER_4_475 ();
 sg13g2_fill_2 FILLER_4_493 ();
 sg13g2_fill_1 FILLER_4_534 ();
 sg13g2_fill_1 FILLER_4_552 ();
 sg13g2_decap_8 FILLER_4_566 ();
 sg13g2_decap_8 FILLER_4_573 ();
 sg13g2_decap_8 FILLER_4_580 ();
 sg13g2_decap_8 FILLER_4_587 ();
 sg13g2_decap_8 FILLER_4_594 ();
 sg13g2_decap_8 FILLER_4_601 ();
 sg13g2_decap_8 FILLER_4_608 ();
 sg13g2_decap_8 FILLER_4_615 ();
 sg13g2_decap_8 FILLER_4_622 ();
 sg13g2_decap_8 FILLER_4_629 ();
 sg13g2_decap_8 FILLER_4_636 ();
 sg13g2_decap_8 FILLER_4_643 ();
 sg13g2_decap_8 FILLER_4_650 ();
 sg13g2_decap_8 FILLER_4_657 ();
 sg13g2_decap_8 FILLER_4_664 ();
 sg13g2_decap_8 FILLER_4_671 ();
 sg13g2_decap_8 FILLER_4_678 ();
 sg13g2_decap_8 FILLER_4_685 ();
 sg13g2_decap_8 FILLER_4_692 ();
 sg13g2_decap_8 FILLER_4_699 ();
 sg13g2_decap_8 FILLER_4_706 ();
 sg13g2_decap_8 FILLER_4_713 ();
 sg13g2_decap_8 FILLER_4_720 ();
 sg13g2_decap_8 FILLER_4_727 ();
 sg13g2_decap_8 FILLER_4_734 ();
 sg13g2_decap_8 FILLER_4_741 ();
 sg13g2_decap_8 FILLER_4_748 ();
 sg13g2_decap_8 FILLER_4_755 ();
 sg13g2_decap_8 FILLER_4_762 ();
 sg13g2_decap_8 FILLER_4_769 ();
 sg13g2_decap_8 FILLER_4_776 ();
 sg13g2_decap_8 FILLER_4_783 ();
 sg13g2_decap_8 FILLER_4_790 ();
 sg13g2_decap_8 FILLER_4_797 ();
 sg13g2_decap_8 FILLER_4_804 ();
 sg13g2_decap_8 FILLER_4_811 ();
 sg13g2_decap_8 FILLER_4_818 ();
 sg13g2_decap_8 FILLER_4_825 ();
 sg13g2_decap_8 FILLER_4_832 ();
 sg13g2_decap_8 FILLER_4_839 ();
 sg13g2_decap_8 FILLER_4_846 ();
 sg13g2_decap_8 FILLER_4_853 ();
 sg13g2_fill_2 FILLER_4_860 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_fill_2 FILLER_5_91 ();
 sg13g2_fill_1 FILLER_5_93 ();
 sg13g2_fill_1 FILLER_5_129 ();
 sg13g2_fill_1 FILLER_5_171 ();
 sg13g2_fill_2 FILLER_5_177 ();
 sg13g2_fill_2 FILLER_5_189 ();
 sg13g2_fill_1 FILLER_5_252 ();
 sg13g2_fill_2 FILLER_5_314 ();
 sg13g2_fill_2 FILLER_5_388 ();
 sg13g2_fill_1 FILLER_5_404 ();
 sg13g2_fill_2 FILLER_5_415 ();
 sg13g2_fill_2 FILLER_5_435 ();
 sg13g2_fill_2 FILLER_5_466 ();
 sg13g2_fill_1 FILLER_5_468 ();
 sg13g2_decap_8 FILLER_5_570 ();
 sg13g2_decap_8 FILLER_5_577 ();
 sg13g2_decap_8 FILLER_5_584 ();
 sg13g2_decap_8 FILLER_5_591 ();
 sg13g2_decap_8 FILLER_5_598 ();
 sg13g2_decap_8 FILLER_5_605 ();
 sg13g2_decap_8 FILLER_5_612 ();
 sg13g2_decap_8 FILLER_5_619 ();
 sg13g2_decap_8 FILLER_5_626 ();
 sg13g2_decap_8 FILLER_5_633 ();
 sg13g2_decap_8 FILLER_5_640 ();
 sg13g2_decap_8 FILLER_5_647 ();
 sg13g2_decap_8 FILLER_5_654 ();
 sg13g2_decap_8 FILLER_5_661 ();
 sg13g2_decap_8 FILLER_5_668 ();
 sg13g2_decap_8 FILLER_5_675 ();
 sg13g2_decap_8 FILLER_5_682 ();
 sg13g2_decap_8 FILLER_5_689 ();
 sg13g2_decap_8 FILLER_5_696 ();
 sg13g2_decap_8 FILLER_5_703 ();
 sg13g2_decap_8 FILLER_5_710 ();
 sg13g2_decap_8 FILLER_5_717 ();
 sg13g2_decap_8 FILLER_5_724 ();
 sg13g2_decap_8 FILLER_5_731 ();
 sg13g2_decap_8 FILLER_5_738 ();
 sg13g2_decap_8 FILLER_5_745 ();
 sg13g2_decap_8 FILLER_5_752 ();
 sg13g2_decap_8 FILLER_5_759 ();
 sg13g2_decap_8 FILLER_5_766 ();
 sg13g2_decap_8 FILLER_5_773 ();
 sg13g2_decap_8 FILLER_5_780 ();
 sg13g2_decap_8 FILLER_5_787 ();
 sg13g2_decap_8 FILLER_5_794 ();
 sg13g2_decap_8 FILLER_5_801 ();
 sg13g2_decap_8 FILLER_5_808 ();
 sg13g2_decap_8 FILLER_5_815 ();
 sg13g2_decap_8 FILLER_5_822 ();
 sg13g2_decap_8 FILLER_5_829 ();
 sg13g2_decap_8 FILLER_5_836 ();
 sg13g2_decap_8 FILLER_5_843 ();
 sg13g2_decap_8 FILLER_5_850 ();
 sg13g2_decap_4 FILLER_5_857 ();
 sg13g2_fill_1 FILLER_5_861 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_fill_2 FILLER_6_91 ();
 sg13g2_fill_1 FILLER_6_152 ();
 sg13g2_fill_2 FILLER_6_175 ();
 sg13g2_fill_1 FILLER_6_206 ();
 sg13g2_fill_1 FILLER_6_237 ();
 sg13g2_fill_1 FILLER_6_315 ();
 sg13g2_fill_2 FILLER_6_361 ();
 sg13g2_fill_2 FILLER_6_407 ();
 sg13g2_fill_1 FILLER_6_432 ();
 sg13g2_fill_1 FILLER_6_523 ();
 sg13g2_fill_2 FILLER_6_529 ();
 sg13g2_fill_1 FILLER_6_539 ();
 sg13g2_fill_1 FILLER_6_549 ();
 sg13g2_decap_8 FILLER_6_578 ();
 sg13g2_decap_8 FILLER_6_585 ();
 sg13g2_decap_8 FILLER_6_592 ();
 sg13g2_decap_8 FILLER_6_599 ();
 sg13g2_decap_8 FILLER_6_606 ();
 sg13g2_decap_8 FILLER_6_613 ();
 sg13g2_decap_8 FILLER_6_620 ();
 sg13g2_decap_8 FILLER_6_627 ();
 sg13g2_decap_8 FILLER_6_634 ();
 sg13g2_decap_8 FILLER_6_641 ();
 sg13g2_decap_8 FILLER_6_648 ();
 sg13g2_decap_8 FILLER_6_655 ();
 sg13g2_decap_8 FILLER_6_662 ();
 sg13g2_decap_8 FILLER_6_669 ();
 sg13g2_decap_8 FILLER_6_676 ();
 sg13g2_decap_8 FILLER_6_683 ();
 sg13g2_decap_8 FILLER_6_690 ();
 sg13g2_decap_8 FILLER_6_697 ();
 sg13g2_decap_8 FILLER_6_704 ();
 sg13g2_decap_8 FILLER_6_711 ();
 sg13g2_decap_8 FILLER_6_718 ();
 sg13g2_decap_8 FILLER_6_725 ();
 sg13g2_decap_8 FILLER_6_732 ();
 sg13g2_decap_8 FILLER_6_739 ();
 sg13g2_decap_8 FILLER_6_746 ();
 sg13g2_decap_8 FILLER_6_753 ();
 sg13g2_decap_8 FILLER_6_760 ();
 sg13g2_decap_8 FILLER_6_767 ();
 sg13g2_decap_8 FILLER_6_774 ();
 sg13g2_decap_8 FILLER_6_781 ();
 sg13g2_decap_8 FILLER_6_788 ();
 sg13g2_decap_8 FILLER_6_795 ();
 sg13g2_decap_8 FILLER_6_802 ();
 sg13g2_decap_8 FILLER_6_809 ();
 sg13g2_decap_8 FILLER_6_816 ();
 sg13g2_decap_8 FILLER_6_823 ();
 sg13g2_decap_8 FILLER_6_830 ();
 sg13g2_decap_8 FILLER_6_837 ();
 sg13g2_decap_8 FILLER_6_844 ();
 sg13g2_decap_8 FILLER_6_851 ();
 sg13g2_decap_4 FILLER_6_858 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_fill_2 FILLER_7_138 ();
 sg13g2_fill_1 FILLER_7_168 ();
 sg13g2_fill_2 FILLER_7_255 ();
 sg13g2_fill_2 FILLER_7_298 ();
 sg13g2_fill_1 FILLER_7_374 ();
 sg13g2_fill_2 FILLER_7_456 ();
 sg13g2_fill_1 FILLER_7_458 ();
 sg13g2_fill_2 FILLER_7_463 ();
 sg13g2_fill_1 FILLER_7_478 ();
 sg13g2_fill_2 FILLER_7_484 ();
 sg13g2_fill_1 FILLER_7_486 ();
 sg13g2_fill_2 FILLER_7_529 ();
 sg13g2_decap_8 FILLER_7_569 ();
 sg13g2_decap_8 FILLER_7_576 ();
 sg13g2_decap_8 FILLER_7_583 ();
 sg13g2_decap_8 FILLER_7_590 ();
 sg13g2_decap_8 FILLER_7_597 ();
 sg13g2_decap_8 FILLER_7_604 ();
 sg13g2_decap_8 FILLER_7_611 ();
 sg13g2_decap_8 FILLER_7_618 ();
 sg13g2_decap_8 FILLER_7_625 ();
 sg13g2_decap_8 FILLER_7_632 ();
 sg13g2_decap_8 FILLER_7_639 ();
 sg13g2_decap_8 FILLER_7_646 ();
 sg13g2_decap_8 FILLER_7_653 ();
 sg13g2_decap_8 FILLER_7_660 ();
 sg13g2_decap_8 FILLER_7_667 ();
 sg13g2_decap_8 FILLER_7_674 ();
 sg13g2_decap_8 FILLER_7_681 ();
 sg13g2_decap_8 FILLER_7_688 ();
 sg13g2_decap_8 FILLER_7_695 ();
 sg13g2_decap_8 FILLER_7_702 ();
 sg13g2_decap_8 FILLER_7_709 ();
 sg13g2_decap_8 FILLER_7_716 ();
 sg13g2_decap_8 FILLER_7_723 ();
 sg13g2_decap_8 FILLER_7_730 ();
 sg13g2_decap_8 FILLER_7_737 ();
 sg13g2_decap_8 FILLER_7_744 ();
 sg13g2_decap_8 FILLER_7_751 ();
 sg13g2_decap_8 FILLER_7_758 ();
 sg13g2_decap_8 FILLER_7_765 ();
 sg13g2_decap_8 FILLER_7_772 ();
 sg13g2_decap_8 FILLER_7_779 ();
 sg13g2_decap_8 FILLER_7_786 ();
 sg13g2_decap_8 FILLER_7_793 ();
 sg13g2_decap_8 FILLER_7_800 ();
 sg13g2_decap_8 FILLER_7_807 ();
 sg13g2_decap_8 FILLER_7_814 ();
 sg13g2_decap_8 FILLER_7_821 ();
 sg13g2_decap_8 FILLER_7_828 ();
 sg13g2_decap_8 FILLER_7_835 ();
 sg13g2_decap_8 FILLER_7_842 ();
 sg13g2_decap_8 FILLER_7_849 ();
 sg13g2_decap_4 FILLER_7_856 ();
 sg13g2_fill_2 FILLER_7_860 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_4 FILLER_8_91 ();
 sg13g2_fill_2 FILLER_8_95 ();
 sg13g2_fill_1 FILLER_8_122 ();
 sg13g2_fill_1 FILLER_8_132 ();
 sg13g2_fill_2 FILLER_8_155 ();
 sg13g2_fill_1 FILLER_8_157 ();
 sg13g2_fill_1 FILLER_8_220 ();
 sg13g2_fill_2 FILLER_8_269 ();
 sg13g2_fill_1 FILLER_8_422 ();
 sg13g2_fill_1 FILLER_8_521 ();
 sg13g2_decap_8 FILLER_8_573 ();
 sg13g2_decap_8 FILLER_8_580 ();
 sg13g2_decap_8 FILLER_8_587 ();
 sg13g2_decap_8 FILLER_8_594 ();
 sg13g2_decap_8 FILLER_8_601 ();
 sg13g2_decap_8 FILLER_8_608 ();
 sg13g2_decap_8 FILLER_8_615 ();
 sg13g2_decap_4 FILLER_8_622 ();
 sg13g2_fill_1 FILLER_8_626 ();
 sg13g2_decap_8 FILLER_8_644 ();
 sg13g2_decap_4 FILLER_8_651 ();
 sg13g2_fill_2 FILLER_8_655 ();
 sg13g2_decap_8 FILLER_8_662 ();
 sg13g2_decap_8 FILLER_8_669 ();
 sg13g2_decap_8 FILLER_8_676 ();
 sg13g2_decap_8 FILLER_8_683 ();
 sg13g2_decap_8 FILLER_8_690 ();
 sg13g2_decap_8 FILLER_8_697 ();
 sg13g2_decap_8 FILLER_8_704 ();
 sg13g2_decap_8 FILLER_8_711 ();
 sg13g2_decap_8 FILLER_8_718 ();
 sg13g2_decap_8 FILLER_8_725 ();
 sg13g2_decap_8 FILLER_8_732 ();
 sg13g2_decap_8 FILLER_8_739 ();
 sg13g2_decap_8 FILLER_8_746 ();
 sg13g2_decap_8 FILLER_8_753 ();
 sg13g2_decap_8 FILLER_8_760 ();
 sg13g2_decap_8 FILLER_8_767 ();
 sg13g2_decap_8 FILLER_8_774 ();
 sg13g2_decap_8 FILLER_8_781 ();
 sg13g2_decap_8 FILLER_8_788 ();
 sg13g2_decap_8 FILLER_8_795 ();
 sg13g2_decap_8 FILLER_8_802 ();
 sg13g2_decap_8 FILLER_8_809 ();
 sg13g2_decap_8 FILLER_8_816 ();
 sg13g2_decap_8 FILLER_8_823 ();
 sg13g2_decap_8 FILLER_8_830 ();
 sg13g2_decap_8 FILLER_8_837 ();
 sg13g2_decap_8 FILLER_8_844 ();
 sg13g2_decap_8 FILLER_8_851 ();
 sg13g2_decap_4 FILLER_8_858 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_fill_1 FILLER_9_188 ();
 sg13g2_fill_1 FILLER_9_222 ();
 sg13g2_fill_1 FILLER_9_250 ();
 sg13g2_fill_2 FILLER_9_299 ();
 sg13g2_fill_1 FILLER_9_301 ();
 sg13g2_fill_2 FILLER_9_334 ();
 sg13g2_fill_2 FILLER_9_438 ();
 sg13g2_fill_2 FILLER_9_504 ();
 sg13g2_fill_1 FILLER_9_506 ();
 sg13g2_fill_2 FILLER_9_539 ();
 sg13g2_decap_8 FILLER_9_572 ();
 sg13g2_fill_2 FILLER_9_579 ();
 sg13g2_decap_4 FILLER_9_588 ();
 sg13g2_fill_2 FILLER_9_592 ();
 sg13g2_decap_8 FILLER_9_602 ();
 sg13g2_decap_8 FILLER_9_609 ();
 sg13g2_decap_4 FILLER_9_616 ();
 sg13g2_fill_1 FILLER_9_620 ();
 sg13g2_decap_4 FILLER_9_649 ();
 sg13g2_fill_1 FILLER_9_653 ();
 sg13g2_decap_8 FILLER_9_674 ();
 sg13g2_fill_2 FILLER_9_681 ();
 sg13g2_decap_8 FILLER_9_688 ();
 sg13g2_fill_2 FILLER_9_695 ();
 sg13g2_decap_8 FILLER_9_710 ();
 sg13g2_decap_8 FILLER_9_717 ();
 sg13g2_decap_8 FILLER_9_724 ();
 sg13g2_decap_8 FILLER_9_731 ();
 sg13g2_decap_8 FILLER_9_738 ();
 sg13g2_decap_8 FILLER_9_745 ();
 sg13g2_decap_8 FILLER_9_752 ();
 sg13g2_decap_8 FILLER_9_759 ();
 sg13g2_decap_8 FILLER_9_766 ();
 sg13g2_decap_8 FILLER_9_773 ();
 sg13g2_decap_8 FILLER_9_780 ();
 sg13g2_decap_8 FILLER_9_787 ();
 sg13g2_decap_8 FILLER_9_794 ();
 sg13g2_decap_8 FILLER_9_801 ();
 sg13g2_decap_8 FILLER_9_808 ();
 sg13g2_decap_8 FILLER_9_815 ();
 sg13g2_decap_8 FILLER_9_822 ();
 sg13g2_decap_8 FILLER_9_829 ();
 sg13g2_decap_8 FILLER_9_836 ();
 sg13g2_decap_8 FILLER_9_843 ();
 sg13g2_decap_8 FILLER_9_850 ();
 sg13g2_decap_4 FILLER_9_857 ();
 sg13g2_fill_1 FILLER_9_861 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_fill_1 FILLER_10_188 ();
 sg13g2_fill_1 FILLER_10_257 ();
 sg13g2_fill_1 FILLER_10_276 ();
 sg13g2_fill_2 FILLER_10_336 ();
 sg13g2_fill_1 FILLER_10_347 ();
 sg13g2_fill_2 FILLER_10_430 ();
 sg13g2_fill_2 FILLER_10_476 ();
 sg13g2_fill_1 FILLER_10_478 ();
 sg13g2_fill_1 FILLER_10_493 ();
 sg13g2_fill_1 FILLER_10_552 ();
 sg13g2_fill_1 FILLER_10_562 ();
 sg13g2_fill_1 FILLER_10_579 ();
 sg13g2_fill_1 FILLER_10_617 ();
 sg13g2_decap_4 FILLER_10_623 ();
 sg13g2_fill_1 FILLER_10_645 ();
 sg13g2_fill_2 FILLER_10_658 ();
 sg13g2_fill_1 FILLER_10_668 ();
 sg13g2_fill_2 FILLER_10_685 ();
 sg13g2_decap_8 FILLER_10_711 ();
 sg13g2_decap_4 FILLER_10_718 ();
 sg13g2_decap_8 FILLER_10_730 ();
 sg13g2_decap_8 FILLER_10_737 ();
 sg13g2_decap_8 FILLER_10_744 ();
 sg13g2_decap_8 FILLER_10_751 ();
 sg13g2_decap_8 FILLER_10_758 ();
 sg13g2_decap_8 FILLER_10_765 ();
 sg13g2_decap_8 FILLER_10_772 ();
 sg13g2_decap_8 FILLER_10_779 ();
 sg13g2_decap_8 FILLER_10_786 ();
 sg13g2_decap_8 FILLER_10_793 ();
 sg13g2_decap_8 FILLER_10_800 ();
 sg13g2_decap_8 FILLER_10_807 ();
 sg13g2_decap_8 FILLER_10_814 ();
 sg13g2_decap_8 FILLER_10_821 ();
 sg13g2_decap_8 FILLER_10_828 ();
 sg13g2_decap_8 FILLER_10_835 ();
 sg13g2_decap_8 FILLER_10_842 ();
 sg13g2_decap_8 FILLER_10_849 ();
 sg13g2_decap_4 FILLER_10_856 ();
 sg13g2_fill_2 FILLER_10_860 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_63 ();
 sg13g2_decap_8 FILLER_11_70 ();
 sg13g2_fill_2 FILLER_11_188 ();
 sg13g2_fill_1 FILLER_11_190 ();
 sg13g2_fill_2 FILLER_11_256 ();
 sg13g2_fill_1 FILLER_11_356 ();
 sg13g2_fill_1 FILLER_11_468 ();
 sg13g2_fill_1 FILLER_11_478 ();
 sg13g2_fill_2 FILLER_11_519 ();
 sg13g2_fill_2 FILLER_11_556 ();
 sg13g2_fill_2 FILLER_11_563 ();
 sg13g2_decap_8 FILLER_11_569 ();
 sg13g2_decap_4 FILLER_11_576 ();
 sg13g2_fill_1 FILLER_11_580 ();
 sg13g2_decap_4 FILLER_11_586 ();
 sg13g2_fill_1 FILLER_11_590 ();
 sg13g2_fill_2 FILLER_11_605 ();
 sg13g2_decap_4 FILLER_11_631 ();
 sg13g2_decap_8 FILLER_11_645 ();
 sg13g2_decap_8 FILLER_11_652 ();
 sg13g2_decap_8 FILLER_11_673 ();
 sg13g2_decap_8 FILLER_11_680 ();
 sg13g2_decap_8 FILLER_11_687 ();
 sg13g2_fill_2 FILLER_11_694 ();
 sg13g2_fill_1 FILLER_11_696 ();
 sg13g2_decap_8 FILLER_11_702 ();
 sg13g2_fill_2 FILLER_11_709 ();
 sg13g2_decap_8 FILLER_11_736 ();
 sg13g2_decap_8 FILLER_11_743 ();
 sg13g2_fill_2 FILLER_11_750 ();
 sg13g2_decap_8 FILLER_11_756 ();
 sg13g2_decap_8 FILLER_11_763 ();
 sg13g2_fill_1 FILLER_11_770 ();
 sg13g2_decap_8 FILLER_11_784 ();
 sg13g2_decap_8 FILLER_11_791 ();
 sg13g2_decap_8 FILLER_11_798 ();
 sg13g2_decap_8 FILLER_11_805 ();
 sg13g2_decap_8 FILLER_11_812 ();
 sg13g2_decap_8 FILLER_11_819 ();
 sg13g2_decap_8 FILLER_11_826 ();
 sg13g2_decap_8 FILLER_11_833 ();
 sg13g2_decap_8 FILLER_11_840 ();
 sg13g2_decap_8 FILLER_11_847 ();
 sg13g2_decap_8 FILLER_11_854 ();
 sg13g2_fill_1 FILLER_11_861 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_decap_8 FILLER_12_56 ();
 sg13g2_decap_8 FILLER_12_63 ();
 sg13g2_decap_8 FILLER_12_70 ();
 sg13g2_fill_1 FILLER_12_224 ();
 sg13g2_fill_1 FILLER_12_296 ();
 sg13g2_fill_2 FILLER_12_395 ();
 sg13g2_fill_2 FILLER_12_403 ();
 sg13g2_fill_1 FILLER_12_405 ();
 sg13g2_fill_1 FILLER_12_490 ();
 sg13g2_fill_2 FILLER_12_541 ();
 sg13g2_fill_1 FILLER_12_561 ();
 sg13g2_decap_4 FILLER_12_586 ();
 sg13g2_fill_1 FILLER_12_602 ();
 sg13g2_fill_2 FILLER_12_615 ();
 sg13g2_decap_4 FILLER_12_621 ();
 sg13g2_fill_2 FILLER_12_625 ();
 sg13g2_fill_1 FILLER_12_675 ();
 sg13g2_decap_8 FILLER_12_710 ();
 sg13g2_decap_4 FILLER_12_717 ();
 sg13g2_fill_1 FILLER_12_721 ();
 sg13g2_decap_4 FILLER_12_732 ();
 sg13g2_fill_2 FILLER_12_736 ();
 sg13g2_fill_1 FILLER_12_792 ();
 sg13g2_decap_8 FILLER_12_805 ();
 sg13g2_decap_8 FILLER_12_812 ();
 sg13g2_decap_8 FILLER_12_819 ();
 sg13g2_decap_8 FILLER_12_826 ();
 sg13g2_decap_8 FILLER_12_833 ();
 sg13g2_decap_8 FILLER_12_840 ();
 sg13g2_decap_8 FILLER_12_847 ();
 sg13g2_decap_8 FILLER_12_854 ();
 sg13g2_fill_1 FILLER_12_861 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_decap_8 FILLER_13_49 ();
 sg13g2_decap_8 FILLER_13_56 ();
 sg13g2_decap_8 FILLER_13_63 ();
 sg13g2_decap_8 FILLER_13_70 ();
 sg13g2_fill_2 FILLER_13_188 ();
 sg13g2_fill_1 FILLER_13_190 ();
 sg13g2_fill_1 FILLER_13_267 ();
 sg13g2_fill_1 FILLER_13_300 ();
 sg13g2_fill_1 FILLER_13_323 ();
 sg13g2_fill_1 FILLER_13_383 ();
 sg13g2_fill_2 FILLER_13_412 ();
 sg13g2_fill_1 FILLER_13_414 ();
 sg13g2_fill_2 FILLER_13_428 ();
 sg13g2_fill_1 FILLER_13_536 ();
 sg13g2_decap_4 FILLER_13_557 ();
 sg13g2_fill_2 FILLER_13_579 ();
 sg13g2_fill_1 FILLER_13_581 ();
 sg13g2_fill_1 FILLER_13_603 ();
 sg13g2_fill_2 FILLER_13_609 ();
 sg13g2_fill_2 FILLER_13_619 ();
 sg13g2_fill_1 FILLER_13_621 ();
 sg13g2_fill_2 FILLER_13_629 ();
 sg13g2_fill_1 FILLER_13_647 ();
 sg13g2_fill_2 FILLER_13_673 ();
 sg13g2_decap_8 FILLER_13_687 ();
 sg13g2_fill_1 FILLER_13_717 ();
 sg13g2_fill_2 FILLER_13_723 ();
 sg13g2_fill_2 FILLER_13_741 ();
 sg13g2_fill_2 FILLER_13_748 ();
 sg13g2_fill_1 FILLER_13_750 ();
 sg13g2_decap_8 FILLER_13_760 ();
 sg13g2_fill_2 FILLER_13_767 ();
 sg13g2_fill_1 FILLER_13_769 ();
 sg13g2_decap_8 FILLER_13_790 ();
 sg13g2_decap_8 FILLER_13_810 ();
 sg13g2_decap_8 FILLER_13_817 ();
 sg13g2_decap_8 FILLER_13_824 ();
 sg13g2_decap_8 FILLER_13_831 ();
 sg13g2_decap_8 FILLER_13_838 ();
 sg13g2_decap_8 FILLER_13_845 ();
 sg13g2_decap_8 FILLER_13_852 ();
 sg13g2_fill_2 FILLER_13_859 ();
 sg13g2_fill_1 FILLER_13_861 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_decap_8 FILLER_14_42 ();
 sg13g2_decap_8 FILLER_14_49 ();
 sg13g2_decap_8 FILLER_14_56 ();
 sg13g2_decap_8 FILLER_14_63 ();
 sg13g2_decap_8 FILLER_14_70 ();
 sg13g2_fill_1 FILLER_14_233 ();
 sg13g2_fill_2 FILLER_14_283 ();
 sg13g2_fill_1 FILLER_14_285 ();
 sg13g2_fill_2 FILLER_14_352 ();
 sg13g2_fill_2 FILLER_14_404 ();
 sg13g2_fill_1 FILLER_14_434 ();
 sg13g2_fill_2 FILLER_14_475 ();
 sg13g2_decap_4 FILLER_14_575 ();
 sg13g2_fill_2 FILLER_14_579 ();
 sg13g2_fill_2 FILLER_14_598 ();
 sg13g2_fill_1 FILLER_14_600 ();
 sg13g2_decap_4 FILLER_14_617 ();
 sg13g2_decap_4 FILLER_14_650 ();
 sg13g2_fill_1 FILLER_14_654 ();
 sg13g2_fill_2 FILLER_14_709 ();
 sg13g2_fill_1 FILLER_14_727 ();
 sg13g2_fill_2 FILLER_14_732 ();
 sg13g2_fill_1 FILLER_14_734 ();
 sg13g2_fill_1 FILLER_14_764 ();
 sg13g2_fill_2 FILLER_14_789 ();
 sg13g2_decap_4 FILLER_14_814 ();
 sg13g2_fill_2 FILLER_14_818 ();
 sg13g2_decap_8 FILLER_14_832 ();
 sg13g2_decap_8 FILLER_14_839 ();
 sg13g2_decap_8 FILLER_14_846 ();
 sg13g2_decap_8 FILLER_14_853 ();
 sg13g2_fill_2 FILLER_14_860 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_8 FILLER_15_35 ();
 sg13g2_decap_8 FILLER_15_42 ();
 sg13g2_decap_8 FILLER_15_49 ();
 sg13g2_decap_8 FILLER_15_56 ();
 sg13g2_decap_8 FILLER_15_63 ();
 sg13g2_decap_8 FILLER_15_70 ();
 sg13g2_fill_2 FILLER_15_223 ();
 sg13g2_fill_1 FILLER_15_331 ();
 sg13g2_fill_1 FILLER_15_530 ();
 sg13g2_fill_1 FILLER_15_561 ();
 sg13g2_fill_2 FILLER_15_575 ();
 sg13g2_fill_1 FILLER_15_598 ();
 sg13g2_decap_8 FILLER_15_650 ();
 sg13g2_decap_8 FILLER_15_657 ();
 sg13g2_fill_2 FILLER_15_664 ();
 sg13g2_decap_8 FILLER_15_673 ();
 sg13g2_decap_4 FILLER_15_680 ();
 sg13g2_fill_1 FILLER_15_684 ();
 sg13g2_decap_4 FILLER_15_700 ();
 sg13g2_fill_2 FILLER_15_704 ();
 sg13g2_fill_2 FILLER_15_729 ();
 sg13g2_fill_1 FILLER_15_731 ();
 sg13g2_fill_1 FILLER_15_736 ();
 sg13g2_decap_8 FILLER_15_742 ();
 sg13g2_fill_2 FILLER_15_749 ();
 sg13g2_decap_4 FILLER_15_763 ();
 sg13g2_fill_1 FILLER_15_767 ();
 sg13g2_decap_4 FILLER_15_795 ();
 sg13g2_fill_1 FILLER_15_799 ();
 sg13g2_decap_4 FILLER_15_812 ();
 sg13g2_decap_8 FILLER_15_837 ();
 sg13g2_decap_8 FILLER_15_844 ();
 sg13g2_decap_8 FILLER_15_851 ();
 sg13g2_decap_4 FILLER_15_858 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_decap_8 FILLER_16_35 ();
 sg13g2_decap_8 FILLER_16_42 ();
 sg13g2_decap_8 FILLER_16_49 ();
 sg13g2_decap_8 FILLER_16_56 ();
 sg13g2_decap_8 FILLER_16_63 ();
 sg13g2_decap_8 FILLER_16_70 ();
 sg13g2_fill_1 FILLER_16_209 ();
 sg13g2_fill_1 FILLER_16_238 ();
 sg13g2_fill_1 FILLER_16_248 ();
 sg13g2_fill_1 FILLER_16_262 ();
 sg13g2_fill_1 FILLER_16_361 ();
 sg13g2_fill_1 FILLER_16_384 ();
 sg13g2_fill_2 FILLER_16_415 ();
 sg13g2_fill_1 FILLER_16_417 ();
 sg13g2_fill_2 FILLER_16_530 ();
 sg13g2_fill_1 FILLER_16_532 ();
 sg13g2_decap_4 FILLER_16_553 ();
 sg13g2_fill_2 FILLER_16_565 ();
 sg13g2_fill_1 FILLER_16_580 ();
 sg13g2_fill_1 FILLER_16_598 ();
 sg13g2_decap_8 FILLER_16_615 ();
 sg13g2_decap_8 FILLER_16_622 ();
 sg13g2_fill_1 FILLER_16_629 ();
 sg13g2_fill_1 FILLER_16_640 ();
 sg13g2_decap_4 FILLER_16_657 ();
 sg13g2_fill_1 FILLER_16_661 ();
 sg13g2_fill_2 FILLER_16_683 ();
 sg13g2_fill_2 FILLER_16_701 ();
 sg13g2_fill_1 FILLER_16_703 ();
 sg13g2_fill_2 FILLER_16_746 ();
 sg13g2_fill_1 FILLER_16_748 ();
 sg13g2_decap_8 FILLER_16_754 ();
 sg13g2_decap_8 FILLER_16_761 ();
 sg13g2_fill_2 FILLER_16_768 ();
 sg13g2_decap_8 FILLER_16_788 ();
 sg13g2_fill_1 FILLER_16_795 ();
 sg13g2_fill_1 FILLER_16_825 ();
 sg13g2_decap_8 FILLER_16_831 ();
 sg13g2_decap_8 FILLER_16_838 ();
 sg13g2_decap_8 FILLER_16_845 ();
 sg13g2_decap_8 FILLER_16_852 ();
 sg13g2_fill_2 FILLER_16_859 ();
 sg13g2_fill_1 FILLER_16_861 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_28 ();
 sg13g2_decap_8 FILLER_17_35 ();
 sg13g2_decap_8 FILLER_17_42 ();
 sg13g2_decap_8 FILLER_17_49 ();
 sg13g2_decap_8 FILLER_17_56 ();
 sg13g2_decap_8 FILLER_17_63 ();
 sg13g2_decap_8 FILLER_17_70 ();
 sg13g2_fill_1 FILLER_17_201 ();
 sg13g2_fill_2 FILLER_17_232 ();
 sg13g2_fill_1 FILLER_17_289 ();
 sg13g2_fill_2 FILLER_17_303 ();
 sg13g2_fill_1 FILLER_17_305 ();
 sg13g2_fill_1 FILLER_17_335 ();
 sg13g2_fill_1 FILLER_17_483 ();
 sg13g2_fill_2 FILLER_17_521 ();
 sg13g2_fill_1 FILLER_17_528 ();
 sg13g2_decap_4 FILLER_17_545 ();
 sg13g2_fill_1 FILLER_17_549 ();
 sg13g2_fill_2 FILLER_17_560 ();
 sg13g2_fill_1 FILLER_17_562 ();
 sg13g2_fill_2 FILLER_17_566 ();
 sg13g2_decap_8 FILLER_17_584 ();
 sg13g2_decap_4 FILLER_17_591 ();
 sg13g2_fill_2 FILLER_17_595 ();
 sg13g2_decap_8 FILLER_17_612 ();
 sg13g2_decap_4 FILLER_17_619 ();
 sg13g2_fill_2 FILLER_17_623 ();
 sg13g2_fill_2 FILLER_17_657 ();
 sg13g2_fill_1 FILLER_17_669 ();
 sg13g2_fill_2 FILLER_17_687 ();
 sg13g2_fill_1 FILLER_17_689 ();
 sg13g2_decap_4 FILLER_17_693 ();
 sg13g2_decap_4 FILLER_17_706 ();
 sg13g2_fill_1 FILLER_17_722 ();
 sg13g2_fill_1 FILLER_17_726 ();
 sg13g2_decap_8 FILLER_17_731 ();
 sg13g2_decap_4 FILLER_17_738 ();
 sg13g2_decap_4 FILLER_17_757 ();
 sg13g2_fill_1 FILLER_17_761 ();
 sg13g2_fill_1 FILLER_17_770 ();
 sg13g2_fill_2 FILLER_17_779 ();
 sg13g2_decap_4 FILLER_17_793 ();
 sg13g2_fill_1 FILLER_17_814 ();
 sg13g2_decap_8 FILLER_17_837 ();
 sg13g2_fill_2 FILLER_17_844 ();
 sg13g2_fill_1 FILLER_17_846 ();
 sg13g2_decap_8 FILLER_17_852 ();
 sg13g2_fill_2 FILLER_17_859 ();
 sg13g2_fill_1 FILLER_17_861 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_21 ();
 sg13g2_decap_8 FILLER_18_28 ();
 sg13g2_decap_8 FILLER_18_35 ();
 sg13g2_decap_8 FILLER_18_42 ();
 sg13g2_decap_8 FILLER_18_49 ();
 sg13g2_decap_8 FILLER_18_56 ();
 sg13g2_decap_8 FILLER_18_63 ();
 sg13g2_decap_4 FILLER_18_70 ();
 sg13g2_fill_2 FILLER_18_74 ();
 sg13g2_fill_2 FILLER_18_130 ();
 sg13g2_fill_1 FILLER_18_147 ();
 sg13g2_fill_2 FILLER_18_175 ();
 sg13g2_fill_1 FILLER_18_247 ();
 sg13g2_fill_2 FILLER_18_283 ();
 sg13g2_fill_1 FILLER_18_374 ();
 sg13g2_fill_2 FILLER_18_417 ();
 sg13g2_fill_1 FILLER_18_419 ();
 sg13g2_fill_1 FILLER_18_426 ();
 sg13g2_fill_2 FILLER_18_446 ();
 sg13g2_fill_2 FILLER_18_470 ();
 sg13g2_fill_1 FILLER_18_522 ();
 sg13g2_decap_8 FILLER_18_541 ();
 sg13g2_decap_4 FILLER_18_548 ();
 sg13g2_decap_4 FILLER_18_565 ();
 sg13g2_fill_1 FILLER_18_574 ();
 sg13g2_decap_4 FILLER_18_591 ();
 sg13g2_fill_1 FILLER_18_595 ();
 sg13g2_fill_1 FILLER_18_610 ();
 sg13g2_decap_8 FILLER_18_647 ();
 sg13g2_decap_4 FILLER_18_654 ();
 sg13g2_fill_1 FILLER_18_658 ();
 sg13g2_decap_4 FILLER_18_663 ();
 sg13g2_fill_2 FILLER_18_667 ();
 sg13g2_decap_8 FILLER_18_682 ();
 sg13g2_fill_2 FILLER_18_689 ();
 sg13g2_decap_4 FILLER_18_712 ();
 sg13g2_fill_2 FILLER_18_716 ();
 sg13g2_fill_2 FILLER_18_739 ();
 sg13g2_fill_1 FILLER_18_741 ();
 sg13g2_fill_1 FILLER_18_756 ();
 sg13g2_decap_8 FILLER_18_760 ();
 sg13g2_fill_1 FILLER_18_767 ();
 sg13g2_fill_2 FILLER_18_772 ();
 sg13g2_fill_2 FILLER_18_791 ();
 sg13g2_fill_1 FILLER_18_793 ();
 sg13g2_decap_4 FILLER_18_806 ();
 sg13g2_decap_4 FILLER_18_815 ();
 sg13g2_decap_8 FILLER_18_855 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_decap_8 FILLER_19_28 ();
 sg13g2_decap_8 FILLER_19_35 ();
 sg13g2_decap_4 FILLER_19_42 ();
 sg13g2_fill_2 FILLER_19_46 ();
 sg13g2_decap_8 FILLER_19_52 ();
 sg13g2_decap_8 FILLER_19_59 ();
 sg13g2_decap_8 FILLER_19_66 ();
 sg13g2_fill_1 FILLER_19_73 ();
 sg13g2_fill_1 FILLER_19_154 ();
 sg13g2_fill_1 FILLER_19_205 ();
 sg13g2_fill_2 FILLER_19_244 ();
 sg13g2_fill_1 FILLER_19_291 ();
 sg13g2_fill_2 FILLER_19_305 ();
 sg13g2_fill_2 FILLER_19_325 ();
 sg13g2_fill_1 FILLER_19_332 ();
 sg13g2_fill_1 FILLER_19_346 ();
 sg13g2_fill_1 FILLER_19_383 ();
 sg13g2_fill_1 FILLER_19_403 ();
 sg13g2_fill_1 FILLER_19_454 ();
 sg13g2_fill_2 FILLER_19_482 ();
 sg13g2_fill_1 FILLER_19_484 ();
 sg13g2_fill_2 FILLER_19_505 ();
 sg13g2_fill_1 FILLER_19_507 ();
 sg13g2_fill_2 FILLER_19_524 ();
 sg13g2_fill_1 FILLER_19_534 ();
 sg13g2_fill_2 FILLER_19_556 ();
 sg13g2_fill_1 FILLER_19_571 ();
 sg13g2_fill_2 FILLER_19_601 ();
 sg13g2_decap_8 FILLER_19_616 ();
 sg13g2_fill_1 FILLER_19_623 ();
 sg13g2_fill_2 FILLER_19_636 ();
 sg13g2_fill_2 FILLER_19_659 ();
 sg13g2_fill_1 FILLER_19_665 ();
 sg13g2_decap_8 FILLER_19_681 ();
 sg13g2_decap_4 FILLER_19_688 ();
 sg13g2_fill_2 FILLER_19_692 ();
 sg13g2_decap_8 FILLER_19_707 ();
 sg13g2_decap_4 FILLER_19_714 ();
 sg13g2_fill_1 FILLER_19_718 ();
 sg13g2_fill_1 FILLER_19_758 ();
 sg13g2_decap_4 FILLER_19_785 ();
 sg13g2_fill_1 FILLER_19_789 ();
 sg13g2_decap_8 FILLER_19_794 ();
 sg13g2_decap_4 FILLER_19_819 ();
 sg13g2_fill_2 FILLER_19_841 ();
 sg13g2_fill_1 FILLER_19_843 ();
 sg13g2_decap_4 FILLER_19_856 ();
 sg13g2_fill_2 FILLER_19_860 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_fill_2 FILLER_20_14 ();
 sg13g2_fill_2 FILLER_20_82 ();
 sg13g2_fill_1 FILLER_20_84 ();
 sg13g2_fill_1 FILLER_20_146 ();
 sg13g2_fill_2 FILLER_20_169 ();
 sg13g2_fill_1 FILLER_20_171 ();
 sg13g2_fill_2 FILLER_20_191 ();
 sg13g2_fill_1 FILLER_20_193 ();
 sg13g2_fill_1 FILLER_20_217 ();
 sg13g2_fill_2 FILLER_20_355 ();
 sg13g2_fill_1 FILLER_20_357 ();
 sg13g2_fill_2 FILLER_20_437 ();
 sg13g2_fill_2 FILLER_20_479 ();
 sg13g2_decap_4 FILLER_20_498 ();
 sg13g2_fill_1 FILLER_20_502 ();
 sg13g2_fill_1 FILLER_20_519 ();
 sg13g2_fill_1 FILLER_20_525 ();
 sg13g2_fill_2 FILLER_20_537 ();
 sg13g2_decap_4 FILLER_20_560 ();
 sg13g2_decap_4 FILLER_20_567 ();
 sg13g2_fill_1 FILLER_20_571 ();
 sg13g2_decap_8 FILLER_20_587 ();
 sg13g2_fill_1 FILLER_20_594 ();
 sg13g2_fill_2 FILLER_20_617 ();
 sg13g2_fill_1 FILLER_20_627 ();
 sg13g2_fill_1 FILLER_20_642 ();
 sg13g2_fill_2 FILLER_20_648 ();
 sg13g2_fill_1 FILLER_20_650 ();
 sg13g2_fill_1 FILLER_20_659 ();
 sg13g2_decap_4 FILLER_20_681 ();
 sg13g2_fill_1 FILLER_20_685 ();
 sg13g2_fill_1 FILLER_20_694 ();
 sg13g2_fill_2 FILLER_20_731 ();
 sg13g2_fill_1 FILLER_20_733 ();
 sg13g2_fill_2 FILLER_20_747 ();
 sg13g2_fill_2 FILLER_20_766 ();
 sg13g2_fill_1 FILLER_20_768 ();
 sg13g2_fill_2 FILLER_20_781 ();
 sg13g2_fill_2 FILLER_20_804 ();
 sg13g2_fill_2 FILLER_20_820 ();
 sg13g2_fill_1 FILLER_20_822 ();
 sg13g2_fill_2 FILLER_20_843 ();
 sg13g2_fill_1 FILLER_20_845 ();
 sg13g2_decap_8 FILLER_20_854 ();
 sg13g2_fill_1 FILLER_20_861 ();
 sg13g2_fill_1 FILLER_21_0 ();
 sg13g2_fill_2 FILLER_21_9 ();
 sg13g2_decap_8 FILLER_21_15 ();
 sg13g2_fill_2 FILLER_21_22 ();
 sg13g2_fill_1 FILLER_21_24 ();
 sg13g2_decap_8 FILLER_21_56 ();
 sg13g2_fill_2 FILLER_21_63 ();
 sg13g2_fill_1 FILLER_21_244 ();
 sg13g2_fill_2 FILLER_21_281 ();
 sg13g2_fill_1 FILLER_21_296 ();
 sg13g2_fill_2 FILLER_21_327 ();
 sg13g2_fill_2 FILLER_21_351 ();
 sg13g2_fill_1 FILLER_21_353 ();
 sg13g2_fill_2 FILLER_21_434 ();
 sg13g2_fill_2 FILLER_21_452 ();
 sg13g2_fill_2 FILLER_21_482 ();
 sg13g2_fill_1 FILLER_21_505 ();
 sg13g2_decap_4 FILLER_21_530 ();
 sg13g2_fill_1 FILLER_21_534 ();
 sg13g2_decap_8 FILLER_21_566 ();
 sg13g2_fill_1 FILLER_21_573 ();
 sg13g2_decap_4 FILLER_21_587 ();
 sg13g2_decap_8 FILLER_21_609 ();
 sg13g2_fill_2 FILLER_21_616 ();
 sg13g2_fill_1 FILLER_21_618 ();
 sg13g2_decap_8 FILLER_21_628 ();
 sg13g2_decap_4 FILLER_21_635 ();
 sg13g2_fill_2 FILLER_21_639 ();
 sg13g2_fill_2 FILLER_21_645 ();
 sg13g2_fill_1 FILLER_21_647 ();
 sg13g2_decap_4 FILLER_21_664 ();
 sg13g2_fill_2 FILLER_21_668 ();
 sg13g2_fill_2 FILLER_21_674 ();
 sg13g2_fill_1 FILLER_21_676 ();
 sg13g2_decap_4 FILLER_21_715 ();
 sg13g2_fill_1 FILLER_21_719 ();
 sg13g2_decap_4 FILLER_21_724 ();
 sg13g2_fill_1 FILLER_21_728 ();
 sg13g2_decap_8 FILLER_21_754 ();
 sg13g2_decap_4 FILLER_21_761 ();
 sg13g2_decap_8 FILLER_21_788 ();
 sg13g2_decap_8 FILLER_21_795 ();
 sg13g2_fill_2 FILLER_21_826 ();
 sg13g2_fill_1 FILLER_21_828 ();
 sg13g2_fill_1 FILLER_21_842 ();
 sg13g2_fill_2 FILLER_21_860 ();
 sg13g2_fill_1 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_32 ();
 sg13g2_fill_2 FILLER_22_39 ();
 sg13g2_fill_1 FILLER_22_68 ();
 sg13g2_fill_2 FILLER_22_117 ();
 sg13g2_fill_2 FILLER_22_158 ();
 sg13g2_fill_1 FILLER_22_160 ();
 sg13g2_fill_2 FILLER_22_180 ();
 sg13g2_fill_1 FILLER_22_182 ();
 sg13g2_fill_1 FILLER_22_201 ();
 sg13g2_fill_1 FILLER_22_239 ();
 sg13g2_fill_1 FILLER_22_270 ();
 sg13g2_fill_2 FILLER_22_280 ();
 sg13g2_fill_2 FILLER_22_295 ();
 sg13g2_fill_1 FILLER_22_297 ();
 sg13g2_fill_2 FILLER_22_343 ();
 sg13g2_fill_1 FILLER_22_345 ();
 sg13g2_fill_1 FILLER_22_413 ();
 sg13g2_decap_4 FILLER_22_446 ();
 sg13g2_fill_2 FILLER_22_450 ();
 sg13g2_fill_1 FILLER_22_460 ();
 sg13g2_decap_4 FILLER_22_474 ();
 sg13g2_fill_1 FILLER_22_478 ();
 sg13g2_fill_1 FILLER_22_487 ();
 sg13g2_decap_4 FILLER_22_509 ();
 sg13g2_decap_8 FILLER_22_529 ();
 sg13g2_fill_2 FILLER_22_536 ();
 sg13g2_fill_1 FILLER_22_538 ();
 sg13g2_decap_4 FILLER_22_559 ();
 sg13g2_fill_2 FILLER_22_615 ();
 sg13g2_decap_4 FILLER_22_667 ();
 sg13g2_fill_1 FILLER_22_671 ();
 sg13g2_fill_2 FILLER_22_710 ();
 sg13g2_decap_4 FILLER_22_725 ();
 sg13g2_fill_2 FILLER_22_737 ();
 sg13g2_fill_1 FILLER_22_739 ();
 sg13g2_decap_4 FILLER_22_756 ();
 sg13g2_decap_4 FILLER_22_768 ();
 sg13g2_fill_2 FILLER_22_772 ();
 sg13g2_decap_4 FILLER_22_792 ();
 sg13g2_fill_2 FILLER_22_806 ();
 sg13g2_fill_1 FILLER_22_808 ();
 sg13g2_fill_1 FILLER_22_814 ();
 sg13g2_fill_2 FILLER_22_820 ();
 sg13g2_decap_4 FILLER_22_834 ();
 sg13g2_fill_2 FILLER_22_846 ();
 sg13g2_fill_1 FILLER_22_848 ();
 sg13g2_decap_8 FILLER_22_854 ();
 sg13g2_fill_1 FILLER_22_861 ();
 sg13g2_decap_4 FILLER_23_39 ();
 sg13g2_decap_8 FILLER_23_51 ();
 sg13g2_decap_4 FILLER_23_58 ();
 sg13g2_fill_1 FILLER_23_62 ();
 sg13g2_fill_2 FILLER_23_126 ();
 sg13g2_fill_2 FILLER_23_180 ();
 sg13g2_fill_2 FILLER_23_224 ();
 sg13g2_fill_2 FILLER_23_238 ();
 sg13g2_fill_2 FILLER_23_256 ();
 sg13g2_fill_2 FILLER_23_296 ();
 sg13g2_fill_2 FILLER_23_304 ();
 sg13g2_fill_2 FILLER_23_322 ();
 sg13g2_fill_1 FILLER_23_364 ();
 sg13g2_fill_1 FILLER_23_373 ();
 sg13g2_fill_2 FILLER_23_383 ();
 sg13g2_fill_1 FILLER_23_385 ();
 sg13g2_fill_2 FILLER_23_418 ();
 sg13g2_fill_1 FILLER_23_420 ();
 sg13g2_fill_1 FILLER_23_449 ();
 sg13g2_decap_4 FILLER_23_484 ();
 sg13g2_fill_2 FILLER_23_511 ();
 sg13g2_fill_1 FILLER_23_513 ();
 sg13g2_fill_1 FILLER_23_535 ();
 sg13g2_fill_2 FILLER_23_557 ();
 sg13g2_fill_1 FILLER_23_559 ();
 sg13g2_fill_1 FILLER_23_591 ();
 sg13g2_fill_2 FILLER_23_627 ();
 sg13g2_fill_1 FILLER_23_629 ();
 sg13g2_fill_2 FILLER_23_643 ();
 sg13g2_fill_1 FILLER_23_645 ();
 sg13g2_fill_2 FILLER_23_653 ();
 sg13g2_fill_1 FILLER_23_675 ();
 sg13g2_fill_2 FILLER_23_684 ();
 sg13g2_decap_4 FILLER_23_716 ();
 sg13g2_decap_8 FILLER_23_724 ();
 sg13g2_fill_1 FILLER_23_731 ();
 sg13g2_decap_4 FILLER_23_737 ();
 sg13g2_decap_8 FILLER_23_770 ();
 sg13g2_fill_1 FILLER_23_777 ();
 sg13g2_decap_8 FILLER_23_791 ();
 sg13g2_fill_1 FILLER_23_806 ();
 sg13g2_fill_1 FILLER_23_815 ();
 sg13g2_decap_8 FILLER_23_827 ();
 sg13g2_decap_4 FILLER_23_857 ();
 sg13g2_fill_1 FILLER_23_861 ();
 sg13g2_fill_2 FILLER_24_14 ();
 sg13g2_fill_2 FILLER_24_36 ();
 sg13g2_fill_2 FILLER_24_43 ();
 sg13g2_fill_1 FILLER_24_45 ();
 sg13g2_fill_2 FILLER_24_94 ();
 sg13g2_fill_1 FILLER_24_132 ();
 sg13g2_fill_1 FILLER_24_181 ();
 sg13g2_fill_1 FILLER_24_334 ();
 sg13g2_fill_2 FILLER_24_350 ();
 sg13g2_fill_1 FILLER_24_397 ();
 sg13g2_fill_2 FILLER_24_404 ();
 sg13g2_fill_1 FILLER_24_411 ();
 sg13g2_decap_8 FILLER_24_444 ();
 sg13g2_fill_2 FILLER_24_451 ();
 sg13g2_fill_1 FILLER_24_474 ();
 sg13g2_decap_4 FILLER_24_480 ();
 sg13g2_fill_1 FILLER_24_488 ();
 sg13g2_decap_8 FILLER_24_503 ();
 sg13g2_fill_1 FILLER_24_510 ();
 sg13g2_decap_8 FILLER_24_529 ();
 sg13g2_fill_2 FILLER_24_536 ();
 sg13g2_fill_2 FILLER_24_563 ();
 sg13g2_fill_1 FILLER_24_565 ();
 sg13g2_fill_1 FILLER_24_571 ();
 sg13g2_decap_8 FILLER_24_586 ();
 sg13g2_fill_2 FILLER_24_593 ();
 sg13g2_fill_1 FILLER_24_595 ();
 sg13g2_decap_4 FILLER_24_617 ();
 sg13g2_fill_2 FILLER_24_621 ();
 sg13g2_fill_1 FILLER_24_626 ();
 sg13g2_fill_1 FILLER_24_657 ();
 sg13g2_decap_4 FILLER_24_662 ();
 sg13g2_fill_1 FILLER_24_666 ();
 sg13g2_fill_1 FILLER_24_689 ();
 sg13g2_decap_8 FILLER_24_706 ();
 sg13g2_fill_2 FILLER_24_713 ();
 sg13g2_fill_1 FILLER_24_715 ();
 sg13g2_decap_8 FILLER_24_732 ();
 sg13g2_decap_8 FILLER_24_739 ();
 sg13g2_fill_1 FILLER_24_746 ();
 sg13g2_fill_2 FILLER_24_752 ();
 sg13g2_fill_1 FILLER_24_754 ();
 sg13g2_fill_2 FILLER_24_760 ();
 sg13g2_fill_1 FILLER_24_762 ();
 sg13g2_fill_2 FILLER_24_795 ();
 sg13g2_fill_1 FILLER_24_797 ();
 sg13g2_decap_8 FILLER_24_806 ();
 sg13g2_decap_8 FILLER_24_813 ();
 sg13g2_decap_4 FILLER_24_820 ();
 sg13g2_fill_1 FILLER_24_836 ();
 sg13g2_fill_2 FILLER_25_12 ();
 sg13g2_fill_2 FILLER_25_50 ();
 sg13g2_fill_1 FILLER_25_52 ();
 sg13g2_fill_1 FILLER_25_80 ();
 sg13g2_fill_2 FILLER_25_224 ();
 sg13g2_fill_2 FILLER_25_249 ();
 sg13g2_fill_1 FILLER_25_379 ();
 sg13g2_decap_4 FILLER_25_440 ();
 sg13g2_fill_1 FILLER_25_444 ();
 sg13g2_decap_4 FILLER_25_469 ();
 sg13g2_fill_2 FILLER_25_493 ();
 sg13g2_fill_2 FILLER_25_499 ();
 sg13g2_fill_2 FILLER_25_510 ();
 sg13g2_fill_2 FILLER_25_527 ();
 sg13g2_fill_1 FILLER_25_529 ();
 sg13g2_fill_2 FILLER_25_533 ();
 sg13g2_decap_4 FILLER_25_543 ();
 sg13g2_fill_1 FILLER_25_556 ();
 sg13g2_fill_2 FILLER_25_565 ();
 sg13g2_fill_1 FILLER_25_567 ();
 sg13g2_decap_4 FILLER_25_580 ();
 sg13g2_fill_1 FILLER_25_584 ();
 sg13g2_fill_2 FILLER_25_604 ();
 sg13g2_fill_1 FILLER_25_606 ();
 sg13g2_fill_2 FILLER_25_616 ();
 sg13g2_fill_1 FILLER_25_631 ();
 sg13g2_decap_4 FILLER_25_657 ();
 sg13g2_fill_2 FILLER_25_661 ();
 sg13g2_fill_1 FILLER_25_671 ();
 sg13g2_fill_1 FILLER_25_684 ();
 sg13g2_fill_2 FILLER_25_698 ();
 sg13g2_fill_1 FILLER_25_700 ();
 sg13g2_fill_1 FILLER_25_721 ();
 sg13g2_fill_2 FILLER_25_735 ();
 sg13g2_fill_2 FILLER_25_763 ();
 sg13g2_fill_2 FILLER_25_773 ();
 sg13g2_decap_4 FILLER_25_789 ();
 sg13g2_fill_2 FILLER_25_813 ();
 sg13g2_fill_2 FILLER_25_840 ();
 sg13g2_fill_1 FILLER_25_842 ();
 sg13g2_fill_2 FILLER_25_860 ();
 sg13g2_fill_1 FILLER_26_0 ();
 sg13g2_fill_2 FILLER_26_9 ();
 sg13g2_fill_1 FILLER_26_49 ();
 sg13g2_fill_2 FILLER_26_103 ();
 sg13g2_fill_1 FILLER_26_105 ();
 sg13g2_fill_2 FILLER_26_152 ();
 sg13g2_fill_1 FILLER_26_164 ();
 sg13g2_fill_1 FILLER_26_171 ();
 sg13g2_fill_2 FILLER_26_181 ();
 sg13g2_fill_2 FILLER_26_285 ();
 sg13g2_fill_2 FILLER_26_301 ();
 sg13g2_fill_1 FILLER_26_303 ();
 sg13g2_fill_2 FILLER_26_311 ();
 sg13g2_fill_1 FILLER_26_313 ();
 sg13g2_fill_2 FILLER_26_339 ();
 sg13g2_fill_2 FILLER_26_353 ();
 sg13g2_fill_1 FILLER_26_407 ();
 sg13g2_fill_2 FILLER_26_441 ();
 sg13g2_fill_1 FILLER_26_443 ();
 sg13g2_fill_2 FILLER_26_458 ();
 sg13g2_fill_2 FILLER_26_482 ();
 sg13g2_fill_1 FILLER_26_484 ();
 sg13g2_fill_2 FILLER_26_510 ();
 sg13g2_fill_1 FILLER_26_518 ();
 sg13g2_decap_8 FILLER_26_523 ();
 sg13g2_fill_2 FILLER_26_547 ();
 sg13g2_decap_8 FILLER_26_652 ();
 sg13g2_fill_2 FILLER_26_659 ();
 sg13g2_fill_2 FILLER_26_674 ();
 sg13g2_fill_1 FILLER_26_689 ();
 sg13g2_decap_8 FILLER_26_695 ();
 sg13g2_decap_8 FILLER_26_702 ();
 sg13g2_fill_2 FILLER_26_709 ();
 sg13g2_fill_1 FILLER_26_711 ();
 sg13g2_fill_2 FILLER_26_729 ();
 sg13g2_decap_4 FILLER_26_756 ();
 sg13g2_fill_2 FILLER_26_760 ();
 sg13g2_fill_2 FILLER_26_769 ();
 sg13g2_decap_8 FILLER_26_801 ();
 sg13g2_decap_4 FILLER_26_808 ();
 sg13g2_decap_8 FILLER_26_829 ();
 sg13g2_decap_4 FILLER_26_836 ();
 sg13g2_fill_2 FILLER_26_845 ();
 sg13g2_fill_1 FILLER_26_847 ();
 sg13g2_fill_1 FILLER_26_861 ();
 sg13g2_fill_1 FILLER_27_0 ();
 sg13g2_fill_1 FILLER_27_29 ();
 sg13g2_fill_1 FILLER_27_52 ();
 sg13g2_fill_1 FILLER_27_80 ();
 sg13g2_fill_2 FILLER_27_110 ();
 sg13g2_fill_1 FILLER_27_112 ();
 sg13g2_fill_1 FILLER_27_131 ();
 sg13g2_fill_1 FILLER_27_177 ();
 sg13g2_fill_1 FILLER_27_297 ();
 sg13g2_fill_1 FILLER_27_326 ();
 sg13g2_fill_1 FILLER_27_335 ();
 sg13g2_fill_1 FILLER_27_385 ();
 sg13g2_fill_2 FILLER_27_391 ();
 sg13g2_fill_1 FILLER_27_400 ();
 sg13g2_fill_2 FILLER_27_409 ();
 sg13g2_fill_1 FILLER_27_411 ();
 sg13g2_fill_2 FILLER_27_430 ();
 sg13g2_fill_1 FILLER_27_432 ();
 sg13g2_fill_2 FILLER_27_490 ();
 sg13g2_fill_1 FILLER_27_492 ();
 sg13g2_fill_1 FILLER_27_506 ();
 sg13g2_decap_4 FILLER_27_515 ();
 sg13g2_decap_8 FILLER_27_544 ();
 sg13g2_fill_1 FILLER_27_551 ();
 sg13g2_fill_2 FILLER_27_569 ();
 sg13g2_decap_8 FILLER_27_575 ();
 sg13g2_fill_2 FILLER_27_582 ();
 sg13g2_fill_1 FILLER_27_584 ();
 sg13g2_fill_2 FILLER_27_607 ();
 sg13g2_fill_1 FILLER_27_609 ();
 sg13g2_fill_1 FILLER_27_614 ();
 sg13g2_fill_2 FILLER_27_623 ();
 sg13g2_decap_4 FILLER_27_639 ();
 sg13g2_fill_2 FILLER_27_643 ();
 sg13g2_decap_8 FILLER_27_658 ();
 sg13g2_fill_2 FILLER_27_682 ();
 sg13g2_decap_8 FILLER_27_689 ();
 sg13g2_fill_1 FILLER_27_696 ();
 sg13g2_fill_2 FILLER_27_717 ();
 sg13g2_fill_1 FILLER_27_728 ();
 sg13g2_fill_2 FILLER_27_737 ();
 sg13g2_fill_1 FILLER_27_739 ();
 sg13g2_decap_8 FILLER_27_745 ();
 sg13g2_decap_8 FILLER_27_765 ();
 sg13g2_fill_1 FILLER_27_784 ();
 sg13g2_fill_2 FILLER_27_806 ();
 sg13g2_fill_1 FILLER_27_831 ();
 sg13g2_fill_1 FILLER_27_861 ();
 sg13g2_fill_1 FILLER_28_0 ();
 sg13g2_fill_1 FILLER_28_81 ();
 sg13g2_fill_2 FILLER_28_110 ();
 sg13g2_fill_1 FILLER_28_112 ();
 sg13g2_fill_2 FILLER_28_134 ();
 sg13g2_fill_1 FILLER_28_136 ();
 sg13g2_fill_2 FILLER_28_165 ();
 sg13g2_fill_1 FILLER_28_167 ();
 sg13g2_fill_2 FILLER_28_214 ();
 sg13g2_fill_1 FILLER_28_277 ();
 sg13g2_fill_1 FILLER_28_360 ();
 sg13g2_fill_1 FILLER_28_369 ();
 sg13g2_fill_2 FILLER_28_384 ();
 sg13g2_fill_2 FILLER_28_438 ();
 sg13g2_decap_4 FILLER_28_457 ();
 sg13g2_fill_1 FILLER_28_474 ();
 sg13g2_fill_1 FILLER_28_488 ();
 sg13g2_fill_1 FILLER_28_526 ();
 sg13g2_decap_8 FILLER_28_540 ();
 sg13g2_fill_1 FILLER_28_547 ();
 sg13g2_fill_2 FILLER_28_560 ();
 sg13g2_fill_2 FILLER_28_583 ();
 sg13g2_fill_1 FILLER_28_585 ();
 sg13g2_decap_8 FILLER_28_599 ();
 sg13g2_decap_4 FILLER_28_606 ();
 sg13g2_fill_2 FILLER_28_634 ();
 sg13g2_fill_1 FILLER_28_644 ();
 sg13g2_fill_2 FILLER_28_658 ();
 sg13g2_fill_1 FILLER_28_660 ();
 sg13g2_decap_4 FILLER_28_711 ();
 sg13g2_fill_2 FILLER_28_739 ();
 sg13g2_fill_2 FILLER_28_767 ();
 sg13g2_fill_1 FILLER_28_773 ();
 sg13g2_decap_4 FILLER_28_791 ();
 sg13g2_fill_1 FILLER_28_795 ();
 sg13g2_fill_2 FILLER_28_801 ();
 sg13g2_fill_1 FILLER_28_824 ();
 sg13g2_decap_8 FILLER_28_828 ();
 sg13g2_decap_8 FILLER_28_835 ();
 sg13g2_fill_2 FILLER_28_842 ();
 sg13g2_decap_4 FILLER_28_856 ();
 sg13g2_fill_2 FILLER_28_860 ();
 sg13g2_fill_1 FILLER_29_0 ();
 sg13g2_fill_1 FILLER_29_34 ();
 sg13g2_fill_2 FILLER_29_46 ();
 sg13g2_fill_2 FILLER_29_94 ();
 sg13g2_fill_1 FILLER_29_128 ();
 sg13g2_fill_1 FILLER_29_161 ();
 sg13g2_fill_1 FILLER_29_201 ();
 sg13g2_fill_1 FILLER_29_211 ();
 sg13g2_fill_2 FILLER_29_243 ();
 sg13g2_fill_2 FILLER_29_294 ();
 sg13g2_fill_1 FILLER_29_296 ();
 sg13g2_fill_1 FILLER_29_319 ();
 sg13g2_fill_2 FILLER_29_333 ();
 sg13g2_fill_1 FILLER_29_335 ();
 sg13g2_fill_1 FILLER_29_353 ();
 sg13g2_fill_2 FILLER_29_386 ();
 sg13g2_fill_1 FILLER_29_418 ();
 sg13g2_fill_2 FILLER_29_424 ();
 sg13g2_fill_1 FILLER_29_426 ();
 sg13g2_fill_1 FILLER_29_451 ();
 sg13g2_decap_4 FILLER_29_464 ();
 sg13g2_fill_1 FILLER_29_468 ();
 sg13g2_decap_8 FILLER_29_478 ();
 sg13g2_decap_4 FILLER_29_485 ();
 sg13g2_fill_2 FILLER_29_489 ();
 sg13g2_decap_8 FILLER_29_503 ();
 sg13g2_fill_2 FILLER_29_510 ();
 sg13g2_decap_4 FILLER_29_516 ();
 sg13g2_fill_1 FILLER_29_524 ();
 sg13g2_fill_2 FILLER_29_538 ();
 sg13g2_fill_1 FILLER_29_540 ();
 sg13g2_decap_4 FILLER_29_554 ();
 sg13g2_fill_2 FILLER_29_558 ();
 sg13g2_decap_4 FILLER_29_605 ();
 sg13g2_fill_1 FILLER_29_613 ();
 sg13g2_fill_2 FILLER_29_624 ();
 sg13g2_fill_2 FILLER_29_656 ();
 sg13g2_fill_1 FILLER_29_658 ();
 sg13g2_fill_1 FILLER_29_676 ();
 sg13g2_fill_2 FILLER_29_690 ();
 sg13g2_fill_1 FILLER_29_692 ();
 sg13g2_decap_4 FILLER_29_720 ();
 sg13g2_fill_1 FILLER_29_724 ();
 sg13g2_fill_2 FILLER_29_730 ();
 sg13g2_fill_2 FILLER_29_741 ();
 sg13g2_fill_1 FILLER_29_743 ();
 sg13g2_decap_8 FILLER_29_785 ();
 sg13g2_fill_1 FILLER_29_808 ();
 sg13g2_fill_2 FILLER_29_838 ();
 sg13g2_fill_1 FILLER_29_840 ();
 sg13g2_decap_4 FILLER_29_857 ();
 sg13g2_fill_1 FILLER_29_861 ();
 sg13g2_fill_2 FILLER_30_0 ();
 sg13g2_fill_2 FILLER_30_14 ();
 sg13g2_fill_1 FILLER_30_44 ();
 sg13g2_fill_2 FILLER_30_72 ();
 sg13g2_fill_2 FILLER_30_262 ();
 sg13g2_fill_1 FILLER_30_270 ();
 sg13g2_fill_1 FILLER_30_348 ();
 sg13g2_fill_2 FILLER_30_370 ();
 sg13g2_fill_2 FILLER_30_438 ();
 sg13g2_decap_8 FILLER_30_458 ();
 sg13g2_fill_1 FILLER_30_465 ();
 sg13g2_fill_2 FILLER_30_512 ();
 sg13g2_decap_4 FILLER_30_535 ();
 sg13g2_decap_4 FILLER_30_572 ();
 sg13g2_decap_4 FILLER_30_594 ();
 sg13g2_fill_2 FILLER_30_607 ();
 sg13g2_fill_1 FILLER_30_622 ();
 sg13g2_fill_1 FILLER_30_647 ();
 sg13g2_decap_8 FILLER_30_657 ();
 sg13g2_decap_8 FILLER_30_664 ();
 sg13g2_fill_2 FILLER_30_671 ();
 sg13g2_fill_2 FILLER_30_686 ();
 sg13g2_fill_1 FILLER_30_688 ();
 sg13g2_decap_8 FILLER_30_764 ();
 sg13g2_fill_2 FILLER_30_771 ();
 sg13g2_fill_2 FILLER_30_805 ();
 sg13g2_fill_1 FILLER_30_807 ();
 sg13g2_fill_1 FILLER_30_821 ();
 sg13g2_fill_2 FILLER_30_834 ();
 sg13g2_fill_1 FILLER_30_836 ();
 sg13g2_decap_4 FILLER_30_857 ();
 sg13g2_fill_1 FILLER_30_861 ();
 sg13g2_fill_2 FILLER_31_27 ();
 sg13g2_fill_2 FILLER_31_56 ();
 sg13g2_fill_2 FILLER_31_75 ();
 sg13g2_fill_2 FILLER_31_146 ();
 sg13g2_fill_1 FILLER_31_190 ();
 sg13g2_fill_1 FILLER_31_219 ();
 sg13g2_fill_1 FILLER_31_236 ();
 sg13g2_fill_1 FILLER_31_245 ();
 sg13g2_fill_1 FILLER_31_391 ();
 sg13g2_fill_1 FILLER_31_418 ();
 sg13g2_fill_2 FILLER_31_441 ();
 sg13g2_fill_1 FILLER_31_443 ();
 sg13g2_decap_4 FILLER_31_454 ();
 sg13g2_decap_8 FILLER_31_486 ();
 sg13g2_fill_2 FILLER_31_498 ();
 sg13g2_fill_2 FILLER_31_516 ();
 sg13g2_decap_4 FILLER_31_531 ();
 sg13g2_fill_1 FILLER_31_535 ();
 sg13g2_fill_1 FILLER_31_554 ();
 sg13g2_fill_2 FILLER_31_560 ();
 sg13g2_fill_1 FILLER_31_562 ();
 sg13g2_decap_4 FILLER_31_622 ();
 sg13g2_fill_1 FILLER_31_626 ();
 sg13g2_decap_8 FILLER_31_637 ();
 sg13g2_fill_1 FILLER_31_665 ();
 sg13g2_fill_1 FILLER_31_675 ();
 sg13g2_fill_2 FILLER_31_686 ();
 sg13g2_fill_1 FILLER_31_704 ();
 sg13g2_decap_8 FILLER_31_722 ();
 sg13g2_decap_4 FILLER_31_729 ();
 sg13g2_decap_8 FILLER_31_747 ();
 sg13g2_fill_2 FILLER_31_793 ();
 sg13g2_fill_1 FILLER_31_795 ();
 sg13g2_fill_1 FILLER_31_800 ();
 sg13g2_decap_8 FILLER_31_822 ();
 sg13g2_fill_1 FILLER_31_829 ();
 sg13g2_decap_4 FILLER_31_856 ();
 sg13g2_fill_2 FILLER_31_860 ();
 sg13g2_fill_1 FILLER_32_0 ();
 sg13g2_fill_2 FILLER_32_17 ();
 sg13g2_fill_2 FILLER_32_46 ();
 sg13g2_fill_2 FILLER_32_71 ();
 sg13g2_fill_2 FILLER_32_92 ();
 sg13g2_fill_1 FILLER_32_94 ();
 sg13g2_fill_1 FILLER_32_114 ();
 sg13g2_fill_2 FILLER_32_176 ();
 sg13g2_fill_2 FILLER_32_184 ();
 sg13g2_fill_1 FILLER_32_186 ();
 sg13g2_fill_2 FILLER_32_257 ();
 sg13g2_fill_1 FILLER_32_360 ();
 sg13g2_fill_1 FILLER_32_408 ();
 sg13g2_decap_8 FILLER_32_447 ();
 sg13g2_decap_4 FILLER_32_459 ();
 sg13g2_fill_1 FILLER_32_463 ();
 sg13g2_fill_1 FILLER_32_476 ();
 sg13g2_decap_4 FILLER_32_484 ();
 sg13g2_fill_1 FILLER_32_488 ();
 sg13g2_decap_8 FILLER_32_523 ();
 sg13g2_fill_2 FILLER_32_543 ();
 sg13g2_fill_1 FILLER_32_545 ();
 sg13g2_decap_8 FILLER_32_580 ();
 sg13g2_decap_8 FILLER_32_591 ();
 sg13g2_fill_1 FILLER_32_598 ();
 sg13g2_decap_4 FILLER_32_612 ();
 sg13g2_fill_1 FILLER_32_616 ();
 sg13g2_decap_4 FILLER_32_644 ();
 sg13g2_fill_2 FILLER_32_656 ();
 sg13g2_fill_1 FILLER_32_658 ();
 sg13g2_fill_1 FILLER_32_681 ();
 sg13g2_decap_4 FILLER_32_691 ();
 sg13g2_fill_1 FILLER_32_695 ();
 sg13g2_decap_4 FILLER_32_721 ();
 sg13g2_fill_1 FILLER_32_725 ();
 sg13g2_fill_2 FILLER_32_734 ();
 sg13g2_fill_2 FILLER_32_757 ();
 sg13g2_decap_4 FILLER_32_763 ();
 sg13g2_decap_4 FILLER_32_770 ();
 sg13g2_decap_8 FILLER_32_786 ();
 sg13g2_decap_4 FILLER_32_793 ();
 sg13g2_decap_8 FILLER_32_818 ();
 sg13g2_fill_2 FILLER_32_825 ();
 sg13g2_decap_4 FILLER_32_840 ();
 sg13g2_fill_1 FILLER_32_844 ();
 sg13g2_decap_4 FILLER_32_857 ();
 sg13g2_fill_1 FILLER_32_861 ();
 sg13g2_fill_1 FILLER_33_0 ();
 sg13g2_fill_2 FILLER_33_67 ();
 sg13g2_fill_2 FILLER_33_82 ();
 sg13g2_fill_2 FILLER_33_121 ();
 sg13g2_fill_2 FILLER_33_213 ();
 sg13g2_fill_2 FILLER_33_230 ();
 sg13g2_fill_1 FILLER_33_232 ();
 sg13g2_fill_2 FILLER_33_259 ();
 sg13g2_fill_1 FILLER_33_294 ();
 sg13g2_fill_2 FILLER_33_356 ();
 sg13g2_fill_1 FILLER_33_376 ();
 sg13g2_fill_2 FILLER_33_417 ();
 sg13g2_decap_8 FILLER_33_440 ();
 sg13g2_decap_4 FILLER_33_475 ();
 sg13g2_fill_1 FILLER_33_479 ();
 sg13g2_fill_1 FILLER_33_493 ();
 sg13g2_fill_2 FILLER_33_518 ();
 sg13g2_decap_8 FILLER_33_543 ();
 sg13g2_decap_4 FILLER_33_550 ();
 sg13g2_decap_4 FILLER_33_566 ();
 sg13g2_decap_4 FILLER_33_574 ();
 sg13g2_fill_1 FILLER_33_578 ();
 sg13g2_decap_4 FILLER_33_583 ();
 sg13g2_fill_1 FILLER_33_587 ();
 sg13g2_decap_4 FILLER_33_613 ();
 sg13g2_fill_1 FILLER_33_617 ();
 sg13g2_decap_4 FILLER_33_645 ();
 sg13g2_fill_2 FILLER_33_649 ();
 sg13g2_fill_2 FILLER_33_663 ();
 sg13g2_fill_1 FILLER_33_665 ();
 sg13g2_fill_2 FILLER_33_674 ();
 sg13g2_decap_8 FILLER_33_697 ();
 sg13g2_fill_1 FILLER_33_704 ();
 sg13g2_fill_2 FILLER_33_740 ();
 sg13g2_decap_4 FILLER_33_746 ();
 sg13g2_fill_1 FILLER_33_750 ();
 sg13g2_decap_4 FILLER_33_764 ();
 sg13g2_decap_4 FILLER_33_785 ();
 sg13g2_decap_4 FILLER_33_811 ();
 sg13g2_fill_1 FILLER_33_818 ();
 sg13g2_fill_2 FILLER_33_835 ();
 sg13g2_fill_1 FILLER_33_837 ();
 sg13g2_fill_2 FILLER_33_859 ();
 sg13g2_fill_1 FILLER_33_861 ();
 sg13g2_fill_1 FILLER_34_4 ();
 sg13g2_fill_1 FILLER_34_9 ();
 sg13g2_fill_2 FILLER_34_25 ();
 sg13g2_fill_2 FILLER_34_54 ();
 sg13g2_fill_1 FILLER_34_56 ();
 sg13g2_fill_1 FILLER_34_67 ();
 sg13g2_fill_2 FILLER_34_73 ();
 sg13g2_fill_1 FILLER_34_75 ();
 sg13g2_fill_2 FILLER_34_102 ();
 sg13g2_fill_1 FILLER_34_141 ();
 sg13g2_fill_2 FILLER_34_229 ();
 sg13g2_fill_2 FILLER_34_274 ();
 sg13g2_fill_2 FILLER_34_289 ();
 sg13g2_fill_1 FILLER_34_291 ();
 sg13g2_fill_1 FILLER_34_396 ();
 sg13g2_fill_2 FILLER_34_431 ();
 sg13g2_fill_1 FILLER_34_441 ();
 sg13g2_fill_2 FILLER_34_463 ();
 sg13g2_decap_8 FILLER_34_478 ();
 sg13g2_decap_4 FILLER_34_485 ();
 sg13g2_fill_1 FILLER_34_489 ();
 sg13g2_decap_4 FILLER_34_502 ();
 sg13g2_fill_1 FILLER_34_536 ();
 sg13g2_fill_2 FILLER_34_546 ();
 sg13g2_fill_1 FILLER_34_548 ();
 sg13g2_decap_4 FILLER_34_562 ();
 sg13g2_decap_4 FILLER_34_592 ();
 sg13g2_fill_1 FILLER_34_596 ();
 sg13g2_fill_2 FILLER_34_622 ();
 sg13g2_fill_2 FILLER_34_645 ();
 sg13g2_fill_1 FILLER_34_655 ();
 sg13g2_fill_1 FILLER_34_667 ();
 sg13g2_decap_8 FILLER_34_671 ();
 sg13g2_fill_1 FILLER_34_678 ();
 sg13g2_decap_8 FILLER_34_688 ();
 sg13g2_decap_8 FILLER_34_695 ();
 sg13g2_decap_4 FILLER_34_702 ();
 sg13g2_decap_4 FILLER_34_722 ();
 sg13g2_fill_2 FILLER_34_734 ();
 sg13g2_fill_2 FILLER_34_760 ();
 sg13g2_fill_1 FILLER_34_762 ();
 sg13g2_fill_1 FILLER_34_799 ();
 sg13g2_decap_8 FILLER_34_805 ();
 sg13g2_decap_4 FILLER_34_812 ();
 sg13g2_fill_2 FILLER_34_821 ();
 sg13g2_fill_1 FILLER_34_823 ();
 sg13g2_fill_2 FILLER_34_845 ();
 sg13g2_fill_2 FILLER_34_859 ();
 sg13g2_fill_1 FILLER_34_861 ();
 sg13g2_fill_2 FILLER_35_8 ();
 sg13g2_fill_1 FILLER_35_32 ();
 sg13g2_fill_2 FILLER_35_85 ();
 sg13g2_fill_2 FILLER_35_111 ();
 sg13g2_fill_1 FILLER_35_151 ();
 sg13g2_decap_4 FILLER_35_201 ();
 sg13g2_fill_1 FILLER_35_205 ();
 sg13g2_fill_2 FILLER_35_229 ();
 sg13g2_fill_2 FILLER_35_239 ();
 sg13g2_fill_1 FILLER_35_260 ();
 sg13g2_fill_2 FILLER_35_282 ();
 sg13g2_fill_1 FILLER_35_284 ();
 sg13g2_fill_2 FILLER_35_344 ();
 sg13g2_fill_1 FILLER_35_372 ();
 sg13g2_fill_2 FILLER_35_390 ();
 sg13g2_decap_8 FILLER_35_477 ();
 sg13g2_fill_2 FILLER_35_484 ();
 sg13g2_fill_2 FILLER_35_521 ();
 sg13g2_fill_2 FILLER_35_531 ();
 sg13g2_decap_4 FILLER_35_549 ();
 sg13g2_fill_1 FILLER_35_553 ();
 sg13g2_fill_2 FILLER_35_581 ();
 sg13g2_fill_1 FILLER_35_583 ();
 sg13g2_fill_2 FILLER_35_614 ();
 sg13g2_fill_2 FILLER_35_638 ();
 sg13g2_fill_1 FILLER_35_640 ();
 sg13g2_decap_4 FILLER_35_662 ();
 sg13g2_fill_1 FILLER_35_666 ();
 sg13g2_fill_2 FILLER_35_708 ();
 sg13g2_fill_1 FILLER_35_710 ();
 sg13g2_fill_2 FILLER_35_716 ();
 sg13g2_decap_8 FILLER_35_730 ();
 sg13g2_fill_2 FILLER_35_737 ();
 sg13g2_fill_1 FILLER_35_739 ();
 sg13g2_fill_1 FILLER_35_750 ();
 sg13g2_decap_8 FILLER_35_759 ();
 sg13g2_fill_2 FILLER_35_766 ();
 sg13g2_fill_1 FILLER_35_781 ();
 sg13g2_fill_2 FILLER_35_811 ();
 sg13g2_fill_2 FILLER_35_837 ();
 sg13g2_fill_1 FILLER_35_839 ();
 sg13g2_fill_1 FILLER_35_861 ();
 sg13g2_fill_1 FILLER_36_0 ();
 sg13g2_fill_2 FILLER_36_49 ();
 sg13g2_fill_2 FILLER_36_60 ();
 sg13g2_fill_2 FILLER_36_67 ();
 sg13g2_fill_1 FILLER_36_69 ();
 sg13g2_fill_1 FILLER_36_80 ();
 sg13g2_fill_1 FILLER_36_85 ();
 sg13g2_fill_2 FILLER_36_98 ();
 sg13g2_fill_1 FILLER_36_100 ();
 sg13g2_fill_1 FILLER_36_122 ();
 sg13g2_fill_2 FILLER_36_174 ();
 sg13g2_fill_2 FILLER_36_184 ();
 sg13g2_fill_1 FILLER_36_186 ();
 sg13g2_decap_8 FILLER_36_191 ();
 sg13g2_decap_4 FILLER_36_198 ();
 sg13g2_fill_2 FILLER_36_202 ();
 sg13g2_fill_2 FILLER_36_216 ();
 sg13g2_fill_2 FILLER_36_239 ();
 sg13g2_fill_1 FILLER_36_258 ();
 sg13g2_fill_2 FILLER_36_268 ();
 sg13g2_fill_2 FILLER_36_301 ();
 sg13g2_fill_1 FILLER_36_303 ();
 sg13g2_fill_1 FILLER_36_319 ();
 sg13g2_fill_2 FILLER_36_333 ();
 sg13g2_fill_1 FILLER_36_335 ();
 sg13g2_fill_2 FILLER_36_371 ();
 sg13g2_fill_2 FILLER_36_399 ();
 sg13g2_decap_4 FILLER_36_404 ();
 sg13g2_fill_1 FILLER_36_433 ();
 sg13g2_fill_2 FILLER_36_452 ();
 sg13g2_fill_1 FILLER_36_454 ();
 sg13g2_decap_4 FILLER_36_463 ();
 sg13g2_fill_2 FILLER_36_476 ();
 sg13g2_decap_8 FILLER_36_487 ();
 sg13g2_decap_4 FILLER_36_494 ();
 sg13g2_fill_2 FILLER_36_511 ();
 sg13g2_fill_1 FILLER_36_513 ();
 sg13g2_fill_1 FILLER_36_518 ();
 sg13g2_decap_4 FILLER_36_535 ();
 sg13g2_fill_1 FILLER_36_539 ();
 sg13g2_fill_1 FILLER_36_548 ();
 sg13g2_decap_8 FILLER_36_578 ();
 sg13g2_decap_4 FILLER_36_585 ();
 sg13g2_fill_1 FILLER_36_589 ();
 sg13g2_fill_2 FILLER_36_598 ();
 sg13g2_fill_1 FILLER_36_600 ();
 sg13g2_decap_4 FILLER_36_615 ();
 sg13g2_decap_8 FILLER_36_631 ();
 sg13g2_fill_2 FILLER_36_638 ();
 sg13g2_fill_1 FILLER_36_645 ();
 sg13g2_decap_8 FILLER_36_656 ();
 sg13g2_fill_1 FILLER_36_663 ();
 sg13g2_fill_2 FILLER_36_688 ();
 sg13g2_fill_1 FILLER_36_715 ();
 sg13g2_decap_8 FILLER_36_726 ();
 sg13g2_decap_8 FILLER_36_733 ();
 sg13g2_fill_2 FILLER_36_740 ();
 sg13g2_fill_2 FILLER_36_763 ();
 sg13g2_fill_1 FILLER_36_765 ();
 sg13g2_fill_1 FILLER_36_783 ();
 sg13g2_fill_2 FILLER_36_792 ();
 sg13g2_fill_1 FILLER_36_798 ();
 sg13g2_decap_8 FILLER_36_804 ();
 sg13g2_decap_4 FILLER_36_811 ();
 sg13g2_fill_2 FILLER_36_834 ();
 sg13g2_fill_1 FILLER_36_836 ();
 sg13g2_decap_8 FILLER_36_853 ();
 sg13g2_fill_2 FILLER_36_860 ();
 sg13g2_fill_2 FILLER_37_0 ();
 sg13g2_fill_1 FILLER_37_42 ();
 sg13g2_fill_1 FILLER_37_74 ();
 sg13g2_fill_2 FILLER_37_100 ();
 sg13g2_fill_1 FILLER_37_102 ();
 sg13g2_fill_1 FILLER_37_154 ();
 sg13g2_fill_2 FILLER_37_185 ();
 sg13g2_fill_1 FILLER_37_187 ();
 sg13g2_fill_2 FILLER_37_211 ();
 sg13g2_fill_1 FILLER_37_213 ();
 sg13g2_fill_2 FILLER_37_226 ();
 sg13g2_decap_4 FILLER_37_235 ();
 sg13g2_fill_1 FILLER_37_273 ();
 sg13g2_decap_8 FILLER_37_306 ();
 sg13g2_fill_1 FILLER_37_313 ();
 sg13g2_fill_2 FILLER_37_327 ();
 sg13g2_fill_2 FILLER_37_392 ();
 sg13g2_fill_1 FILLER_37_421 ();
 sg13g2_fill_2 FILLER_37_468 ();
 sg13g2_fill_1 FILLER_37_470 ();
 sg13g2_fill_1 FILLER_37_502 ();
 sg13g2_decap_4 FILLER_37_507 ();
 sg13g2_fill_1 FILLER_37_511 ();
 sg13g2_fill_1 FILLER_37_520 ();
 sg13g2_fill_1 FILLER_37_542 ();
 sg13g2_decap_8 FILLER_37_572 ();
 sg13g2_decap_4 FILLER_37_579 ();
 sg13g2_decap_4 FILLER_37_607 ();
 sg13g2_fill_1 FILLER_37_611 ();
 sg13g2_fill_1 FILLER_37_632 ();
 sg13g2_decap_4 FILLER_37_653 ();
 sg13g2_fill_2 FILLER_37_657 ();
 sg13g2_fill_2 FILLER_37_662 ();
 sg13g2_decap_4 FILLER_37_681 ();
 sg13g2_fill_1 FILLER_37_685 ();
 sg13g2_decap_4 FILLER_37_699 ();
 sg13g2_fill_2 FILLER_37_719 ();
 sg13g2_decap_4 FILLER_37_729 ();
 sg13g2_decap_4 FILLER_37_759 ();
 sg13g2_fill_2 FILLER_37_763 ();
 sg13g2_decap_8 FILLER_37_790 ();
 sg13g2_fill_2 FILLER_37_805 ();
 sg13g2_decap_8 FILLER_37_828 ();
 sg13g2_fill_2 FILLER_37_840 ();
 sg13g2_fill_1 FILLER_37_842 ();
 sg13g2_fill_2 FILLER_37_860 ();
 sg13g2_fill_2 FILLER_38_0 ();
 sg13g2_fill_2 FILLER_38_33 ();
 sg13g2_fill_2 FILLER_38_53 ();
 sg13g2_fill_1 FILLER_38_98 ();
 sg13g2_fill_2 FILLER_38_126 ();
 sg13g2_fill_2 FILLER_38_136 ();
 sg13g2_fill_1 FILLER_38_152 ();
 sg13g2_fill_2 FILLER_38_161 ();
 sg13g2_fill_1 FILLER_38_215 ();
 sg13g2_fill_1 FILLER_38_228 ();
 sg13g2_fill_1 FILLER_38_234 ();
 sg13g2_fill_2 FILLER_38_271 ();
 sg13g2_fill_1 FILLER_38_273 ();
 sg13g2_fill_2 FILLER_38_282 ();
 sg13g2_decap_4 FILLER_38_438 ();
 sg13g2_fill_2 FILLER_38_478 ();
 sg13g2_decap_4 FILLER_38_501 ();
 sg13g2_fill_2 FILLER_38_538 ();
 sg13g2_fill_1 FILLER_38_540 ();
 sg13g2_fill_2 FILLER_38_561 ();
 sg13g2_fill_2 FILLER_38_567 ();
 sg13g2_fill_2 FILLER_38_574 ();
 sg13g2_decap_8 FILLER_38_601 ();
 sg13g2_fill_1 FILLER_38_608 ();
 sg13g2_fill_1 FILLER_38_622 ();
 sg13g2_decap_4 FILLER_38_637 ();
 sg13g2_fill_2 FILLER_38_641 ();
 sg13g2_fill_2 FILLER_38_650 ();
 sg13g2_fill_1 FILLER_38_652 ();
 sg13g2_fill_2 FILLER_38_678 ();
 sg13g2_fill_1 FILLER_38_680 ();
 sg13g2_fill_2 FILLER_38_698 ();
 sg13g2_fill_2 FILLER_38_704 ();
 sg13g2_decap_8 FILLER_38_728 ();
 sg13g2_decap_8 FILLER_38_735 ();
 sg13g2_fill_2 FILLER_38_749 ();
 sg13g2_fill_1 FILLER_38_751 ();
 sg13g2_fill_2 FILLER_38_760 ();
 sg13g2_fill_1 FILLER_38_762 ();
 sg13g2_fill_2 FILLER_38_784 ();
 sg13g2_fill_1 FILLER_38_786 ();
 sg13g2_fill_2 FILLER_38_822 ();
 sg13g2_fill_1 FILLER_38_824 ();
 sg13g2_fill_2 FILLER_38_846 ();
 sg13g2_fill_2 FILLER_38_860 ();
 sg13g2_fill_2 FILLER_39_4 ();
 sg13g2_fill_1 FILLER_39_27 ();
 sg13g2_fill_2 FILLER_39_71 ();
 sg13g2_fill_2 FILLER_39_107 ();
 sg13g2_fill_2 FILLER_39_133 ();
 sg13g2_fill_2 FILLER_39_158 ();
 sg13g2_fill_2 FILLER_39_206 ();
 sg13g2_fill_1 FILLER_39_208 ();
 sg13g2_fill_1 FILLER_39_214 ();
 sg13g2_fill_2 FILLER_39_240 ();
 sg13g2_fill_2 FILLER_39_270 ();
 sg13g2_fill_1 FILLER_39_329 ();
 sg13g2_fill_1 FILLER_39_403 ();
 sg13g2_fill_1 FILLER_39_413 ();
 sg13g2_fill_1 FILLER_39_441 ();
 sg13g2_decap_8 FILLER_39_483 ();
 sg13g2_fill_2 FILLER_39_519 ();
 sg13g2_fill_1 FILLER_39_531 ();
 sg13g2_decap_4 FILLER_39_553 ();
 sg13g2_fill_1 FILLER_39_557 ();
 sg13g2_fill_2 FILLER_39_579 ();
 sg13g2_decap_8 FILLER_39_624 ();
 sg13g2_fill_1 FILLER_39_631 ();
 sg13g2_decap_8 FILLER_39_647 ();
 sg13g2_decap_4 FILLER_39_654 ();
 sg13g2_fill_1 FILLER_39_662 ();
 sg13g2_fill_1 FILLER_39_667 ();
 sg13g2_decap_8 FILLER_39_692 ();
 sg13g2_fill_1 FILLER_39_717 ();
 sg13g2_fill_2 FILLER_39_748 ();
 sg13g2_fill_2 FILLER_39_759 ();
 sg13g2_fill_1 FILLER_39_761 ();
 sg13g2_fill_1 FILLER_39_766 ();
 sg13g2_fill_2 FILLER_39_781 ();
 sg13g2_decap_4 FILLER_39_788 ();
 sg13g2_fill_2 FILLER_39_797 ();
 sg13g2_decap_4 FILLER_39_817 ();
 sg13g2_fill_2 FILLER_39_833 ();
 sg13g2_fill_1 FILLER_39_847 ();
 sg13g2_fill_2 FILLER_39_860 ();
 sg13g2_fill_1 FILLER_40_26 ();
 sg13g2_fill_1 FILLER_40_52 ();
 sg13g2_fill_2 FILLER_40_76 ();
 sg13g2_fill_1 FILLER_40_78 ();
 sg13g2_fill_2 FILLER_40_100 ();
 sg13g2_fill_1 FILLER_40_102 ();
 sg13g2_fill_2 FILLER_40_107 ();
 sg13g2_fill_1 FILLER_40_131 ();
 sg13g2_fill_2 FILLER_40_201 ();
 sg13g2_fill_1 FILLER_40_243 ();
 sg13g2_fill_2 FILLER_40_292 ();
 sg13g2_fill_1 FILLER_40_294 ();
 sg13g2_fill_2 FILLER_40_315 ();
 sg13g2_fill_2 FILLER_40_335 ();
 sg13g2_fill_2 FILLER_40_355 ();
 sg13g2_fill_1 FILLER_40_357 ();
 sg13g2_fill_1 FILLER_40_413 ();
 sg13g2_fill_2 FILLER_40_459 ();
 sg13g2_decap_4 FILLER_40_474 ();
 sg13g2_fill_1 FILLER_40_478 ();
 sg13g2_fill_2 FILLER_40_500 ();
 sg13g2_fill_1 FILLER_40_502 ();
 sg13g2_decap_8 FILLER_40_548 ();
 sg13g2_fill_1 FILLER_40_555 ();
 sg13g2_fill_2 FILLER_40_568 ();
 sg13g2_fill_2 FILLER_40_574 ();
 sg13g2_fill_1 FILLER_40_576 ();
 sg13g2_fill_2 FILLER_40_581 ();
 sg13g2_fill_1 FILLER_40_583 ();
 sg13g2_fill_2 FILLER_40_596 ();
 sg13g2_fill_2 FILLER_40_632 ();
 sg13g2_decap_8 FILLER_40_673 ();
 sg13g2_fill_1 FILLER_40_680 ();
 sg13g2_decap_4 FILLER_40_686 ();
 sg13g2_fill_1 FILLER_40_690 ();
 sg13g2_fill_1 FILLER_40_704 ();
 sg13g2_fill_2 FILLER_40_731 ();
 sg13g2_fill_1 FILLER_40_746 ();
 sg13g2_fill_1 FILLER_40_760 ();
 sg13g2_decap_4 FILLER_40_797 ();
 sg13g2_fill_2 FILLER_40_801 ();
 sg13g2_fill_2 FILLER_40_839 ();
 sg13g2_fill_1 FILLER_40_841 ();
 sg13g2_fill_2 FILLER_40_860 ();
 sg13g2_fill_1 FILLER_41_0 ();
 sg13g2_fill_1 FILLER_41_11 ();
 sg13g2_fill_1 FILLER_41_30 ();
 sg13g2_fill_2 FILLER_41_97 ();
 sg13g2_fill_2 FILLER_41_121 ();
 sg13g2_fill_1 FILLER_41_175 ();
 sg13g2_fill_2 FILLER_41_208 ();
 sg13g2_fill_1 FILLER_41_210 ();
 sg13g2_fill_1 FILLER_41_275 ();
 sg13g2_fill_2 FILLER_41_399 ();
 sg13g2_fill_2 FILLER_41_441 ();
 sg13g2_fill_1 FILLER_41_443 ();
 sg13g2_fill_2 FILLER_41_457 ();
 sg13g2_fill_1 FILLER_41_459 ();
 sg13g2_fill_2 FILLER_41_488 ();
 sg13g2_decap_4 FILLER_41_534 ();
 sg13g2_fill_2 FILLER_41_538 ();
 sg13g2_decap_4 FILLER_41_544 ();
 sg13g2_fill_2 FILLER_41_548 ();
 sg13g2_fill_2 FILLER_41_578 ();
 sg13g2_fill_1 FILLER_41_580 ();
 sg13g2_decap_4 FILLER_41_588 ();
 sg13g2_fill_1 FILLER_41_592 ();
 sg13g2_decap_4 FILLER_41_606 ();
 sg13g2_fill_2 FILLER_41_631 ();
 sg13g2_fill_1 FILLER_41_651 ();
 sg13g2_decap_8 FILLER_41_678 ();
 sg13g2_fill_2 FILLER_41_689 ();
 sg13g2_fill_1 FILLER_41_691 ();
 sg13g2_fill_1 FILLER_41_740 ();
 sg13g2_decap_8 FILLER_41_755 ();
 sg13g2_fill_2 FILLER_41_770 ();
 sg13g2_fill_2 FILLER_41_776 ();
 sg13g2_fill_1 FILLER_41_778 ();
 sg13g2_decap_4 FILLER_41_795 ();
 sg13g2_decap_8 FILLER_41_822 ();
 sg13g2_fill_2 FILLER_41_833 ();
 sg13g2_fill_1 FILLER_41_835 ();
 sg13g2_fill_2 FILLER_41_841 ();
 sg13g2_fill_1 FILLER_41_843 ();
 sg13g2_decap_8 FILLER_41_854 ();
 sg13g2_fill_1 FILLER_41_861 ();
 sg13g2_fill_1 FILLER_42_0 ();
 sg13g2_fill_1 FILLER_42_27 ();
 sg13g2_fill_1 FILLER_42_61 ();
 sg13g2_fill_2 FILLER_42_67 ();
 sg13g2_fill_2 FILLER_42_78 ();
 sg13g2_fill_1 FILLER_42_100 ();
 sg13g2_fill_1 FILLER_42_130 ();
 sg13g2_fill_1 FILLER_42_143 ();
 sg13g2_fill_2 FILLER_42_149 ();
 sg13g2_fill_2 FILLER_42_164 ();
 sg13g2_fill_2 FILLER_42_184 ();
 sg13g2_fill_1 FILLER_42_218 ();
 sg13g2_fill_2 FILLER_42_311 ();
 sg13g2_fill_1 FILLER_42_313 ();
 sg13g2_fill_2 FILLER_42_340 ();
 sg13g2_fill_2 FILLER_42_351 ();
 sg13g2_fill_2 FILLER_42_421 ();
 sg13g2_fill_2 FILLER_42_432 ();
 sg13g2_fill_1 FILLER_42_434 ();
 sg13g2_fill_2 FILLER_42_460 ();
 sg13g2_fill_1 FILLER_42_462 ();
 sg13g2_fill_2 FILLER_42_472 ();
 sg13g2_fill_1 FILLER_42_474 ();
 sg13g2_fill_2 FILLER_42_510 ();
 sg13g2_fill_1 FILLER_42_542 ();
 sg13g2_fill_2 FILLER_42_551 ();
 sg13g2_fill_1 FILLER_42_553 ();
 sg13g2_fill_2 FILLER_42_572 ();
 sg13g2_fill_1 FILLER_42_574 ();
 sg13g2_fill_1 FILLER_42_596 ();
 sg13g2_decap_8 FILLER_42_613 ();
 sg13g2_fill_1 FILLER_42_620 ();
 sg13g2_decap_4 FILLER_42_662 ();
 sg13g2_fill_2 FILLER_42_674 ();
 sg13g2_fill_1 FILLER_42_676 ();
 sg13g2_decap_4 FILLER_42_689 ();
 sg13g2_fill_2 FILLER_42_693 ();
 sg13g2_fill_2 FILLER_42_720 ();
 sg13g2_fill_2 FILLER_42_725 ();
 sg13g2_fill_1 FILLER_42_727 ();
 sg13g2_decap_4 FILLER_42_741 ();
 sg13g2_decap_8 FILLER_42_749 ();
 sg13g2_fill_1 FILLER_42_756 ();
 sg13g2_fill_2 FILLER_42_786 ();
 sg13g2_decap_8 FILLER_42_794 ();
 sg13g2_decap_8 FILLER_42_801 ();
 sg13g2_fill_1 FILLER_42_808 ();
 sg13g2_decap_4 FILLER_42_824 ();
 sg13g2_fill_2 FILLER_42_828 ();
 sg13g2_fill_1 FILLER_42_861 ();
 sg13g2_fill_1 FILLER_43_0 ();
 sg13g2_fill_2 FILLER_43_5 ();
 sg13g2_fill_2 FILLER_43_27 ();
 sg13g2_fill_1 FILLER_43_52 ();
 sg13g2_fill_2 FILLER_43_101 ();
 sg13g2_fill_1 FILLER_43_103 ();
 sg13g2_fill_1 FILLER_43_121 ();
 sg13g2_fill_2 FILLER_43_141 ();
 sg13g2_fill_1 FILLER_43_143 ();
 sg13g2_fill_1 FILLER_43_155 ();
 sg13g2_fill_1 FILLER_43_213 ();
 sg13g2_fill_2 FILLER_43_243 ();
 sg13g2_fill_2 FILLER_43_290 ();
 sg13g2_fill_1 FILLER_43_297 ();
 sg13g2_fill_2 FILLER_43_340 ();
 sg13g2_fill_1 FILLER_43_368 ();
 sg13g2_fill_2 FILLER_43_437 ();
 sg13g2_fill_1 FILLER_43_439 ();
 sg13g2_fill_2 FILLER_43_459 ();
 sg13g2_fill_1 FILLER_43_461 ();
 sg13g2_fill_2 FILLER_43_480 ();
 sg13g2_fill_1 FILLER_43_482 ();
 sg13g2_fill_1 FILLER_43_507 ();
 sg13g2_decap_4 FILLER_43_588 ();
 sg13g2_fill_1 FILLER_43_592 ();
 sg13g2_decap_8 FILLER_43_609 ();
 sg13g2_fill_2 FILLER_43_616 ();
 sg13g2_decap_8 FILLER_43_661 ();
 sg13g2_fill_1 FILLER_43_720 ();
 sg13g2_decap_8 FILLER_43_741 ();
 sg13g2_fill_1 FILLER_43_748 ();
 sg13g2_fill_2 FILLER_43_759 ();
 sg13g2_fill_2 FILLER_43_784 ();
 sg13g2_fill_1 FILLER_43_786 ();
 sg13g2_decap_8 FILLER_43_792 ();
 sg13g2_fill_2 FILLER_43_799 ();
 sg13g2_fill_1 FILLER_43_820 ();
 sg13g2_fill_2 FILLER_43_845 ();
 sg13g2_decap_8 FILLER_43_852 ();
 sg13g2_fill_2 FILLER_43_859 ();
 sg13g2_fill_1 FILLER_43_861 ();
 sg13g2_fill_2 FILLER_44_0 ();
 sg13g2_fill_1 FILLER_44_25 ();
 sg13g2_fill_1 FILLER_44_30 ();
 sg13g2_fill_2 FILLER_44_50 ();
 sg13g2_fill_1 FILLER_44_52 ();
 sg13g2_fill_1 FILLER_44_71 ();
 sg13g2_fill_1 FILLER_44_134 ();
 sg13g2_fill_2 FILLER_44_164 ();
 sg13g2_fill_1 FILLER_44_166 ();
 sg13g2_fill_1 FILLER_44_180 ();
 sg13g2_fill_1 FILLER_44_193 ();
 sg13g2_fill_2 FILLER_44_199 ();
 sg13g2_fill_1 FILLER_44_205 ();
 sg13g2_fill_1 FILLER_44_216 ();
 sg13g2_fill_1 FILLER_44_257 ();
 sg13g2_fill_2 FILLER_44_271 ();
 sg13g2_fill_2 FILLER_44_278 ();
 sg13g2_fill_1 FILLER_44_294 ();
 sg13g2_fill_2 FILLER_44_311 ();
 sg13g2_fill_1 FILLER_44_321 ();
 sg13g2_fill_1 FILLER_44_345 ();
 sg13g2_fill_2 FILLER_44_385 ();
 sg13g2_fill_2 FILLER_44_465 ();
 sg13g2_fill_1 FILLER_44_479 ();
 sg13g2_fill_2 FILLER_44_509 ();
 sg13g2_fill_1 FILLER_44_549 ();
 sg13g2_fill_1 FILLER_44_563 ();
 sg13g2_fill_1 FILLER_44_581 ();
 sg13g2_fill_2 FILLER_44_643 ();
 sg13g2_fill_1 FILLER_44_645 ();
 sg13g2_fill_1 FILLER_44_650 ();
 sg13g2_fill_1 FILLER_44_656 ();
 sg13g2_fill_2 FILLER_44_662 ();
 sg13g2_fill_2 FILLER_44_670 ();
 sg13g2_fill_1 FILLER_44_672 ();
 sg13g2_fill_2 FILLER_44_686 ();
 sg13g2_fill_2 FILLER_44_695 ();
 sg13g2_fill_1 FILLER_44_697 ();
 sg13g2_decap_8 FILLER_44_704 ();
 sg13g2_fill_1 FILLER_44_711 ();
 sg13g2_fill_2 FILLER_44_730 ();
 sg13g2_fill_1 FILLER_44_732 ();
 sg13g2_fill_1 FILLER_44_762 ();
 sg13g2_fill_2 FILLER_44_772 ();
 sg13g2_fill_1 FILLER_44_786 ();
 sg13g2_fill_1 FILLER_44_812 ();
 sg13g2_decap_4 FILLER_44_823 ();
 sg13g2_fill_1 FILLER_44_827 ();
 sg13g2_decap_4 FILLER_44_844 ();
 sg13g2_fill_1 FILLER_44_848 ();
 sg13g2_decap_8 FILLER_44_854 ();
 sg13g2_fill_1 FILLER_44_861 ();
 sg13g2_fill_2 FILLER_45_5 ();
 sg13g2_fill_1 FILLER_45_7 ();
 sg13g2_fill_1 FILLER_45_27 ();
 sg13g2_fill_2 FILLER_45_61 ();
 sg13g2_fill_1 FILLER_45_63 ();
 sg13g2_fill_2 FILLER_45_68 ();
 sg13g2_fill_1 FILLER_45_70 ();
 sg13g2_fill_1 FILLER_45_75 ();
 sg13g2_fill_2 FILLER_45_91 ();
 sg13g2_fill_1 FILLER_45_93 ();
 sg13g2_fill_2 FILLER_45_102 ();
 sg13g2_fill_2 FILLER_45_116 ();
 sg13g2_fill_1 FILLER_45_118 ();
 sg13g2_fill_2 FILLER_45_128 ();
 sg13g2_fill_1 FILLER_45_130 ();
 sg13g2_fill_2 FILLER_45_162 ();
 sg13g2_fill_1 FILLER_45_172 ();
 sg13g2_fill_1 FILLER_45_197 ();
 sg13g2_fill_2 FILLER_45_232 ();
 sg13g2_fill_2 FILLER_45_284 ();
 sg13g2_fill_1 FILLER_45_290 ();
 sg13g2_fill_2 FILLER_45_313 ();
 sg13g2_fill_1 FILLER_45_327 ();
 sg13g2_fill_2 FILLER_45_350 ();
 sg13g2_fill_2 FILLER_45_398 ();
 sg13g2_fill_1 FILLER_45_404 ();
 sg13g2_fill_1 FILLER_45_413 ();
 sg13g2_fill_2 FILLER_45_465 ();
 sg13g2_fill_2 FILLER_45_481 ();
 sg13g2_fill_1 FILLER_45_483 ();
 sg13g2_fill_1 FILLER_45_516 ();
 sg13g2_fill_2 FILLER_45_539 ();
 sg13g2_fill_1 FILLER_45_581 ();
 sg13g2_fill_2 FILLER_45_639 ();
 sg13g2_fill_1 FILLER_45_675 ();
 sg13g2_fill_2 FILLER_45_696 ();
 sg13g2_fill_1 FILLER_45_715 ();
 sg13g2_decap_4 FILLER_45_729 ();
 sg13g2_decap_4 FILLER_45_745 ();
 sg13g2_fill_1 FILLER_45_749 ();
 sg13g2_decap_4 FILLER_45_754 ();
 sg13g2_fill_2 FILLER_45_771 ();
 sg13g2_fill_1 FILLER_45_773 ();
 sg13g2_decap_4 FILLER_45_808 ();
 sg13g2_fill_2 FILLER_45_812 ();
 sg13g2_fill_2 FILLER_45_818 ();
 sg13g2_fill_1 FILLER_45_820 ();
 sg13g2_fill_2 FILLER_45_860 ();
 sg13g2_fill_1 FILLER_46_0 ();
 sg13g2_fill_2 FILLER_46_22 ();
 sg13g2_fill_1 FILLER_46_78 ();
 sg13g2_fill_2 FILLER_46_109 ();
 sg13g2_fill_1 FILLER_46_111 ();
 sg13g2_fill_2 FILLER_46_163 ();
 sg13g2_fill_2 FILLER_46_228 ();
 sg13g2_fill_2 FILLER_46_279 ();
 sg13g2_fill_1 FILLER_46_309 ();
 sg13g2_fill_2 FILLER_46_349 ();
 sg13g2_fill_2 FILLER_46_375 ();
 sg13g2_fill_1 FILLER_46_448 ();
 sg13g2_fill_1 FILLER_46_528 ();
 sg13g2_fill_2 FILLER_46_534 ();
 sg13g2_fill_2 FILLER_46_576 ();
 sg13g2_fill_1 FILLER_46_578 ();
 sg13g2_fill_2 FILLER_46_614 ();
 sg13g2_fill_2 FILLER_46_674 ();
 sg13g2_fill_1 FILLER_46_676 ();
 sg13g2_fill_2 FILLER_46_708 ();
 sg13g2_fill_1 FILLER_46_710 ();
 sg13g2_decap_8 FILLER_46_728 ();
 sg13g2_fill_1 FILLER_46_753 ();
 sg13g2_fill_1 FILLER_46_770 ();
 sg13g2_decap_4 FILLER_46_775 ();
 sg13g2_fill_2 FILLER_46_779 ();
 sg13g2_decap_8 FILLER_46_785 ();
 sg13g2_fill_2 FILLER_46_806 ();
 sg13g2_fill_1 FILLER_46_808 ();
 sg13g2_fill_2 FILLER_46_831 ();
 sg13g2_fill_1 FILLER_46_833 ();
 sg13g2_decap_4 FILLER_46_858 ();
 sg13g2_fill_2 FILLER_47_25 ();
 sg13g2_fill_1 FILLER_47_32 ();
 sg13g2_fill_1 FILLER_47_107 ();
 sg13g2_fill_2 FILLER_47_112 ();
 sg13g2_fill_1 FILLER_47_114 ();
 sg13g2_fill_2 FILLER_47_160 ();
 sg13g2_fill_1 FILLER_47_162 ();
 sg13g2_fill_1 FILLER_47_174 ();
 sg13g2_fill_1 FILLER_47_183 ();
 sg13g2_fill_1 FILLER_47_211 ();
 sg13g2_fill_2 FILLER_47_220 ();
 sg13g2_fill_1 FILLER_47_222 ();
 sg13g2_fill_1 FILLER_47_258 ();
 sg13g2_fill_1 FILLER_47_343 ();
 sg13g2_fill_1 FILLER_47_364 ();
 sg13g2_fill_2 FILLER_47_436 ();
 sg13g2_fill_1 FILLER_47_438 ();
 sg13g2_fill_1 FILLER_47_497 ();
 sg13g2_fill_1 FILLER_47_540 ();
 sg13g2_fill_2 FILLER_47_560 ();
 sg13g2_fill_1 FILLER_47_562 ();
 sg13g2_fill_2 FILLER_47_597 ();
 sg13g2_fill_1 FILLER_47_599 ();
 sg13g2_fill_2 FILLER_47_618 ();
 sg13g2_fill_1 FILLER_47_620 ();
 sg13g2_fill_2 FILLER_47_634 ();
 sg13g2_decap_4 FILLER_47_653 ();
 sg13g2_decap_4 FILLER_47_673 ();
 sg13g2_fill_1 FILLER_47_677 ();
 sg13g2_fill_1 FILLER_47_700 ();
 sg13g2_fill_2 FILLER_47_715 ();
 sg13g2_fill_2 FILLER_47_721 ();
 sg13g2_fill_1 FILLER_47_723 ();
 sg13g2_fill_1 FILLER_47_747 ();
 sg13g2_fill_1 FILLER_47_778 ();
 sg13g2_fill_2 FILLER_47_789 ();
 sg13g2_fill_2 FILLER_47_824 ();
 sg13g2_fill_1 FILLER_47_826 ();
 sg13g2_fill_2 FILLER_47_840 ();
 sg13g2_fill_2 FILLER_47_859 ();
 sg13g2_fill_1 FILLER_47_861 ();
 sg13g2_fill_1 FILLER_48_0 ();
 sg13g2_fill_2 FILLER_48_22 ();
 sg13g2_fill_1 FILLER_48_49 ();
 sg13g2_fill_2 FILLER_48_54 ();
 sg13g2_fill_1 FILLER_48_56 ();
 sg13g2_fill_2 FILLER_48_67 ();
 sg13g2_fill_1 FILLER_48_69 ();
 sg13g2_fill_1 FILLER_48_96 ();
 sg13g2_fill_2 FILLER_48_160 ();
 sg13g2_fill_2 FILLER_48_205 ();
 sg13g2_fill_2 FILLER_48_239 ();
 sg13g2_fill_2 FILLER_48_262 ();
 sg13g2_fill_1 FILLER_48_264 ();
 sg13g2_fill_2 FILLER_48_278 ();
 sg13g2_fill_1 FILLER_48_312 ();
 sg13g2_fill_1 FILLER_48_340 ();
 sg13g2_fill_1 FILLER_48_360 ();
 sg13g2_fill_1 FILLER_48_381 ();
 sg13g2_fill_2 FILLER_48_462 ();
 sg13g2_fill_1 FILLER_48_596 ();
 sg13g2_fill_2 FILLER_48_625 ();
 sg13g2_fill_2 FILLER_48_649 ();
 sg13g2_decap_8 FILLER_48_656 ();
 sg13g2_decap_4 FILLER_48_663 ();
 sg13g2_fill_2 FILLER_48_667 ();
 sg13g2_fill_2 FILLER_48_674 ();
 sg13g2_fill_1 FILLER_48_676 ();
 sg13g2_decap_4 FILLER_48_702 ();
 sg13g2_fill_2 FILLER_48_706 ();
 sg13g2_fill_2 FILLER_48_713 ();
 sg13g2_fill_1 FILLER_48_777 ();
 sg13g2_decap_4 FILLER_48_785 ();
 sg13g2_fill_2 FILLER_48_789 ();
 sg13g2_fill_1 FILLER_48_815 ();
 sg13g2_decap_4 FILLER_48_821 ();
 sg13g2_fill_2 FILLER_48_825 ();
 sg13g2_decap_4 FILLER_48_857 ();
 sg13g2_fill_1 FILLER_48_861 ();
 sg13g2_fill_1 FILLER_49_56 ();
 sg13g2_fill_2 FILLER_49_82 ();
 sg13g2_fill_2 FILLER_49_105 ();
 sg13g2_fill_1 FILLER_49_107 ();
 sg13g2_fill_2 FILLER_49_119 ();
 sg13g2_fill_2 FILLER_49_136 ();
 sg13g2_fill_1 FILLER_49_151 ();
 sg13g2_fill_2 FILLER_49_169 ();
 sg13g2_fill_1 FILLER_49_171 ();
 sg13g2_fill_1 FILLER_49_181 ();
 sg13g2_fill_2 FILLER_49_187 ();
 sg13g2_fill_1 FILLER_49_189 ();
 sg13g2_fill_2 FILLER_49_200 ();
 sg13g2_fill_2 FILLER_49_256 ();
 sg13g2_fill_2 FILLER_49_267 ();
 sg13g2_fill_1 FILLER_49_269 ();
 sg13g2_fill_1 FILLER_49_365 ();
 sg13g2_fill_2 FILLER_49_371 ();
 sg13g2_fill_1 FILLER_49_373 ();
 sg13g2_fill_1 FILLER_49_388 ();
 sg13g2_fill_1 FILLER_49_422 ();
 sg13g2_fill_1 FILLER_49_442 ();
 sg13g2_fill_2 FILLER_49_542 ();
 sg13g2_fill_2 FILLER_49_571 ();
 sg13g2_fill_2 FILLER_49_630 ();
 sg13g2_fill_2 FILLER_49_664 ();
 sg13g2_fill_1 FILLER_49_666 ();
 sg13g2_decap_4 FILLER_49_695 ();
 sg13g2_decap_4 FILLER_49_711 ();
 sg13g2_fill_2 FILLER_49_727 ();
 sg13g2_fill_1 FILLER_49_741 ();
 sg13g2_decap_8 FILLER_49_771 ();
 sg13g2_decap_4 FILLER_49_778 ();
 sg13g2_fill_2 FILLER_49_787 ();
 sg13g2_fill_1 FILLER_49_789 ();
 sg13g2_fill_2 FILLER_49_811 ();
 sg13g2_fill_2 FILLER_49_825 ();
 sg13g2_decap_8 FILLER_49_855 ();
 sg13g2_fill_1 FILLER_50_0 ();
 sg13g2_fill_2 FILLER_50_24 ();
 sg13g2_fill_1 FILLER_50_70 ();
 sg13g2_fill_2 FILLER_50_102 ();
 sg13g2_fill_1 FILLER_50_125 ();
 sg13g2_fill_2 FILLER_50_134 ();
 sg13g2_fill_2 FILLER_50_140 ();
 sg13g2_fill_2 FILLER_50_179 ();
 sg13g2_fill_1 FILLER_50_181 ();
 sg13g2_fill_2 FILLER_50_205 ();
 sg13g2_fill_1 FILLER_50_213 ();
 sg13g2_fill_2 FILLER_50_294 ();
 sg13g2_fill_1 FILLER_50_296 ();
 sg13g2_fill_2 FILLER_50_302 ();
 sg13g2_fill_1 FILLER_50_304 ();
 sg13g2_fill_1 FILLER_50_315 ();
 sg13g2_fill_2 FILLER_50_343 ();
 sg13g2_fill_1 FILLER_50_345 ();
 sg13g2_fill_2 FILLER_50_459 ();
 sg13g2_fill_2 FILLER_50_477 ();
 sg13g2_fill_2 FILLER_50_546 ();
 sg13g2_fill_1 FILLER_50_548 ();
 sg13g2_decap_8 FILLER_50_651 ();
 sg13g2_fill_2 FILLER_50_671 ();
 sg13g2_decap_8 FILLER_50_682 ();
 sg13g2_decap_8 FILLER_50_710 ();
 sg13g2_decap_4 FILLER_50_725 ();
 sg13g2_fill_1 FILLER_50_742 ();
 sg13g2_fill_2 FILLER_50_765 ();
 sg13g2_fill_1 FILLER_50_775 ();
 sg13g2_fill_2 FILLER_50_793 ();
 sg13g2_fill_1 FILLER_50_795 ();
 sg13g2_decap_8 FILLER_50_819 ();
 sg13g2_fill_2 FILLER_50_826 ();
 sg13g2_fill_1 FILLER_50_828 ();
 sg13g2_fill_1 FILLER_50_848 ();
 sg13g2_fill_1 FILLER_51_56 ();
 sg13g2_fill_1 FILLER_51_99 ();
 sg13g2_fill_2 FILLER_51_126 ();
 sg13g2_fill_1 FILLER_51_128 ();
 sg13g2_fill_2 FILLER_51_173 ();
 sg13g2_fill_1 FILLER_51_215 ();
 sg13g2_fill_2 FILLER_51_246 ();
 sg13g2_fill_2 FILLER_51_258 ();
 sg13g2_fill_1 FILLER_51_301 ();
 sg13g2_fill_2 FILLER_51_330 ();
 sg13g2_fill_1 FILLER_51_360 ();
 sg13g2_fill_2 FILLER_51_367 ();
 sg13g2_fill_1 FILLER_51_369 ();
 sg13g2_fill_1 FILLER_51_405 ();
 sg13g2_fill_1 FILLER_51_442 ();
 sg13g2_fill_2 FILLER_51_453 ();
 sg13g2_fill_2 FILLER_51_482 ();
 sg13g2_fill_2 FILLER_51_595 ();
 sg13g2_fill_2 FILLER_51_672 ();
 sg13g2_fill_2 FILLER_51_686 ();
 sg13g2_fill_1 FILLER_51_688 ();
 sg13g2_fill_2 FILLER_51_697 ();
 sg13g2_fill_1 FILLER_51_699 ();
 sg13g2_decap_8 FILLER_51_705 ();
 sg13g2_fill_2 FILLER_51_735 ();
 sg13g2_fill_1 FILLER_51_737 ();
 sg13g2_fill_2 FILLER_51_764 ();
 sg13g2_fill_2 FILLER_51_814 ();
 sg13g2_fill_2 FILLER_51_821 ();
 sg13g2_fill_1 FILLER_51_823 ();
 sg13g2_decap_8 FILLER_51_841 ();
 sg13g2_decap_8 FILLER_51_853 ();
 sg13g2_fill_2 FILLER_51_860 ();
 sg13g2_fill_1 FILLER_52_87 ();
 sg13g2_fill_2 FILLER_52_130 ();
 sg13g2_fill_1 FILLER_52_172 ();
 sg13g2_fill_1 FILLER_52_182 ();
 sg13g2_fill_2 FILLER_52_198 ();
 sg13g2_fill_1 FILLER_52_200 ();
 sg13g2_fill_2 FILLER_52_219 ();
 sg13g2_fill_1 FILLER_52_239 ();
 sg13g2_fill_1 FILLER_52_250 ();
 sg13g2_fill_1 FILLER_52_266 ();
 sg13g2_fill_2 FILLER_52_290 ();
 sg13g2_fill_2 FILLER_52_368 ();
 sg13g2_fill_2 FILLER_52_475 ();
 sg13g2_fill_2 FILLER_52_572 ();
 sg13g2_fill_1 FILLER_52_574 ();
 sg13g2_fill_1 FILLER_52_618 ();
 sg13g2_fill_1 FILLER_52_628 ();
 sg13g2_fill_2 FILLER_52_634 ();
 sg13g2_fill_2 FILLER_52_666 ();
 sg13g2_decap_8 FILLER_52_694 ();
 sg13g2_fill_1 FILLER_52_701 ();
 sg13g2_fill_2 FILLER_52_719 ();
 sg13g2_fill_2 FILLER_52_728 ();
 sg13g2_fill_1 FILLER_52_742 ();
 sg13g2_fill_2 FILLER_52_772 ();
 sg13g2_fill_1 FILLER_52_774 ();
 sg13g2_fill_2 FILLER_52_785 ();
 sg13g2_fill_1 FILLER_52_787 ();
 sg13g2_fill_2 FILLER_52_806 ();
 sg13g2_decap_4 FILLER_52_820 ();
 sg13g2_fill_2 FILLER_52_860 ();
 sg13g2_fill_1 FILLER_53_0 ();
 sg13g2_fill_1 FILLER_53_27 ();
 sg13g2_fill_2 FILLER_53_103 ();
 sg13g2_fill_2 FILLER_53_125 ();
 sg13g2_fill_1 FILLER_53_127 ();
 sg13g2_fill_2 FILLER_53_133 ();
 sg13g2_fill_2 FILLER_53_163 ();
 sg13g2_fill_1 FILLER_53_165 ();
 sg13g2_fill_2 FILLER_53_201 ();
 sg13g2_fill_1 FILLER_53_216 ();
 sg13g2_fill_2 FILLER_53_271 ();
 sg13g2_fill_1 FILLER_53_273 ();
 sg13g2_fill_2 FILLER_53_291 ();
 sg13g2_fill_1 FILLER_53_293 ();
 sg13g2_fill_2 FILLER_53_309 ();
 sg13g2_fill_1 FILLER_53_324 ();
 sg13g2_fill_2 FILLER_53_348 ();
 sg13g2_fill_2 FILLER_53_378 ();
 sg13g2_fill_2 FILLER_53_413 ();
 sg13g2_fill_1 FILLER_53_521 ();
 sg13g2_fill_2 FILLER_53_623 ();
 sg13g2_fill_1 FILLER_53_645 ();
 sg13g2_decap_4 FILLER_53_681 ();
 sg13g2_fill_1 FILLER_53_685 ();
 sg13g2_fill_2 FILLER_53_706 ();
 sg13g2_fill_2 FILLER_53_713 ();
 sg13g2_decap_8 FILLER_53_732 ();
 sg13g2_fill_1 FILLER_53_739 ();
 sg13g2_fill_2 FILLER_53_757 ();
 sg13g2_fill_1 FILLER_53_772 ();
 sg13g2_fill_2 FILLER_53_790 ();
 sg13g2_fill_1 FILLER_53_792 ();
 sg13g2_decap_4 FILLER_53_816 ();
 sg13g2_fill_2 FILLER_53_820 ();
 sg13g2_fill_2 FILLER_53_838 ();
 sg13g2_fill_1 FILLER_53_840 ();
 sg13g2_fill_2 FILLER_54_0 ();
 sg13g2_fill_2 FILLER_54_75 ();
 sg13g2_fill_1 FILLER_54_77 ();
 sg13g2_fill_2 FILLER_54_91 ();
 sg13g2_fill_1 FILLER_54_93 ();
 sg13g2_fill_1 FILLER_54_110 ();
 sg13g2_fill_2 FILLER_54_137 ();
 sg13g2_fill_2 FILLER_54_151 ();
 sg13g2_fill_1 FILLER_54_158 ();
 sg13g2_fill_1 FILLER_54_172 ();
 sg13g2_fill_1 FILLER_54_203 ();
 sg13g2_fill_1 FILLER_54_209 ();
 sg13g2_fill_1 FILLER_54_215 ();
 sg13g2_fill_1 FILLER_54_239 ();
 sg13g2_fill_1 FILLER_54_249 ();
 sg13g2_fill_1 FILLER_54_321 ();
 sg13g2_fill_2 FILLER_54_396 ();
 sg13g2_fill_1 FILLER_54_445 ();
 sg13g2_fill_1 FILLER_54_566 ();
 sg13g2_fill_1 FILLER_54_609 ();
 sg13g2_fill_2 FILLER_54_645 ();
 sg13g2_fill_2 FILLER_54_683 ();
 sg13g2_decap_4 FILLER_54_700 ();
 sg13g2_fill_2 FILLER_54_704 ();
 sg13g2_decap_8 FILLER_54_727 ();
 sg13g2_decap_4 FILLER_54_734 ();
 sg13g2_fill_2 FILLER_54_738 ();
 sg13g2_decap_4 FILLER_54_755 ();
 sg13g2_decap_8 FILLER_54_786 ();
 sg13g2_fill_2 FILLER_54_793 ();
 sg13g2_fill_2 FILLER_54_814 ();
 sg13g2_fill_1 FILLER_54_816 ();
 sg13g2_fill_2 FILLER_54_834 ();
 sg13g2_fill_1 FILLER_54_836 ();
 sg13g2_decap_4 FILLER_54_858 ();
 sg13g2_fill_2 FILLER_55_0 ();
 sg13g2_fill_2 FILLER_55_61 ();
 sg13g2_fill_1 FILLER_55_73 ();
 sg13g2_fill_2 FILLER_55_84 ();
 sg13g2_fill_1 FILLER_55_86 ();
 sg13g2_fill_1 FILLER_55_94 ();
 sg13g2_fill_2 FILLER_55_110 ();
 sg13g2_fill_1 FILLER_55_138 ();
 sg13g2_fill_2 FILLER_55_169 ();
 sg13g2_fill_1 FILLER_55_171 ();
 sg13g2_fill_1 FILLER_55_201 ();
 sg13g2_fill_1 FILLER_55_225 ();
 sg13g2_fill_1 FILLER_55_411 ();
 sg13g2_fill_1 FILLER_55_475 ();
 sg13g2_fill_2 FILLER_55_507 ();
 sg13g2_fill_1 FILLER_55_656 ();
 sg13g2_fill_1 FILLER_55_676 ();
 sg13g2_fill_1 FILLER_55_697 ();
 sg13g2_decap_4 FILLER_55_707 ();
 sg13g2_fill_2 FILLER_55_711 ();
 sg13g2_fill_1 FILLER_55_734 ();
 sg13g2_fill_2 FILLER_55_754 ();
 sg13g2_fill_1 FILLER_55_756 ();
 sg13g2_fill_2 FILLER_55_771 ();
 sg13g2_fill_1 FILLER_55_773 ();
 sg13g2_fill_1 FILLER_55_777 ();
 sg13g2_decap_8 FILLER_55_783 ();
 sg13g2_decap_4 FILLER_55_790 ();
 sg13g2_fill_2 FILLER_55_794 ();
 sg13g2_fill_2 FILLER_55_806 ();
 sg13g2_fill_1 FILLER_55_808 ();
 sg13g2_decap_8 FILLER_55_831 ();
 sg13g2_fill_1 FILLER_55_838 ();
 sg13g2_fill_1 FILLER_55_848 ();
 sg13g2_fill_2 FILLER_56_0 ();
 sg13g2_fill_1 FILLER_56_2 ();
 sg13g2_fill_2 FILLER_56_27 ();
 sg13g2_fill_2 FILLER_56_36 ();
 sg13g2_fill_1 FILLER_56_82 ();
 sg13g2_fill_1 FILLER_56_121 ();
 sg13g2_fill_2 FILLER_56_155 ();
 sg13g2_fill_2 FILLER_56_205 ();
 sg13g2_fill_1 FILLER_56_251 ();
 sg13g2_fill_1 FILLER_56_458 ();
 sg13g2_fill_2 FILLER_56_557 ();
 sg13g2_fill_2 FILLER_56_572 ();
 sg13g2_fill_2 FILLER_56_596 ();
 sg13g2_fill_2 FILLER_56_707 ();
 sg13g2_fill_1 FILLER_56_709 ();
 sg13g2_fill_1 FILLER_56_715 ();
 sg13g2_fill_2 FILLER_56_724 ();
 sg13g2_fill_1 FILLER_56_726 ();
 sg13g2_fill_1 FILLER_56_732 ();
 sg13g2_fill_2 FILLER_56_774 ();
 sg13g2_fill_2 FILLER_56_792 ();
 sg13g2_fill_1 FILLER_56_794 ();
 sg13g2_fill_2 FILLER_56_807 ();
 sg13g2_fill_1 FILLER_56_809 ();
 sg13g2_decap_8 FILLER_56_817 ();
 sg13g2_decap_8 FILLER_56_824 ();
 sg13g2_fill_2 FILLER_56_831 ();
 sg13g2_fill_1 FILLER_56_833 ();
 sg13g2_decap_4 FILLER_56_856 ();
 sg13g2_fill_2 FILLER_56_860 ();
 sg13g2_fill_1 FILLER_57_100 ();
 sg13g2_fill_1 FILLER_57_162 ();
 sg13g2_fill_2 FILLER_57_207 ();
 sg13g2_fill_2 FILLER_57_308 ();
 sg13g2_fill_2 FILLER_57_332 ();
 sg13g2_fill_1 FILLER_57_334 ();
 sg13g2_fill_2 FILLER_57_353 ();
 sg13g2_fill_1 FILLER_57_355 ();
 sg13g2_fill_1 FILLER_57_415 ();
 sg13g2_fill_2 FILLER_57_443 ();
 sg13g2_fill_1 FILLER_57_617 ();
 sg13g2_fill_1 FILLER_57_650 ();
 sg13g2_fill_1 FILLER_57_675 ();
 sg13g2_fill_2 FILLER_57_684 ();
 sg13g2_fill_2 FILLER_57_698 ();
 sg13g2_decap_4 FILLER_57_720 ();
 sg13g2_fill_2 FILLER_57_757 ();
 sg13g2_fill_1 FILLER_57_759 ();
 sg13g2_fill_1 FILLER_57_821 ();
 sg13g2_fill_2 FILLER_57_860 ();
 sg13g2_fill_2 FILLER_58_65 ();
 sg13g2_fill_2 FILLER_58_121 ();
 sg13g2_fill_2 FILLER_58_147 ();
 sg13g2_fill_1 FILLER_58_162 ();
 sg13g2_fill_1 FILLER_58_394 ();
 sg13g2_fill_2 FILLER_58_409 ();
 sg13g2_fill_2 FILLER_58_425 ();
 sg13g2_fill_2 FILLER_58_618 ();
 sg13g2_fill_1 FILLER_58_620 ();
 sg13g2_fill_2 FILLER_58_631 ();
 sg13g2_fill_1 FILLER_58_633 ();
 sg13g2_fill_2 FILLER_58_655 ();
 sg13g2_decap_4 FILLER_58_714 ();
 sg13g2_fill_2 FILLER_58_718 ();
 sg13g2_fill_2 FILLER_58_724 ();
 sg13g2_decap_8 FILLER_58_734 ();
 sg13g2_fill_2 FILLER_58_741 ();
 sg13g2_fill_1 FILLER_58_743 ();
 sg13g2_decap_4 FILLER_58_754 ();
 sg13g2_fill_2 FILLER_58_778 ();
 sg13g2_fill_1 FILLER_58_808 ();
 sg13g2_fill_1 FILLER_58_833 ();
 sg13g2_decap_4 FILLER_58_856 ();
 sg13g2_fill_2 FILLER_58_860 ();
 sg13g2_fill_2 FILLER_59_223 ();
 sg13g2_fill_1 FILLER_59_265 ();
 sg13g2_fill_1 FILLER_59_299 ();
 sg13g2_fill_2 FILLER_59_378 ();
 sg13g2_fill_2 FILLER_59_427 ();
 sg13g2_fill_1 FILLER_59_429 ();
 sg13g2_fill_1 FILLER_59_690 ();
 sg13g2_fill_1 FILLER_59_717 ();
 sg13g2_decap_4 FILLER_59_734 ();
 sg13g2_decap_4 FILLER_59_757 ();
 sg13g2_fill_1 FILLER_59_761 ();
 sg13g2_fill_1 FILLER_59_770 ();
 sg13g2_decap_4 FILLER_59_776 ();
 sg13g2_decap_8 FILLER_59_787 ();
 sg13g2_fill_2 FILLER_59_794 ();
 sg13g2_decap_8 FILLER_59_823 ();
 sg13g2_fill_1 FILLER_59_861 ();
 sg13g2_fill_2 FILLER_60_0 ();
 sg13g2_fill_2 FILLER_60_57 ();
 sg13g2_fill_2 FILLER_60_68 ();
 sg13g2_fill_2 FILLER_60_161 ();
 sg13g2_fill_2 FILLER_60_194 ();
 sg13g2_fill_1 FILLER_60_385 ();
 sg13g2_fill_2 FILLER_60_395 ();
 sg13g2_fill_1 FILLER_60_500 ();
 sg13g2_fill_2 FILLER_60_542 ();
 sg13g2_fill_2 FILLER_60_649 ();
 sg13g2_fill_2 FILLER_60_681 ();
 sg13g2_fill_2 FILLER_60_720 ();
 sg13g2_fill_1 FILLER_60_722 ();
 sg13g2_fill_2 FILLER_60_728 ();
 sg13g2_decap_8 FILLER_60_751 ();
 sg13g2_fill_1 FILLER_60_758 ();
 sg13g2_decap_8 FILLER_60_784 ();
 sg13g2_fill_2 FILLER_60_803 ();
 sg13g2_fill_1 FILLER_60_805 ();
 sg13g2_decap_8 FILLER_60_815 ();
 sg13g2_decap_4 FILLER_60_822 ();
 sg13g2_fill_2 FILLER_60_830 ();
 sg13g2_decap_8 FILLER_60_853 ();
 sg13g2_fill_2 FILLER_60_860 ();
 sg13g2_fill_2 FILLER_61_0 ();
 sg13g2_fill_1 FILLER_61_112 ();
 sg13g2_fill_2 FILLER_61_129 ();
 sg13g2_fill_2 FILLER_61_212 ();
 sg13g2_fill_1 FILLER_61_238 ();
 sg13g2_fill_1 FILLER_61_410 ();
 sg13g2_fill_2 FILLER_61_433 ();
 sg13g2_fill_1 FILLER_61_511 ();
 sg13g2_fill_2 FILLER_61_594 ();
 sg13g2_fill_2 FILLER_61_635 ();
 sg13g2_fill_1 FILLER_61_637 ();
 sg13g2_fill_2 FILLER_61_643 ();
 sg13g2_fill_2 FILLER_61_679 ();
 sg13g2_fill_2 FILLER_61_707 ();
 sg13g2_fill_1 FILLER_61_709 ();
 sg13g2_fill_2 FILLER_61_725 ();
 sg13g2_fill_2 FILLER_61_732 ();
 sg13g2_decap_4 FILLER_61_747 ();
 sg13g2_fill_2 FILLER_61_751 ();
 sg13g2_fill_2 FILLER_61_758 ();
 sg13g2_decap_4 FILLER_61_765 ();
 sg13g2_decap_4 FILLER_61_786 ();
 sg13g2_fill_2 FILLER_61_802 ();
 sg13g2_fill_1 FILLER_61_804 ();
 sg13g2_fill_2 FILLER_61_821 ();
 sg13g2_fill_1 FILLER_61_823 ();
 sg13g2_fill_1 FILLER_61_861 ();
 sg13g2_fill_2 FILLER_62_42 ();
 sg13g2_fill_1 FILLER_62_57 ();
 sg13g2_fill_1 FILLER_62_73 ();
 sg13g2_fill_1 FILLER_62_141 ();
 sg13g2_fill_2 FILLER_62_192 ();
 sg13g2_fill_2 FILLER_62_284 ();
 sg13g2_fill_1 FILLER_62_286 ();
 sg13g2_fill_1 FILLER_62_402 ();
 sg13g2_fill_2 FILLER_62_524 ();
 sg13g2_fill_1 FILLER_62_618 ();
 sg13g2_fill_2 FILLER_62_640 ();
 sg13g2_fill_1 FILLER_62_642 ();
 sg13g2_fill_2 FILLER_62_648 ();
 sg13g2_fill_1 FILLER_62_664 ();
 sg13g2_fill_2 FILLER_62_698 ();
 sg13g2_fill_1 FILLER_62_700 ();
 sg13g2_fill_2 FILLER_62_716 ();
 sg13g2_fill_1 FILLER_62_718 ();
 sg13g2_fill_2 FILLER_62_748 ();
 sg13g2_fill_1 FILLER_62_758 ();
 sg13g2_fill_2 FILLER_62_766 ();
 sg13g2_decap_8 FILLER_62_780 ();
 sg13g2_decap_4 FILLER_62_787 ();
 sg13g2_fill_2 FILLER_62_814 ();
 sg13g2_fill_2 FILLER_62_833 ();
 sg13g2_fill_1 FILLER_62_835 ();
 sg13g2_fill_2 FILLER_62_860 ();
 sg13g2_fill_2 FILLER_63_32 ();
 sg13g2_fill_1 FILLER_63_203 ();
 sg13g2_fill_1 FILLER_63_231 ();
 sg13g2_fill_2 FILLER_63_272 ();
 sg13g2_fill_2 FILLER_63_326 ();
 sg13g2_fill_2 FILLER_63_400 ();
 sg13g2_fill_1 FILLER_63_536 ();
 sg13g2_fill_1 FILLER_63_585 ();
 sg13g2_fill_2 FILLER_63_628 ();
 sg13g2_fill_1 FILLER_63_684 ();
 sg13g2_fill_2 FILLER_63_691 ();
 sg13g2_fill_1 FILLER_63_693 ();
 sg13g2_fill_2 FILLER_63_727 ();
 sg13g2_fill_1 FILLER_63_736 ();
 sg13g2_fill_1 FILLER_63_749 ();
 sg13g2_decap_4 FILLER_63_755 ();
 sg13g2_fill_2 FILLER_63_768 ();
 sg13g2_fill_2 FILLER_63_775 ();
 sg13g2_fill_1 FILLER_63_777 ();
 sg13g2_fill_2 FILLER_63_783 ();
 sg13g2_fill_1 FILLER_63_785 ();
 sg13g2_decap_8 FILLER_63_830 ();
 sg13g2_fill_1 FILLER_64_38 ();
 sg13g2_fill_1 FILLER_64_100 ();
 sg13g2_fill_1 FILLER_64_137 ();
 sg13g2_fill_1 FILLER_64_236 ();
 sg13g2_fill_2 FILLER_64_295 ();
 sg13g2_fill_2 FILLER_64_379 ();
 sg13g2_fill_1 FILLER_64_482 ();
 sg13g2_fill_1 FILLER_64_502 ();
 sg13g2_fill_2 FILLER_64_639 ();
 sg13g2_fill_1 FILLER_64_641 ();
 sg13g2_fill_1 FILLER_64_666 ();
 sg13g2_fill_2 FILLER_64_708 ();
 sg13g2_fill_1 FILLER_64_710 ();
 sg13g2_fill_2 FILLER_64_727 ();
 sg13g2_fill_2 FILLER_64_737 ();
 sg13g2_fill_1 FILLER_64_739 ();
 sg13g2_fill_2 FILLER_64_764 ();
 sg13g2_fill_1 FILLER_64_766 ();
 sg13g2_decap_4 FILLER_64_782 ();
 sg13g2_decap_8 FILLER_64_798 ();
 sg13g2_fill_1 FILLER_64_805 ();
 sg13g2_decap_4 FILLER_64_811 ();
 sg13g2_fill_2 FILLER_64_815 ();
 sg13g2_decap_8 FILLER_64_822 ();
 sg13g2_fill_2 FILLER_64_829 ();
 sg13g2_decap_4 FILLER_64_856 ();
 sg13g2_fill_2 FILLER_64_860 ();
 sg13g2_fill_1 FILLER_65_0 ();
 sg13g2_fill_1 FILLER_65_33 ();
 sg13g2_fill_1 FILLER_65_388 ();
 sg13g2_fill_2 FILLER_65_491 ();
 sg13g2_fill_2 FILLER_65_534 ();
 sg13g2_fill_1 FILLER_65_536 ();
 sg13g2_fill_2 FILLER_65_565 ();
 sg13g2_fill_2 FILLER_65_626 ();
 sg13g2_fill_1 FILLER_65_717 ();
 sg13g2_fill_1 FILLER_65_725 ();
 sg13g2_fill_2 FILLER_65_751 ();
 sg13g2_fill_2 FILLER_65_758 ();
 sg13g2_fill_2 FILLER_65_765 ();
 sg13g2_fill_1 FILLER_65_798 ();
 sg13g2_decap_4 FILLER_65_804 ();
 sg13g2_fill_1 FILLER_65_808 ();
 sg13g2_fill_2 FILLER_65_821 ();
 sg13g2_fill_1 FILLER_65_823 ();
 sg13g2_decap_8 FILLER_65_849 ();
 sg13g2_decap_4 FILLER_65_856 ();
 sg13g2_fill_2 FILLER_65_860 ();
 sg13g2_fill_2 FILLER_66_32 ();
 sg13g2_fill_1 FILLER_66_43 ();
 sg13g2_fill_1 FILLER_66_72 ();
 sg13g2_fill_1 FILLER_66_141 ();
 sg13g2_fill_1 FILLER_66_212 ();
 sg13g2_fill_2 FILLER_66_317 ();
 sg13g2_fill_1 FILLER_66_332 ();
 sg13g2_fill_2 FILLER_66_460 ();
 sg13g2_fill_2 FILLER_66_544 ();
 sg13g2_fill_1 FILLER_66_546 ();
 sg13g2_fill_1 FILLER_66_560 ();
 sg13g2_fill_1 FILLER_66_574 ();
 sg13g2_fill_1 FILLER_66_580 ();
 sg13g2_fill_2 FILLER_66_609 ();
 sg13g2_fill_1 FILLER_66_611 ();
 sg13g2_fill_2 FILLER_66_623 ();
 sg13g2_fill_1 FILLER_66_625 ();
 sg13g2_fill_1 FILLER_66_652 ();
 sg13g2_fill_1 FILLER_66_680 ();
 sg13g2_fill_1 FILLER_66_685 ();
 sg13g2_fill_2 FILLER_66_691 ();
 sg13g2_fill_1 FILLER_66_693 ();
 sg13g2_fill_1 FILLER_66_711 ();
 sg13g2_fill_2 FILLER_66_727 ();
 sg13g2_fill_2 FILLER_66_741 ();
 sg13g2_fill_1 FILLER_66_743 ();
 sg13g2_fill_2 FILLER_66_785 ();
 sg13g2_fill_1 FILLER_66_787 ();
 sg13g2_fill_2 FILLER_66_795 ();
 sg13g2_fill_1 FILLER_66_797 ();
 sg13g2_fill_1 FILLER_66_822 ();
 sg13g2_fill_2 FILLER_66_841 ();
 sg13g2_fill_1 FILLER_66_843 ();
 sg13g2_decap_8 FILLER_66_855 ();
 sg13g2_fill_2 FILLER_67_32 ();
 sg13g2_fill_1 FILLER_67_43 ();
 sg13g2_fill_2 FILLER_67_59 ();
 sg13g2_fill_1 FILLER_67_70 ();
 sg13g2_fill_1 FILLER_67_89 ();
 sg13g2_fill_1 FILLER_67_142 ();
 sg13g2_fill_2 FILLER_67_248 ();
 sg13g2_fill_1 FILLER_67_314 ();
 sg13g2_fill_1 FILLER_67_464 ();
 sg13g2_fill_2 FILLER_67_602 ();
 sg13g2_fill_1 FILLER_67_604 ();
 sg13g2_fill_2 FILLER_67_634 ();
 sg13g2_fill_2 FILLER_67_642 ();
 sg13g2_fill_2 FILLER_67_663 ();
 sg13g2_fill_1 FILLER_67_665 ();
 sg13g2_fill_1 FILLER_67_704 ();
 sg13g2_fill_1 FILLER_67_713 ();
 sg13g2_fill_1 FILLER_67_719 ();
 sg13g2_fill_1 FILLER_67_729 ();
 sg13g2_fill_2 FILLER_67_751 ();
 sg13g2_fill_1 FILLER_67_753 ();
 sg13g2_fill_2 FILLER_67_771 ();
 sg13g2_decap_8 FILLER_67_786 ();
 sg13g2_decap_4 FILLER_67_793 ();
 sg13g2_decap_8 FILLER_67_810 ();
 sg13g2_decap_8 FILLER_67_817 ();
 sg13g2_fill_1 FILLER_68_41 ();
 sg13g2_fill_2 FILLER_68_181 ();
 sg13g2_fill_2 FILLER_68_196 ();
 sg13g2_fill_1 FILLER_68_230 ();
 sg13g2_fill_2 FILLER_68_318 ();
 sg13g2_fill_1 FILLER_68_379 ();
 sg13g2_fill_2 FILLER_68_389 ();
 sg13g2_fill_1 FILLER_68_546 ();
 sg13g2_fill_2 FILLER_68_643 ();
 sg13g2_fill_1 FILLER_68_720 ();
 sg13g2_fill_2 FILLER_68_759 ();
 sg13g2_fill_1 FILLER_68_761 ();
 sg13g2_fill_2 FILLER_68_784 ();
 sg13g2_fill_1 FILLER_68_786 ();
 sg13g2_fill_2 FILLER_68_795 ();
 sg13g2_decap_4 FILLER_68_818 ();
 sg13g2_fill_2 FILLER_68_822 ();
 sg13g2_fill_2 FILLER_68_832 ();
 sg13g2_decap_4 FILLER_68_858 ();
 sg13g2_fill_2 FILLER_69_31 ();
 sg13g2_fill_2 FILLER_69_87 ();
 sg13g2_fill_1 FILLER_69_154 ();
 sg13g2_fill_1 FILLER_69_183 ();
 sg13g2_fill_2 FILLER_69_211 ();
 sg13g2_fill_1 FILLER_69_460 ();
 sg13g2_fill_1 FILLER_69_554 ();
 sg13g2_fill_2 FILLER_69_574 ();
 sg13g2_fill_2 FILLER_69_606 ();
 sg13g2_fill_2 FILLER_69_637 ();
 sg13g2_fill_2 FILLER_69_665 ();
 sg13g2_fill_1 FILLER_69_667 ();
 sg13g2_fill_1 FILLER_69_686 ();
 sg13g2_fill_1 FILLER_69_708 ();
 sg13g2_fill_2 FILLER_69_714 ();
 sg13g2_fill_1 FILLER_69_721 ();
 sg13g2_fill_2 FILLER_69_741 ();
 sg13g2_fill_1 FILLER_69_764 ();
 sg13g2_fill_2 FILLER_69_782 ();
 sg13g2_fill_1 FILLER_69_784 ();
 sg13g2_decap_8 FILLER_69_822 ();
 sg13g2_decap_4 FILLER_69_829 ();
 sg13g2_fill_2 FILLER_69_859 ();
 sg13g2_fill_1 FILLER_69_861 ();
 sg13g2_fill_1 FILLER_70_51 ();
 sg13g2_fill_2 FILLER_70_184 ();
 sg13g2_fill_1 FILLER_70_199 ();
 sg13g2_fill_2 FILLER_70_233 ();
 sg13g2_fill_1 FILLER_70_414 ();
 sg13g2_fill_1 FILLER_70_433 ();
 sg13g2_fill_1 FILLER_70_447 ();
 sg13g2_fill_2 FILLER_70_483 ();
 sg13g2_fill_1 FILLER_70_533 ();
 sg13g2_fill_2 FILLER_70_540 ();
 sg13g2_fill_1 FILLER_70_571 ();
 sg13g2_fill_1 FILLER_70_603 ();
 sg13g2_fill_1 FILLER_70_617 ();
 sg13g2_fill_2 FILLER_70_650 ();
 sg13g2_fill_1 FILLER_70_652 ();
 sg13g2_fill_1 FILLER_70_666 ();
 sg13g2_fill_2 FILLER_70_696 ();
 sg13g2_fill_1 FILLER_70_766 ();
 sg13g2_fill_1 FILLER_70_771 ();
 sg13g2_fill_2 FILLER_70_785 ();
 sg13g2_fill_2 FILLER_70_808 ();
 sg13g2_fill_2 FILLER_70_826 ();
 sg13g2_fill_2 FILLER_70_840 ();
 sg13g2_fill_1 FILLER_71_72 ();
 sg13g2_fill_2 FILLER_71_87 ();
 sg13g2_fill_2 FILLER_71_104 ();
 sg13g2_fill_2 FILLER_71_156 ();
 sg13g2_fill_2 FILLER_71_194 ();
 sg13g2_fill_1 FILLER_71_209 ();
 sg13g2_fill_1 FILLER_71_255 ();
 sg13g2_fill_1 FILLER_71_321 ();
 sg13g2_fill_2 FILLER_71_365 ();
 sg13g2_fill_2 FILLER_71_376 ();
 sg13g2_fill_2 FILLER_71_432 ();
 sg13g2_fill_2 FILLER_71_503 ();
 sg13g2_fill_2 FILLER_71_548 ();
 sg13g2_fill_2 FILLER_71_596 ();
 sg13g2_fill_2 FILLER_71_622 ();
 sg13g2_fill_1 FILLER_71_624 ();
 sg13g2_fill_2 FILLER_71_706 ();
 sg13g2_fill_2 FILLER_71_721 ();
 sg13g2_fill_1 FILLER_71_723 ();
 sg13g2_fill_2 FILLER_71_733 ();
 sg13g2_fill_2 FILLER_71_743 ();
 sg13g2_fill_1 FILLER_71_750 ();
 sg13g2_fill_2 FILLER_71_759 ();
 sg13g2_fill_2 FILLER_71_795 ();
 sg13g2_fill_2 FILLER_71_809 ();
 sg13g2_decap_8 FILLER_71_834 ();
 sg13g2_fill_1 FILLER_71_841 ();
 sg13g2_decap_8 FILLER_71_854 ();
 sg13g2_fill_1 FILLER_71_861 ();
 sg13g2_fill_1 FILLER_72_30 ();
 sg13g2_fill_1 FILLER_72_86 ();
 sg13g2_fill_2 FILLER_72_155 ();
 sg13g2_fill_2 FILLER_72_264 ();
 sg13g2_fill_1 FILLER_72_419 ();
 sg13g2_fill_2 FILLER_72_484 ();
 sg13g2_fill_1 FILLER_72_564 ();
 sg13g2_fill_1 FILLER_72_601 ();
 sg13g2_fill_1 FILLER_72_619 ();
 sg13g2_fill_2 FILLER_72_638 ();
 sg13g2_fill_1 FILLER_72_657 ();
 sg13g2_fill_2 FILLER_72_671 ();
 sg13g2_fill_2 FILLER_72_686 ();
 sg13g2_fill_1 FILLER_72_688 ();
 sg13g2_fill_1 FILLER_72_712 ();
 sg13g2_fill_2 FILLER_72_717 ();
 sg13g2_fill_2 FILLER_72_754 ();
 sg13g2_fill_1 FILLER_72_756 ();
 sg13g2_fill_1 FILLER_72_778 ();
 sg13g2_fill_1 FILLER_72_787 ();
 sg13g2_fill_1 FILLER_72_811 ();
 sg13g2_fill_1 FILLER_72_840 ();
 sg13g2_fill_1 FILLER_72_855 ();
 sg13g2_fill_2 FILLER_72_860 ();
 sg13g2_fill_1 FILLER_73_0 ();
 sg13g2_fill_1 FILLER_73_40 ();
 sg13g2_fill_2 FILLER_73_67 ();
 sg13g2_fill_1 FILLER_73_124 ();
 sg13g2_fill_1 FILLER_73_212 ();
 sg13g2_fill_1 FILLER_73_289 ();
 sg13g2_fill_2 FILLER_73_433 ();
 sg13g2_fill_2 FILLER_73_489 ();
 sg13g2_fill_1 FILLER_73_527 ();
 sg13g2_fill_2 FILLER_73_541 ();
 sg13g2_fill_1 FILLER_73_543 ();
 sg13g2_fill_2 FILLER_73_591 ();
 sg13g2_fill_2 FILLER_73_621 ();
 sg13g2_fill_2 FILLER_73_635 ();
 sg13g2_fill_1 FILLER_73_637 ();
 sg13g2_fill_2 FILLER_73_653 ();
 sg13g2_fill_1 FILLER_73_655 ();
 sg13g2_fill_2 FILLER_73_664 ();
 sg13g2_fill_1 FILLER_73_666 ();
 sg13g2_fill_2 FILLER_73_680 ();
 sg13g2_fill_1 FILLER_73_682 ();
 sg13g2_fill_2 FILLER_73_688 ();
 sg13g2_fill_2 FILLER_73_694 ();
 sg13g2_fill_1 FILLER_73_710 ();
 sg13g2_fill_2 FILLER_73_784 ();
 sg13g2_fill_1 FILLER_73_804 ();
 sg13g2_fill_2 FILLER_73_820 ();
 sg13g2_fill_1 FILLER_73_822 ();
 sg13g2_fill_1 FILLER_73_861 ();
 sg13g2_fill_2 FILLER_74_0 ();
 sg13g2_fill_1 FILLER_74_77 ();
 sg13g2_fill_2 FILLER_74_121 ();
 sg13g2_fill_1 FILLER_74_139 ();
 sg13g2_fill_1 FILLER_74_184 ();
 sg13g2_fill_2 FILLER_74_211 ();
 sg13g2_fill_1 FILLER_74_237 ();
 sg13g2_fill_1 FILLER_74_293 ();
 sg13g2_fill_1 FILLER_74_385 ();
 sg13g2_fill_2 FILLER_74_408 ();
 sg13g2_fill_2 FILLER_74_595 ();
 sg13g2_fill_2 FILLER_74_611 ();
 sg13g2_fill_1 FILLER_74_626 ();
 sg13g2_fill_1 FILLER_74_648 ();
 sg13g2_fill_1 FILLER_74_673 ();
 sg13g2_fill_1 FILLER_74_705 ();
 sg13g2_fill_1 FILLER_74_716 ();
 sg13g2_fill_2 FILLER_74_729 ();
 sg13g2_fill_2 FILLER_74_789 ();
 sg13g2_fill_1 FILLER_74_791 ();
 sg13g2_fill_2 FILLER_74_834 ();
 sg13g2_fill_1 FILLER_74_836 ();
 sg13g2_fill_1 FILLER_74_861 ();
 sg13g2_fill_2 FILLER_75_120 ();
 sg13g2_fill_2 FILLER_75_146 ();
 sg13g2_fill_1 FILLER_75_172 ();
 sg13g2_fill_1 FILLER_75_218 ();
 sg13g2_fill_2 FILLER_75_295 ();
 sg13g2_fill_1 FILLER_75_421 ();
 sg13g2_fill_2 FILLER_75_541 ();
 sg13g2_fill_1 FILLER_75_543 ();
 sg13g2_fill_2 FILLER_75_584 ();
 sg13g2_fill_2 FILLER_75_627 ();
 sg13g2_fill_1 FILLER_75_629 ();
 sg13g2_fill_2 FILLER_75_655 ();
 sg13g2_fill_2 FILLER_75_677 ();
 sg13g2_fill_1 FILLER_75_679 ();
 sg13g2_fill_1 FILLER_75_687 ();
 sg13g2_fill_2 FILLER_75_700 ();
 sg13g2_fill_1 FILLER_75_702 ();
 sg13g2_fill_1 FILLER_75_711 ();
 sg13g2_fill_2 FILLER_75_717 ();
 sg13g2_fill_1 FILLER_75_744 ();
 sg13g2_fill_2 FILLER_75_754 ();
 sg13g2_fill_1 FILLER_75_812 ();
 sg13g2_fill_1 FILLER_75_830 ();
 sg13g2_fill_2 FILLER_75_860 ();
 sg13g2_fill_2 FILLER_76_46 ();
 sg13g2_fill_2 FILLER_76_213 ();
 sg13g2_fill_2 FILLER_76_258 ();
 sg13g2_fill_2 FILLER_76_285 ();
 sg13g2_fill_2 FILLER_76_363 ();
 sg13g2_fill_2 FILLER_76_459 ();
 sg13g2_fill_2 FILLER_76_529 ();
 sg13g2_fill_1 FILLER_76_562 ();
 sg13g2_fill_2 FILLER_76_579 ();
 sg13g2_fill_2 FILLER_76_592 ();
 sg13g2_fill_2 FILLER_76_601 ();
 sg13g2_fill_1 FILLER_76_603 ();
 sg13g2_fill_1 FILLER_76_628 ();
 sg13g2_fill_1 FILLER_76_646 ();
 sg13g2_fill_2 FILLER_76_676 ();
 sg13g2_fill_2 FILLER_76_699 ();
 sg13g2_fill_1 FILLER_76_705 ();
 sg13g2_fill_2 FILLER_76_753 ();
 sg13g2_fill_2 FILLER_76_767 ();
 sg13g2_fill_1 FILLER_76_769 ();
 sg13g2_fill_2 FILLER_76_775 ();
 sg13g2_fill_2 FILLER_76_793 ();
 sg13g2_fill_1 FILLER_76_809 ();
 sg13g2_fill_2 FILLER_76_859 ();
 sg13g2_fill_1 FILLER_76_861 ();
 sg13g2_fill_2 FILLER_77_105 ();
 sg13g2_fill_1 FILLER_77_135 ();
 sg13g2_fill_2 FILLER_77_150 ();
 sg13g2_fill_2 FILLER_77_314 ();
 sg13g2_fill_2 FILLER_77_344 ();
 sg13g2_fill_1 FILLER_77_383 ();
 sg13g2_fill_2 FILLER_77_523 ();
 sg13g2_fill_1 FILLER_77_525 ();
 sg13g2_fill_2 FILLER_77_534 ();
 sg13g2_fill_1 FILLER_77_554 ();
 sg13g2_fill_2 FILLER_77_594 ();
 sg13g2_fill_1 FILLER_77_596 ();
 sg13g2_fill_1 FILLER_77_636 ();
 sg13g2_fill_2 FILLER_77_653 ();
 sg13g2_fill_1 FILLER_77_680 ();
 sg13g2_fill_2 FILLER_77_709 ();
 sg13g2_fill_1 FILLER_77_711 ();
 sg13g2_fill_1 FILLER_77_724 ();
 sg13g2_fill_2 FILLER_77_754 ();
 sg13g2_fill_2 FILLER_77_797 ();
 sg13g2_fill_1 FILLER_77_812 ();
 sg13g2_fill_1 FILLER_77_818 ();
 sg13g2_fill_2 FILLER_77_830 ();
 sg13g2_fill_1 FILLER_77_832 ();
 sg13g2_fill_1 FILLER_77_839 ();
 sg13g2_fill_2 FILLER_77_860 ();
 sg13g2_fill_1 FILLER_78_0 ();
 sg13g2_fill_1 FILLER_78_95 ();
 sg13g2_fill_1 FILLER_78_129 ();
 sg13g2_fill_1 FILLER_78_222 ();
 sg13g2_fill_2 FILLER_78_341 ();
 sg13g2_fill_2 FILLER_78_459 ();
 sg13g2_fill_2 FILLER_78_533 ();
 sg13g2_fill_2 FILLER_78_579 ();
 sg13g2_fill_2 FILLER_78_598 ();
 sg13g2_fill_2 FILLER_78_605 ();
 sg13g2_fill_2 FILLER_78_614 ();
 sg13g2_fill_1 FILLER_78_623 ();
 sg13g2_fill_2 FILLER_78_630 ();
 sg13g2_fill_1 FILLER_78_632 ();
 sg13g2_fill_1 FILLER_78_651 ();
 sg13g2_fill_2 FILLER_78_685 ();
 sg13g2_fill_2 FILLER_78_692 ();
 sg13g2_fill_1 FILLER_78_694 ();
 sg13g2_fill_1 FILLER_78_712 ();
 sg13g2_fill_2 FILLER_78_726 ();
 sg13g2_fill_1 FILLER_78_728 ();
 sg13g2_fill_1 FILLER_78_759 ();
 sg13g2_fill_1 FILLER_78_843 ();
 sg13g2_fill_1 FILLER_78_861 ();
 sg13g2_fill_2 FILLER_79_0 ();
 sg13g2_fill_1 FILLER_79_2 ();
 sg13g2_fill_2 FILLER_79_13 ();
 sg13g2_fill_2 FILLER_79_85 ();
 sg13g2_fill_1 FILLER_79_216 ();
 sg13g2_fill_2 FILLER_79_280 ();
 sg13g2_fill_2 FILLER_79_551 ();
 sg13g2_fill_2 FILLER_79_560 ();
 sg13g2_fill_1 FILLER_79_562 ();
 sg13g2_fill_2 FILLER_79_581 ();
 sg13g2_fill_1 FILLER_79_619 ();
 sg13g2_fill_2 FILLER_79_648 ();
 sg13g2_fill_1 FILLER_79_650 ();
 sg13g2_fill_2 FILLER_79_658 ();
 sg13g2_fill_1 FILLER_79_660 ();
 sg13g2_fill_1 FILLER_79_676 ();
 sg13g2_fill_1 FILLER_79_697 ();
 sg13g2_fill_2 FILLER_79_719 ();
 sg13g2_fill_1 FILLER_79_745 ();
 sg13g2_fill_2 FILLER_79_761 ();
 sg13g2_fill_2 FILLER_79_795 ();
 sg13g2_fill_1 FILLER_79_797 ();
 sg13g2_fill_2 FILLER_80_15 ();
 sg13g2_fill_1 FILLER_80_119 ();
 sg13g2_fill_2 FILLER_80_184 ();
 sg13g2_fill_1 FILLER_80_215 ();
 sg13g2_fill_2 FILLER_80_261 ();
 sg13g2_fill_2 FILLER_80_421 ();
 sg13g2_fill_1 FILLER_80_510 ();
 sg13g2_fill_1 FILLER_80_583 ();
 sg13g2_fill_2 FILLER_80_602 ();
 sg13g2_fill_1 FILLER_80_604 ();
 sg13g2_fill_2 FILLER_80_614 ();
 sg13g2_fill_1 FILLER_80_616 ();
 sg13g2_fill_2 FILLER_80_622 ();
 sg13g2_fill_2 FILLER_80_633 ();
 sg13g2_fill_1 FILLER_80_635 ();
 sg13g2_fill_1 FILLER_80_649 ();
 sg13g2_fill_2 FILLER_80_662 ();
 sg13g2_fill_2 FILLER_80_690 ();
 sg13g2_fill_1 FILLER_80_692 ();
 sg13g2_fill_1 FILLER_80_730 ();
 sg13g2_fill_2 FILLER_80_749 ();
 sg13g2_fill_1 FILLER_80_751 ();
 sg13g2_fill_2 FILLER_80_757 ();
 sg13g2_fill_1 FILLER_80_759 ();
 sg13g2_fill_2 FILLER_80_777 ();
 sg13g2_fill_2 FILLER_80_791 ();
 sg13g2_fill_1 FILLER_80_805 ();
 sg13g2_fill_1 FILLER_80_840 ();
 sg13g2_fill_2 FILLER_80_860 ();
 assign uio_oe[0] = net11;
 assign uio_oe[1] = net12;
 assign uio_oe[2] = net13;
 assign uio_oe[3] = net14;
 assign uio_oe[4] = net15;
 assign uio_oe[5] = net16;
 assign uio_oe[6] = net17;
 assign uio_oe[7] = net18;
 assign uio_out[0] = net19;
 assign uio_out[1] = net20;
 assign uio_out[2] = net21;
 assign uio_out[3] = net22;
 assign uio_out[4] = net23;
 assign uio_out[5] = net24;
 assign uio_out[6] = net25;
 assign uio_out[7] = net26;
endmodule
