module tt_um_crockpotveggies_neuron (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _160_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _164_;
 wire _165_;
 wire _166_;
 wire _167_;
 wire _168_;
 wire _169_;
 wire _170_;
 wire _171_;
 wire _172_;
 wire _173_;
 wire _174_;
 wire _175_;
 wire _176_;
 wire _177_;
 wire _178_;
 wire _179_;
 wire _180_;
 wire _181_;
 wire _182_;
 wire _183_;
 wire _184_;
 wire _185_;
 wire _186_;
 wire _187_;
 wire _188_;
 wire _189_;
 wire _190_;
 wire _191_;
 wire _192_;
 wire _193_;
 wire _194_;
 wire _195_;
 wire _196_;
 wire _197_;
 wire _198_;
 wire _199_;
 wire _200_;
 wire _201_;
 wire _202_;
 wire _203_;
 wire _204_;
 wire _205_;
 wire _206_;
 wire _207_;
 wire _208_;
 wire _209_;
 wire _210_;
 wire _211_;
 wire _212_;
 wire _213_;
 wire _214_;
 wire _215_;
 wire _216_;
 wire _217_;
 wire _218_;
 wire _219_;
 wire _220_;
 wire _221_;
 wire _222_;
 wire _223_;
 wire _224_;
 wire _225_;
 wire _226_;
 wire _227_;
 wire _228_;
 wire _229_;
 wire _230_;
 wire _231_;
 wire _232_;
 wire _233_;
 wire _234_;
 wire _235_;
 wire _236_;
 wire _237_;
 wire _238_;
 wire _239_;
 wire _240_;
 wire _241_;
 wire _242_;
 wire _243_;
 wire _244_;
 wire _245_;
 wire _246_;
 wire _247_;
 wire \u_neuron.addr[0] ;
 wire \u_neuron.addr[1] ;
 wire \u_neuron.addr[2] ;
 wire \u_neuron.addr[3] ;
 wire \u_neuron.addr[4] ;
 wire \u_neuron.addr[5] ;
 wire \u_neuron.arm_event ;
 wire \u_neuron.cfg_arg[0] ;
 wire \u_neuron.cfg_arg[1] ;
 wire \u_neuron.cfg_arg[2] ;
 wire \u_neuron.cfg_arg[3] ;
 wire \u_neuron.cfg_op[0] ;
 wire \u_neuron.cfg_op[1] ;
 wire \u_neuron.conv_emit_data[0] ;
 wire \u_neuron.conv_emit_data[1] ;
 wire \u_neuron.conv_emit_data[2] ;
 wire net18;
 wire \u_neuron.conv_emit_data[4] ;
 wire net19;
 wire \u_neuron.conv_emit_data[6] ;
 wire net38;
 wire \u_neuron.conv_emit_valid ;
 wire \u_neuron.conv_last_sum[0] ;
 wire \u_neuron.conv_last_sum[1] ;
 wire \u_neuron.conv_last_sum[2] ;
 wire \u_neuron.conv_last_sum_next[0] ;
 wire \u_neuron.conv_last_sum_next[1] ;
 wire \u_neuron.conv_last_sum_next[2] ;
 wire net20;
 wire \u_neuron.conv_post_spike ;
 wire \u_neuron.conv_shift[0] ;
 wire \u_neuron.conv_shift[1] ;
 wire \u_neuron.conv_shift[2] ;
 wire \u_neuron.conv_shift[3] ;
 wire \u_neuron.conv_shift_next[0] ;
 wire \u_neuron.conv_shift_next[1] ;
 wire \u_neuron.conv_shift_next[2] ;
 wire \u_neuron.conv_shift_next[3] ;
 wire \u_neuron.fst_armed ;
 wire \u_neuron.fst_armed_next ;
 wire \u_neuron.fst_emit_data[0] ;
 wire \u_neuron.fst_emit_data[1] ;
 wire \u_neuron.fst_emit_data[2] ;
 wire \u_neuron.fst_emit_data[3] ;
 wire \u_neuron.fst_emit_data[4] ;
 wire net33;
 wire \u_neuron.fst_emit_data[6] ;
 wire net41;
 wire \u_neuron.fst_emit_valid ;
 wire \u_neuron.fst_last_t[0] ;
 wire \u_neuron.fst_last_t[1] ;
 wire \u_neuron.fst_last_t[2] ;
 wire \u_neuron.fst_last_t[3] ;
 wire \u_neuron.fst_last_t[4] ;
 wire \u_neuron.fst_last_t[5] ;
 wire \u_neuron.fst_last_t[6] ;
 wire \u_neuron.fst_last_t[7] ;
 wire \u_neuron.fst_last_t_next[0] ;
 wire \u_neuron.fst_last_t_next[1] ;
 wire \u_neuron.fst_last_t_next[2] ;
 wire \u_neuron.fst_last_t_next[3] ;
 wire \u_neuron.fst_last_t_next[4] ;
 wire \u_neuron.fst_last_t_next[5] ;
 wire \u_neuron.fst_last_t_next[6] ;
 wire \u_neuron.fst_last_t_next[7] ;
 wire net34;
 wire \u_neuron.fst_post_spike ;
 wire \u_neuron.fst_t[0] ;
 wire \u_neuron.fst_t[1] ;
 wire \u_neuron.fst_t[2] ;
 wire \u_neuron.fst_t[3] ;
 wire \u_neuron.fst_t[4] ;
 wire \u_neuron.fst_t[5] ;
 wire \u_neuron.fst_t[6] ;
 wire \u_neuron.fst_t[7] ;
 wire \u_neuron.fst_t_next[0] ;
 wire \u_neuron.fst_t_next[1] ;
 wire \u_neuron.fst_t_next[2] ;
 wire \u_neuron.fst_t_next[3] ;
 wire \u_neuron.fst_t_next[4] ;
 wire \u_neuron.fst_t_next[5] ;
 wire \u_neuron.fst_t_next[6] ;
 wire \u_neuron.fst_t_next[7] ;
 wire \u_neuron.have_out ;
 wire \u_neuron.in_ack ;
 wire \u_neuron.in_data[0] ;
 wire \u_neuron.in_data[1] ;
 wire \u_neuron.in_data[2] ;
 wire \u_neuron.in_data[3] ;
 wire \u_neuron.in_data[4] ;
 wire \u_neuron.in_data[5] ;
 wire \u_neuron.in_data[6] ;
 wire \u_neuron.in_data[7] ;
 wire \u_neuron.in_fire ;
 wire \u_neuron.in_req_seen ;
 wire \u_neuron.is_arm_cmd ;
 wire \u_neuron.is_cfg_cmd ;
 wire \u_neuron.is_prog_addr ;
 wire \u_neuron.is_reset_cmd ;
 wire \u_neuron.is_special_cmd ;
 wire \u_neuron.is_tick ;
 wire \u_neuron.learn_en ;
 wire \u_neuron.learn_pending ;
 wire \u_neuron.learn_ptr[0] ;
 wire \u_neuron.learn_ptr[1] ;
 wire \u_neuron.learn_ptr[2] ;
 wire \u_neuron.learn_ptr[3] ;
 wire \u_neuron.lif_V[0] ;
 wire \u_neuron.lif_V[1] ;
 wire \u_neuron.lif_V[2] ;
 wire \u_neuron.lif_V[3] ;
 wire \u_neuron.lif_V[4] ;
 wire \u_neuron.lif_V[5] ;
 wire \u_neuron.lif_V[6] ;
 wire \u_neuron.lif_V[7] ;
 wire \u_neuron.lif_V_next[0] ;
 wire \u_neuron.lif_V_next[1] ;
 wire \u_neuron.lif_V_next[2] ;
 wire \u_neuron.lif_V_next[3] ;
 wire \u_neuron.lif_V_next[4] ;
 wire \u_neuron.lif_V_next[5] ;
 wire \u_neuron.lif_V_next[6] ;
 wire \u_neuron.lif_V_next[7] ;
 wire \u_neuron.lif_emit_data[0] ;
 wire \u_neuron.lif_emit_data[1] ;
 wire \u_neuron.lif_emit_data[2] ;
 wire \u_neuron.lif_emit_data[3] ;
 wire \u_neuron.lif_emit_data[4] ;
 wire net35;
 wire \u_neuron.lif_emit_data[6] ;
 wire net42;
 wire \u_neuron.lif_emit_valid ;
 wire \u_neuron.lif_learn_start ;
 wire \u_neuron.lif_post_spike ;
 wire \u_neuron.ltd_idx[0] ;
 wire \u_neuron.ltd_idx[1] ;
 wire \u_neuron.ltd_idx[2] ;
 wire \u_neuron.ltd_idx[3] ;
 wire \u_neuron.ltd_wdata[0] ;
 wire \u_neuron.ltd_wdata[1] ;
 wire \u_neuron.ltd_we ;
 wire \u_neuron.ltp_idx[0] ;
 wire \u_neuron.ltp_idx[1] ;
 wire \u_neuron.ltp_idx[2] ;
 wire \u_neuron.ltp_idx[3] ;
 wire \u_neuron.ltp_wdata[0] ;
 wire \u_neuron.ltp_wdata[1] ;
 wire \u_neuron.ltp_we ;
 wire \u_neuron.mode[0] ;
 wire \u_neuron.mode[1] ;
 wire \u_neuron.mode_conv_evt ;
 wire \u_neuron.mode_emit_data[0] ;
 wire \u_neuron.mode_emit_data[1] ;
 wire \u_neuron.mode_emit_data[2] ;
 wire \u_neuron.mode_emit_data[3] ;
 wire \u_neuron.mode_emit_data[4] ;
 wire \u_neuron.mode_emit_data[5] ;
 wire \u_neuron.mode_emit_data[6] ;
 wire \u_neuron.mode_emit_data[7] ;
 wire \u_neuron.mode_emit_valid ;
 wire \u_neuron.mode_fst_evt ;
 wire \u_neuron.mode_learn_start ;
 wire \u_neuron.mode_lif_evt ;
 wire \u_neuron.mode_post_spike ;
 wire \u_neuron.mode_td_evt ;
 wire \u_neuron.normal_event ;
 wire \u_neuron.out_fire ;
 wire \u_neuron.out_req ;
 wire \u_neuron.pending_widx[0] ;
 wire \u_neuron.pending_widx[1] ;
 wire \u_neuron.pending_widx[2] ;
 wire \u_neuron.pending_widx[3] ;
 wire \u_neuron.polarity ;
 wire \u_neuron.post_trace ;
 wire \u_neuron.pre_trace[0] ;
 wire \u_neuron.pre_trace[10] ;
 wire \u_neuron.pre_trace[11] ;
 wire \u_neuron.pre_trace[12] ;
 wire \u_neuron.pre_trace[13] ;
 wire \u_neuron.pre_trace[14] ;
 wire \u_neuron.pre_trace[15] ;
 wire \u_neuron.pre_trace[1] ;
 wire \u_neuron.pre_trace[2] ;
 wire \u_neuron.pre_trace[3] ;
 wire \u_neuron.pre_trace[4] ;
 wire \u_neuron.pre_trace[5] ;
 wire \u_neuron.pre_trace[6] ;
 wire \u_neuron.pre_trace[7] ;
 wire \u_neuron.pre_trace[8] ;
 wire \u_neuron.pre_trace[9] ;
 wire \u_neuron.soft_reset_fire ;
 wire \u_neuron.spike_seen_this_tick ;
 wire \u_neuron.spike_seen_this_tick_next ;
 wire \u_neuron.stream_act ;
 wire \u_neuron.td_curr[0] ;
 wire \u_neuron.td_curr[1] ;
 wire \u_neuron.td_curr[2] ;
 wire \u_neuron.td_curr[3] ;
 wire \u_neuron.td_curr[4] ;
 wire \u_neuron.td_curr[5] ;
 wire \u_neuron.td_curr[6] ;
 wire \u_neuron.td_curr[7] ;
 wire \u_neuron.td_curr_next[0] ;
 wire \u_neuron.td_curr_next[1] ;
 wire \u_neuron.td_curr_next[2] ;
 wire \u_neuron.td_curr_next[3] ;
 wire \u_neuron.td_curr_next[4] ;
 wire \u_neuron.td_curr_next[5] ;
 wire \u_neuron.td_curr_next[6] ;
 wire \u_neuron.td_curr_next[7] ;
 wire \u_neuron.td_emit_data[0] ;
 wire \u_neuron.td_emit_data[1] ;
 wire \u_neuron.td_emit_data[2] ;
 wire \u_neuron.td_emit_data[3] ;
 wire \u_neuron.td_emit_data[4] ;
 wire net36;
 wire \u_neuron.td_emit_data[6] ;
 wire clknet_0_clk;
 wire \u_neuron.td_emit_valid ;
 wire \u_neuron.td_last_diff[0] ;
 wire \u_neuron.td_last_diff[1] ;
 wire \u_neuron.td_last_diff[2] ;
 wire \u_neuron.td_last_diff[3] ;
 wire \u_neuron.td_last_diff[4] ;
 wire \u_neuron.td_last_diff[5] ;
 wire \u_neuron.td_last_diff[6] ;
 wire \u_neuron.td_last_diff[7] ;
 wire \u_neuron.td_last_diff_next[0] ;
 wire \u_neuron.td_last_diff_next[1] ;
 wire \u_neuron.td_last_diff_next[2] ;
 wire \u_neuron.td_last_diff_next[3] ;
 wire \u_neuron.td_last_diff_next[4] ;
 wire \u_neuron.td_last_diff_next[5] ;
 wire \u_neuron.td_last_diff_next[6] ;
 wire \u_neuron.td_last_diff_next[7] ;
 wire net37;
 wire \u_neuron.td_post_spike ;
 wire \u_neuron.td_prev[0] ;
 wire \u_neuron.td_prev[1] ;
 wire \u_neuron.td_prev[2] ;
 wire \u_neuron.td_prev[3] ;
 wire \u_neuron.td_prev[4] ;
 wire \u_neuron.td_prev[5] ;
 wire \u_neuron.td_prev[6] ;
 wire \u_neuron.td_prev[7] ;
 wire \u_neuron.td_prev_next[0] ;
 wire \u_neuron.td_prev_next[1] ;
 wire \u_neuron.td_prev_next[2] ;
 wire \u_neuron.td_prev_next[3] ;
 wire \u_neuron.td_prev_next[4] ;
 wire \u_neuron.td_prev_next[5] ;
 wire \u_neuron.td_prev_next[6] ;
 wire \u_neuron.td_prev_next[7] ;
 wire \u_neuron.uio_in_sync[0] ;
 wire \u_neuron.uio_in_sync[1] ;
 wire \u_neuron.uio_in_sync[2] ;
 wire \u_neuron.uio_in_sync[3] ;
 wire \u_neuron.uio_in_sync[4] ;
 wire \u_neuron.uio_in_sync[5] ;
 wire \u_neuron.uio_in_sync[6] ;
 wire \u_neuron.uio_in_sync[7] ;
 wire \u_neuron.w_addr_curr[0] ;
 wire \u_neuron.w_addr_curr[1] ;
 wire \u_neuron.w_eff[0] ;
 wire \u_neuron.w_eff[1] ;
 wire \u_neuron.w_ptr_curr[0] ;
 wire \u_neuron.w_ptr_curr[1] ;
 wire \u_neuron.wtab[0] ;
 wire \u_neuron.wtab[10] ;
 wire \u_neuron.wtab[11] ;
 wire \u_neuron.wtab[12] ;
 wire \u_neuron.wtab[13] ;
 wire \u_neuron.wtab[14] ;
 wire \u_neuron.wtab[15] ;
 wire \u_neuron.wtab[16] ;
 wire \u_neuron.wtab[17] ;
 wire \u_neuron.wtab[18] ;
 wire \u_neuron.wtab[19] ;
 wire \u_neuron.wtab[1] ;
 wire \u_neuron.wtab[20] ;
 wire \u_neuron.wtab[21] ;
 wire \u_neuron.wtab[22] ;
 wire \u_neuron.wtab[23] ;
 wire \u_neuron.wtab[24] ;
 wire \u_neuron.wtab[25] ;
 wire \u_neuron.wtab[26] ;
 wire \u_neuron.wtab[27] ;
 wire \u_neuron.wtab[28] ;
 wire \u_neuron.wtab[29] ;
 wire \u_neuron.wtab[2] ;
 wire \u_neuron.wtab[30] ;
 wire \u_neuron.wtab[31] ;
 wire \u_neuron.wtab[3] ;
 wire \u_neuron.wtab[4] ;
 wire \u_neuron.wtab[5] ;
 wire \u_neuron.wtab[6] ;
 wire \u_neuron.wtab[7] ;
 wire \u_neuron.wtab[8] ;
 wire \u_neuron.wtab[9] ;
 wire net39;
 wire net40;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire \u_neuron.u_conv/_00_ ;
 wire \u_neuron.u_conv/_01_ ;
 wire \u_neuron.u_conv/_02_ ;
 wire \u_neuron.u_conv/_03_ ;
 wire \u_neuron.u_conv/_04_ ;
 wire \u_neuron.u_conv/_05_ ;
 wire \u_neuron.u_conv/_06_ ;
 wire \u_neuron.u_conv/_07_ ;
 wire \u_neuron.u_decode/_00_ ;
 wire \u_neuron.u_decode/_01_ ;
 wire \u_neuron.u_decode/_02_ ;
 wire \u_neuron.u_decode/_03_ ;
 wire \u_neuron.u_frontend/_00_ ;
 wire \u_neuron.u_frontend/_01_ ;
 wire \u_neuron.u_frontend/_02_ ;
 wire \u_neuron.u_frontend/_03_ ;
 wire \u_neuron.u_frontend/in_req ;
 wire \u_neuron.u_frontend/out_ack ;
 wire \u_neuron.u_frontend/ui_in_meta[0] ;
 wire \u_neuron.u_frontend/ui_in_meta[1] ;
 wire \u_neuron.u_frontend/ui_in_meta[2] ;
 wire \u_neuron.u_frontend/ui_in_meta[3] ;
 wire \u_neuron.u_frontend/ui_in_meta[4] ;
 wire \u_neuron.u_frontend/ui_in_meta[5] ;
 wire \u_neuron.u_frontend/ui_in_meta[6] ;
 wire \u_neuron.u_frontend/ui_in_meta[7] ;
 wire \u_neuron.u_frontend/uio_in_meta[0] ;
 wire \u_neuron.u_frontend/uio_in_meta[1] ;
 wire \u_neuron.u_frontend/uio_in_meta[2] ;
 wire \u_neuron.u_frontend/uio_in_meta[3] ;
 wire \u_neuron.u_frontend/uio_in_meta[4] ;
 wire \u_neuron.u_frontend/uio_in_meta[5] ;
 wire \u_neuron.u_frontend/uio_in_meta[6] ;
 wire \u_neuron.u_frontend/uio_in_meta[7] ;
 wire \u_neuron.u_fst/_000_ ;
 wire \u_neuron.u_fst/_001_ ;
 wire \u_neuron.u_fst/_002_ ;
 wire \u_neuron.u_fst/_003_ ;
 wire \u_neuron.u_fst/_004_ ;
 wire \u_neuron.u_fst/_005_ ;
 wire \u_neuron.u_fst/_006_ ;
 wire \u_neuron.u_fst/_007_ ;
 wire \u_neuron.u_fst/_008_ ;
 wire \u_neuron.u_fst/_009_ ;
 wire \u_neuron.u_fst/_010_ ;
 wire \u_neuron.u_fst/_011_ ;
 wire \u_neuron.u_fst/_012_ ;
 wire \u_neuron.u_fst/_013_ ;
 wire \u_neuron.u_fst/_014_ ;
 wire \u_neuron.u_fst/_015_ ;
 wire \u_neuron.u_fst/_016_ ;
 wire \u_neuron.u_fst/_017_ ;
 wire \u_neuron.u_fst/_018_ ;
 wire \u_neuron.u_fst/_019_ ;
 wire \u_neuron.u_fst/_020_ ;
 wire \u_neuron.u_fst/_021_ ;
 wire \u_neuron.u_fst/_022_ ;
 wire \u_neuron.u_fst/_023_ ;
 wire \u_neuron.u_fst/_024_ ;
 wire \u_neuron.u_fst/_025_ ;
 wire \u_neuron.u_fst/_026_ ;
 wire \u_neuron.u_fst/_027_ ;
 wire \u_neuron.u_fst/_028_ ;
 wire \u_neuron.u_fst/_029_ ;
 wire \u_neuron.u_fst/_030_ ;
 wire \u_neuron.u_fst/_031_ ;
 wire \u_neuron.u_fst/_032_ ;
 wire \u_neuron.u_fst/_033_ ;
 wire \u_neuron.u_fst/_034_ ;
 wire \u_neuron.u_fst/_035_ ;
 wire \u_neuron.u_fst/_036_ ;
 wire \u_neuron.u_fst/_037_ ;
 wire \u_neuron.u_fst/_038_ ;
 wire \u_neuron.u_fst/_039_ ;
 wire \u_neuron.u_fst/_040_ ;
 wire \u_neuron.u_fst/_041_ ;
 wire \u_neuron.u_fst/_042_ ;
 wire \u_neuron.u_fst/_043_ ;
 wire \u_neuron.u_fst/_044_ ;
 wire \u_neuron.u_fst/_045_ ;
 wire \u_neuron.u_fst/_046_ ;
 wire \u_neuron.u_fst/_047_ ;
 wire \u_neuron.u_learning/_000_ ;
 wire \u_neuron.u_learning/_001_ ;
 wire \u_neuron.u_learning/_002_ ;
 wire \u_neuron.u_learning/_003_ ;
 wire \u_neuron.u_learning/_004_ ;
 wire \u_neuron.u_learning/_005_ ;
 wire \u_neuron.u_learning/_006_ ;
 wire \u_neuron.u_learning/_007_ ;
 wire \u_neuron.u_learning/_008_ ;
 wire \u_neuron.u_learning/_009_ ;
 wire \u_neuron.u_learning/_010_ ;
 wire \u_neuron.u_learning/_011_ ;
 wire \u_neuron.u_learning/_012_ ;
 wire \u_neuron.u_learning/_013_ ;
 wire \u_neuron.u_learning/_014_ ;
 wire \u_neuron.u_learning/_015_ ;
 wire \u_neuron.u_learning/_016_ ;
 wire \u_neuron.u_learning/_017_ ;
 wire \u_neuron.u_learning/_018_ ;
 wire \u_neuron.u_learning/_019_ ;
 wire \u_neuron.u_learning/_020_ ;
 wire \u_neuron.u_learning/_021_ ;
 wire \u_neuron.u_learning/_022_ ;
 wire \u_neuron.u_learning/_023_ ;
 wire \u_neuron.u_learning/_024_ ;
 wire \u_neuron.u_learning/_025_ ;
 wire \u_neuron.u_learning/_026_ ;
 wire \u_neuron.u_learning/_027_ ;
 wire \u_neuron.u_learning/_028_ ;
 wire \u_neuron.u_learning/_029_ ;
 wire \u_neuron.u_learning/_030_ ;
 wire \u_neuron.u_learning/_031_ ;
 wire \u_neuron.u_learning/_032_ ;
 wire \u_neuron.u_learning/_033_ ;
 wire \u_neuron.u_learning/_034_ ;
 wire \u_neuron.u_learning/_035_ ;
 wire \u_neuron.u_learning/_036_ ;
 wire \u_neuron.u_learning/_037_ ;
 wire \u_neuron.u_learning/_038_ ;
 wire \u_neuron.u_learning/_039_ ;
 wire \u_neuron.u_learning/_040_ ;
 wire \u_neuron.u_learning/_041_ ;
 wire \u_neuron.u_learning/_042_ ;
 wire \u_neuron.u_learning/_043_ ;
 wire \u_neuron.u_learning/_044_ ;
 wire \u_neuron.u_learning/_045_ ;
 wire \u_neuron.u_learning/_046_ ;
 wire \u_neuron.u_learning/_047_ ;
 wire \u_neuron.u_learning/_048_ ;
 wire \u_neuron.u_learning/_049_ ;
 wire \u_neuron.u_learning/_050_ ;
 wire \u_neuron.u_learning/_051_ ;
 wire \u_neuron.u_learning/_052_ ;
 wire \u_neuron.u_learning/_053_ ;
 wire \u_neuron.u_learning/_054_ ;
 wire \u_neuron.u_learning/_055_ ;
 wire \u_neuron.u_learning/_056_ ;
 wire \u_neuron.u_learning/_057_ ;
 wire \u_neuron.u_learning/_058_ ;
 wire \u_neuron.u_learning/_059_ ;
 wire \u_neuron.u_learning/_060_ ;
 wire \u_neuron.u_learning/_061_ ;
 wire \u_neuron.u_learning/_062_ ;
 wire \u_neuron.u_learning/_063_ ;
 wire \u_neuron.u_learning/_064_ ;
 wire \u_neuron.u_learning/_065_ ;
 wire \u_neuron.u_learning/_066_ ;
 wire \u_neuron.u_learning/_067_ ;
 wire \u_neuron.u_learning/_068_ ;
 wire \u_neuron.u_learning/_069_ ;
 wire \u_neuron.u_learning/_070_ ;
 wire \u_neuron.u_learning/_071_ ;
 wire \u_neuron.u_learning/_072_ ;
 wire \u_neuron.u_learning/_073_ ;
 wire \u_neuron.u_learning/_074_ ;
 wire \u_neuron.u_learning/_075_ ;
 wire \u_neuron.u_learning/_076_ ;
 wire \u_neuron.u_learning/_077_ ;
 wire \u_neuron.u_learning/_078_ ;
 wire \u_neuron.u_learning/_079_ ;
 wire \u_neuron.u_learning/_080_ ;
 wire \u_neuron.u_learning/_081_ ;
 wire \u_neuron.u_learning/_082_ ;
 wire \u_neuron.u_learning/_083_ ;
 wire \u_neuron.u_learning/_084_ ;
 wire \u_neuron.u_learning/_085_ ;
 wire \u_neuron.u_learning/_086_ ;
 wire \u_neuron.u_learning/_087_ ;
 wire \u_neuron.u_learning/_088_ ;
 wire \u_neuron.u_learning/_089_ ;
 wire \u_neuron.u_learning/_090_ ;
 wire \u_neuron.u_learning/_091_ ;
 wire \u_neuron.u_learning/_092_ ;
 wire \u_neuron.u_learning/_093_ ;
 wire \u_neuron.u_learning/_094_ ;
 wire \u_neuron.u_learning/_095_ ;
 wire \u_neuron.u_learning/_096_ ;
 wire \u_neuron.u_learning/_097_ ;
 wire \u_neuron.u_learning/_098_ ;
 wire \u_neuron.u_learning/_099_ ;
 wire \u_neuron.u_learning/_100_ ;
 wire \u_neuron.u_learning/_101_ ;
 wire \u_neuron.u_learning/_102_ ;
 wire \u_neuron.u_learning/_103_ ;
 wire \u_neuron.u_learning/_104_ ;
 wire \u_neuron.u_learning/_105_ ;
 wire \u_neuron.u_learning/_106_ ;
 wire \u_neuron.u_learning/_107_ ;
 wire \u_neuron.u_learning/_108_ ;
 wire \u_neuron.u_learning/_109_ ;
 wire \u_neuron.u_learning/_110_ ;
 wire \u_neuron.u_learning/_111_ ;
 wire \u_neuron.u_learning/_112_ ;
 wire \u_neuron.u_learning/_113_ ;
 wire \u_neuron.u_learning/_114_ ;
 wire \u_neuron.u_learning/_115_ ;
 wire \u_neuron.u_learning/_116_ ;
 wire \u_neuron.u_learning/_117_ ;
 wire \u_neuron.u_learning/_118_ ;
 wire \u_neuron.u_learning/_119_ ;
 wire \u_neuron.u_learning/_120_ ;
 wire \u_neuron.u_learning/_121_ ;
 wire \u_neuron.u_learning/_122_ ;
 wire \u_neuron.u_learning/_123_ ;
 wire \u_neuron.u_learning/_124_ ;
 wire \u_neuron.u_learning/_125_ ;
 wire \u_neuron.u_learning/_126_ ;
 wire \u_neuron.u_learning/_127_ ;
 wire \u_neuron.u_learning/_128_ ;
 wire \u_neuron.u_learning/_129_ ;
 wire \u_neuron.u_learning/_130_ ;
 wire \u_neuron.u_learning/_131_ ;
 wire \u_neuron.u_learning/_132_ ;
 wire \u_neuron.u_learning/_133_ ;
 wire \u_neuron.u_learning/_134_ ;
 wire \u_neuron.u_learning/_135_ ;
 wire \u_neuron.u_learning/_136_ ;
 wire \u_neuron.u_learning/_137_ ;
 wire \u_neuron.u_learning/_138_ ;
 wire \u_neuron.u_learning/_139_ ;
 wire \u_neuron.u_learning/_140_ ;
 wire \u_neuron.u_learning/_141_ ;
 wire \u_neuron.u_learning/_142_ ;
 wire \u_neuron.u_learning/_143_ ;
 wire \u_neuron.u_learning/_144_ ;
 wire \u_neuron.u_learning/_145_ ;
 wire \u_neuron.u_learning/_146_ ;
 wire \u_neuron.u_learning/_147_ ;
 wire \u_neuron.u_learning/_148_ ;
 wire \u_neuron.u_learning/_149_ ;
 wire \u_neuron.u_learning/_150_ ;
 wire \u_neuron.u_lif/_000_ ;
 wire \u_neuron.u_lif/_001_ ;
 wire \u_neuron.u_lif/_002_ ;
 wire \u_neuron.u_lif/_003_ ;
 wire \u_neuron.u_lif/_004_ ;
 wire \u_neuron.u_lif/_005_ ;
 wire \u_neuron.u_lif/_006_ ;
 wire \u_neuron.u_lif/_007_ ;
 wire \u_neuron.u_lif/_008_ ;
 wire \u_neuron.u_lif/_009_ ;
 wire \u_neuron.u_lif/_010_ ;
 wire \u_neuron.u_lif/_011_ ;
 wire \u_neuron.u_lif/_012_ ;
 wire \u_neuron.u_lif/_013_ ;
 wire \u_neuron.u_lif/_014_ ;
 wire \u_neuron.u_lif/_015_ ;
 wire \u_neuron.u_lif/_016_ ;
 wire \u_neuron.u_lif/_017_ ;
 wire \u_neuron.u_lif/_018_ ;
 wire \u_neuron.u_lif/_019_ ;
 wire \u_neuron.u_lif/_020_ ;
 wire \u_neuron.u_lif/_021_ ;
 wire \u_neuron.u_lif/_022_ ;
 wire \u_neuron.u_lif/_023_ ;
 wire \u_neuron.u_lif/_024_ ;
 wire \u_neuron.u_lif/_025_ ;
 wire \u_neuron.u_lif/_026_ ;
 wire \u_neuron.u_lif/_027_ ;
 wire \u_neuron.u_lif/_028_ ;
 wire \u_neuron.u_lif/_029_ ;
 wire \u_neuron.u_lif/_030_ ;
 wire \u_neuron.u_lif/_031_ ;
 wire \u_neuron.u_lif/_032_ ;
 wire \u_neuron.u_lif/_033_ ;
 wire \u_neuron.u_lif/_034_ ;
 wire \u_neuron.u_lif/_035_ ;
 wire \u_neuron.u_lif/_036_ ;
 wire \u_neuron.u_lif/_037_ ;
 wire \u_neuron.u_lif/_038_ ;
 wire \u_neuron.u_lif/_039_ ;
 wire \u_neuron.u_lif/_040_ ;
 wire \u_neuron.u_lif/_041_ ;
 wire \u_neuron.u_lif/_042_ ;
 wire \u_neuron.u_lif/_043_ ;
 wire \u_neuron.u_lif/_044_ ;
 wire \u_neuron.u_lif/_045_ ;
 wire \u_neuron.u_lif/_046_ ;
 wire \u_neuron.u_lif/_047_ ;
 wire \u_neuron.u_lif/_048_ ;
 wire \u_neuron.u_lif/_049_ ;
 wire \u_neuron.u_lif/_050_ ;
 wire \u_neuron.u_lif/_051_ ;
 wire \u_neuron.u_lif/_052_ ;
 wire \u_neuron.u_lif/_053_ ;
 wire \u_neuron.u_lif/_054_ ;
 wire \u_neuron.u_lif/_055_ ;
 wire \u_neuron.u_lif/_056_ ;
 wire \u_neuron.u_lif/_057_ ;
 wire \u_neuron.u_lif/_058_ ;
 wire \u_neuron.u_lif/_059_ ;
 wire \u_neuron.u_lif/_060_ ;
 wire \u_neuron.u_outq/_00_ ;
 wire \u_neuron.u_outq/_01_ ;
 wire \u_neuron.u_outq/_02_ ;
 wire \u_neuron.u_outq/_03_ ;
 wire \u_neuron.u_outq/_04_ ;
 wire \u_neuron.u_outq/_05_ ;
 wire \u_neuron.u_outq/_06_ ;
 wire \u_neuron.u_outq/_07_ ;
 wire \u_neuron.u_outq/_08_ ;
 wire \u_neuron.u_outq/_09_ ;
 wire \u_neuron.u_outq/_10_ ;
 wire \u_neuron.u_outq/_11_ ;
 wire \u_neuron.u_outq/_12_ ;
 wire \u_neuron.u_outq/_13_ ;
 wire \u_neuron.u_outq/_14_ ;
 wire \u_neuron.u_outq/_15_ ;
 wire \u_neuron.u_outq/_16_ ;
 wire \u_neuron.u_outq/_17_ ;
 wire \u_neuron.u_outq/_18_ ;
 wire \u_neuron.u_outq/_19_ ;
 wire \u_neuron.u_outq/_20_ ;
 wire \u_neuron.u_outq/_21_ ;
 wire \u_neuron.u_outq/_22_ ;
 wire \u_neuron.u_outq/_23_ ;
 wire \u_neuron.u_outq/_24_ ;
 wire \u_neuron.u_outq/_25_ ;
 wire \u_neuron.u_outq/_26_ ;
 wire \u_neuron.u_outq/_27_ ;
 wire \u_neuron.u_outq/_28_ ;
 wire \u_neuron.u_syn/_000_ ;
 wire \u_neuron.u_syn/_001_ ;
 wire \u_neuron.u_syn/_002_ ;
 wire \u_neuron.u_syn/_003_ ;
 wire \u_neuron.u_syn/_004_ ;
 wire \u_neuron.u_syn/_005_ ;
 wire \u_neuron.u_syn/_006_ ;
 wire \u_neuron.u_syn/_007_ ;
 wire \u_neuron.u_syn/_008_ ;
 wire \u_neuron.u_syn/_009_ ;
 wire \u_neuron.u_syn/_010_ ;
 wire \u_neuron.u_syn/_011_ ;
 wire \u_neuron.u_syn/_012_ ;
 wire \u_neuron.u_syn/_013_ ;
 wire \u_neuron.u_syn/_014_ ;
 wire \u_neuron.u_syn/_015_ ;
 wire \u_neuron.u_syn/_016_ ;
 wire \u_neuron.u_syn/_017_ ;
 wire \u_neuron.u_syn/_018_ ;
 wire \u_neuron.u_syn/_019_ ;
 wire \u_neuron.u_syn/_020_ ;
 wire \u_neuron.u_syn/_021_ ;
 wire \u_neuron.u_syn/_022_ ;
 wire \u_neuron.u_syn/_023_ ;
 wire \u_neuron.u_syn/_024_ ;
 wire \u_neuron.u_syn/_025_ ;
 wire \u_neuron.u_syn/_026_ ;
 wire \u_neuron.u_syn/_027_ ;
 wire \u_neuron.u_syn/_028_ ;
 wire \u_neuron.u_syn/_029_ ;
 wire \u_neuron.u_syn/_030_ ;
 wire \u_neuron.u_syn/_031_ ;
 wire \u_neuron.u_syn/_032_ ;
 wire \u_neuron.u_syn/_033_ ;
 wire \u_neuron.u_syn/_034_ ;
 wire \u_neuron.u_syn/_035_ ;
 wire \u_neuron.u_syn/_036_ ;
 wire \u_neuron.u_syn/_037_ ;
 wire \u_neuron.u_syn/_038_ ;
 wire \u_neuron.u_syn/_039_ ;
 wire \u_neuron.u_syn/_040_ ;
 wire \u_neuron.u_syn/_041_ ;
 wire \u_neuron.u_syn/_042_ ;
 wire \u_neuron.u_syn/_043_ ;
 wire \u_neuron.u_syn/_044_ ;
 wire \u_neuron.u_syn/_045_ ;
 wire \u_neuron.u_syn/_046_ ;
 wire \u_neuron.u_syn/_047_ ;
 wire \u_neuron.u_syn/_048_ ;
 wire \u_neuron.u_syn/_049_ ;
 wire \u_neuron.u_syn/_050_ ;
 wire \u_neuron.u_syn/_051_ ;
 wire \u_neuron.u_syn/_052_ ;
 wire \u_neuron.u_syn/_053_ ;
 wire \u_neuron.u_syn/_054_ ;
 wire \u_neuron.u_syn/_055_ ;
 wire \u_neuron.u_syn/_056_ ;
 wire \u_neuron.u_syn/_057_ ;
 wire \u_neuron.u_syn/_058_ ;
 wire \u_neuron.u_syn/_059_ ;
 wire \u_neuron.u_syn/_060_ ;
 wire \u_neuron.u_syn/_061_ ;
 wire \u_neuron.u_syn/_062_ ;
 wire \u_neuron.u_syn/_063_ ;
 wire \u_neuron.u_syn/_064_ ;
 wire \u_neuron.u_syn/_065_ ;
 wire \u_neuron.u_syn/_066_ ;
 wire \u_neuron.u_syn/_067_ ;
 wire \u_neuron.u_syn/_068_ ;
 wire \u_neuron.u_syn/_069_ ;
 wire \u_neuron.u_syn/_070_ ;
 wire \u_neuron.u_syn/_071_ ;
 wire \u_neuron.u_syn/_072_ ;
 wire \u_neuron.u_syn/_073_ ;
 wire \u_neuron.u_syn/_074_ ;
 wire \u_neuron.u_syn/_075_ ;
 wire \u_neuron.u_syn/_076_ ;
 wire \u_neuron.u_syn/_077_ ;
 wire \u_neuron.u_syn/_078_ ;
 wire \u_neuron.u_syn/_079_ ;
 wire \u_neuron.u_syn/_080_ ;
 wire \u_neuron.u_syn/_081_ ;
 wire \u_neuron.u_syn/_082_ ;
 wire \u_neuron.u_syn/_083_ ;
 wire \u_neuron.u_syn/_084_ ;
 wire \u_neuron.u_syn/_085_ ;
 wire \u_neuron.u_syn/_086_ ;
 wire \u_neuron.u_syn/_087_ ;
 wire \u_neuron.u_syn/_088_ ;
 wire \u_neuron.u_syn/_089_ ;
 wire \u_neuron.u_syn/_090_ ;
 wire \u_neuron.u_syn/_091_ ;
 wire \u_neuron.u_syn/_092_ ;
 wire \u_neuron.u_syn/_093_ ;
 wire \u_neuron.u_syn/_094_ ;
 wire \u_neuron.u_syn/_095_ ;
 wire \u_neuron.u_syn/_096_ ;
 wire \u_neuron.u_syn/_097_ ;
 wire \u_neuron.u_syn/_098_ ;
 wire \u_neuron.u_syn/_099_ ;
 wire \u_neuron.u_syn/_100_ ;
 wire \u_neuron.u_syn/_101_ ;
 wire \u_neuron.u_syn/_102_ ;
 wire \u_neuron.u_syn/_103_ ;
 wire \u_neuron.u_syn/_104_ ;
 wire \u_neuron.u_syn/_105_ ;
 wire \u_neuron.u_syn/_106_ ;
 wire \u_neuron.u_syn/_107_ ;
 wire \u_neuron.u_syn/_108_ ;
 wire \u_neuron.u_syn/_109_ ;
 wire \u_neuron.u_syn/_110_ ;
 wire \u_neuron.u_syn/_111_ ;
 wire \u_neuron.u_syn/_112_ ;
 wire \u_neuron.u_syn/_113_ ;
 wire \u_neuron.u_syn/_114_ ;
 wire \u_neuron.u_syn/_115_ ;
 wire \u_neuron.u_syn/_116_ ;
 wire \u_neuron.u_syn/_117_ ;
 wire \u_neuron.u_syn/_118_ ;
 wire \u_neuron.u_syn/_119_ ;
 wire \u_neuron.u_syn/_120_ ;
 wire \u_neuron.u_syn/_121_ ;
 wire \u_neuron.u_syn/_122_ ;
 wire \u_neuron.u_syn/_123_ ;
 wire \u_neuron.u_syn/_124_ ;
 wire \u_neuron.u_syn/_125_ ;
 wire \u_neuron.u_syn/_126_ ;
 wire \u_neuron.u_syn/_127_ ;
 wire \u_neuron.u_syn/_128_ ;
 wire \u_neuron.u_syn/_129_ ;
 wire \u_neuron.u_syn/_130_ ;
 wire \u_neuron.u_syn/_131_ ;
 wire \u_neuron.u_syn/_132_ ;
 wire \u_neuron.u_syn/_133_ ;
 wire \u_neuron.u_syn/_134_ ;
 wire \u_neuron.u_syn/_135_ ;
 wire \u_neuron.u_syn/_136_ ;
 wire \u_neuron.u_syn/_137_ ;
 wire \u_neuron.u_syn/_138_ ;
 wire \u_neuron.u_syn/_139_ ;
 wire \u_neuron.u_syn/_140_ ;
 wire \u_neuron.u_syn/_141_ ;
 wire \u_neuron.u_syn/_142_ ;
 wire \u_neuron.u_syn/_143_ ;
 wire \u_neuron.u_syn/_144_ ;
 wire \u_neuron.u_syn/_145_ ;
 wire \u_neuron.u_syn/_146_ ;
 wire \u_neuron.u_syn/_147_ ;
 wire \u_neuron.u_syn/_148_ ;
 wire \u_neuron.u_syn/_149_ ;
 wire \u_neuron.u_syn/_150_ ;
 wire \u_neuron.u_syn/_151_ ;
 wire \u_neuron.u_syn/_152_ ;
 wire \u_neuron.u_syn/_153_ ;
 wire \u_neuron.u_syn/_154_ ;
 wire \u_neuron.u_syn/_155_ ;
 wire \u_neuron.u_syn/_156_ ;
 wire \u_neuron.u_syn/_157_ ;
 wire \u_neuron.u_syn/_158_ ;
 wire \u_neuron.u_syn/_159_ ;
 wire \u_neuron.u_syn/_160_ ;
 wire \u_neuron.u_syn/_161_ ;
 wire \u_neuron.u_syn/_162_ ;
 wire \u_neuron.u_syn/_163_ ;
 wire \u_neuron.u_syn/_164_ ;
 wire \u_neuron.u_syn/_165_ ;
 wire \u_neuron.u_syn/_166_ ;
 wire \u_neuron.u_syn/_167_ ;
 wire \u_neuron.u_syn/_168_ ;
 wire \u_neuron.u_syn/_169_ ;
 wire \u_neuron.u_syn/_170_ ;
 wire \u_neuron.u_syn/_171_ ;
 wire \u_neuron.u_syn/_172_ ;
 wire \u_neuron.u_syn/_173_ ;
 wire \u_neuron.u_syn/_174_ ;
 wire \u_neuron.u_syn/_175_ ;
 wire \u_neuron.u_syn/_176_ ;
 wire \u_neuron.u_syn/_177_ ;
 wire \u_neuron.u_syn/_178_ ;
 wire \u_neuron.u_syn/_179_ ;
 wire \u_neuron.u_syn/_180_ ;
 wire \u_neuron.u_syn/_181_ ;
 wire \u_neuron.u_syn/_182_ ;
 wire \u_neuron.u_syn/_183_ ;
 wire \u_neuron.u_syn/_184_ ;
 wire \u_neuron.u_syn/_185_ ;
 wire \u_neuron.u_syn/_186_ ;
 wire \u_neuron.u_syn/_187_ ;
 wire \u_neuron.u_syn/_188_ ;
 wire \u_neuron.u_syn/_189_ ;
 wire \u_neuron.u_syn/_190_ ;
 wire \u_neuron.u_syn/_191_ ;
 wire \u_neuron.u_syn/_192_ ;
 wire \u_neuron.u_syn/_193_ ;
 wire \u_neuron.u_syn/_194_ ;
 wire \u_neuron.u_syn/_195_ ;
 wire \u_neuron.u_syn/_196_ ;
 wire \u_neuron.u_syn/_197_ ;
 wire \u_neuron.u_syn/_198_ ;
 wire \u_neuron.u_syn/_199_ ;
 wire \u_neuron.u_syn/_200_ ;
 wire \u_neuron.u_syn/_201_ ;
 wire \u_neuron.u_syn/_202_ ;
 wire \u_neuron.u_syn/_203_ ;
 wire \u_neuron.u_syn/_204_ ;
 wire \u_neuron.u_syn/_205_ ;
 wire \u_neuron.u_syn/_206_ ;
 wire \u_neuron.u_syn/_207_ ;
 wire \u_neuron.u_syn/_208_ ;
 wire \u_neuron.u_syn/_209_ ;
 wire \u_neuron.u_syn/_210_ ;
 wire \u_neuron.u_syn/_211_ ;
 wire \u_neuron.u_syn/_212_ ;
 wire \u_neuron.u_syn/_213_ ;
 wire \u_neuron.u_syn/_214_ ;
 wire \u_neuron.u_syn/_215_ ;
 wire \u_neuron.u_syn/_216_ ;
 wire \u_neuron.u_syn/_217_ ;
 wire \u_neuron.u_syn/_218_ ;
 wire \u_neuron.u_syn/_219_ ;
 wire \u_neuron.u_syn/_220_ ;
 wire \u_neuron.u_syn/_221_ ;
 wire \u_neuron.u_syn/_222_ ;
 wire \u_neuron.u_syn/_223_ ;
 wire \u_neuron.u_syn/_224_ ;
 wire \u_neuron.u_syn/_225_ ;
 wire \u_neuron.u_syn/_226_ ;
 wire \u_neuron.u_syn/_227_ ;
 wire \u_neuron.u_syn/_228_ ;
 wire \u_neuron.u_syn/_229_ ;
 wire \u_neuron.u_syn/_230_ ;
 wire \u_neuron.u_syn/_231_ ;
 wire \u_neuron.u_syn/_232_ ;
 wire \u_neuron.u_syn/_233_ ;
 wire \u_neuron.u_syn/_234_ ;
 wire \u_neuron.u_syn/_235_ ;
 wire \u_neuron.u_syn/_236_ ;
 wire \u_neuron.u_syn/_237_ ;
 wire \u_neuron.u_syn/_238_ ;
 wire \u_neuron.u_syn/_239_ ;
 wire \u_neuron.u_syn/_240_ ;
 wire \u_neuron.u_syn/_241_ ;
 wire \u_neuron.u_syn/_242_ ;
 wire \u_neuron.u_syn/_243_ ;
 wire \u_neuron.u_syn/_244_ ;
 wire \u_neuron.u_syn/_245_ ;
 wire \u_neuron.u_syn/_246_ ;
 wire \u_neuron.u_syn/_247_ ;
 wire \u_neuron.u_syn/_248_ ;
 wire \u_neuron.u_syn/_249_ ;
 wire \u_neuron.u_syn/_250_ ;
 wire \u_neuron.u_syn/_251_ ;
 wire \u_neuron.u_syn/_252_ ;
 wire \u_neuron.u_syn/_253_ ;
 wire \u_neuron.u_syn/_254_ ;
 wire \u_neuron.u_syn/_255_ ;
 wire \u_neuron.u_syn/_256_ ;
 wire \u_neuron.u_syn/_257_ ;
 wire \u_neuron.u_syn/_258_ ;
 wire \u_neuron.u_syn/_259_ ;
 wire \u_neuron.u_syn/_260_ ;
 wire \u_neuron.u_syn/_261_ ;
 wire \u_neuron.u_syn/_262_ ;
 wire \u_neuron.u_syn/_263_ ;
 wire \u_neuron.u_syn/_264_ ;
 wire \u_neuron.u_syn/_265_ ;
 wire \u_neuron.u_syn/_266_ ;
 wire \u_neuron.u_syn/_267_ ;
 wire \u_neuron.u_syn/_268_ ;
 wire \u_neuron.u_syn/_269_ ;
 wire \u_neuron.u_syn/_270_ ;
 wire \u_neuron.u_syn/_271_ ;
 wire \u_neuron.u_syn/_272_ ;
 wire \u_neuron.u_syn/_273_ ;
 wire \u_neuron.u_syn/_274_ ;
 wire \u_neuron.u_syn/_275_ ;
 wire \u_neuron.u_syn/_276_ ;
 wire \u_neuron.u_syn/_277_ ;
 wire \u_neuron.u_syn/_278_ ;
 wire \u_neuron.u_syn/_279_ ;
 wire \u_neuron.u_syn/_280_ ;
 wire \u_neuron.u_syn/_281_ ;
 wire \u_neuron.u_syn/_282_ ;
 wire \u_neuron.u_syn/_283_ ;
 wire \u_neuron.u_syn/_284_ ;
 wire \u_neuron.u_syn/_285_ ;
 wire \u_neuron.u_syn/_286_ ;
 wire \u_neuron.u_syn/_287_ ;
 wire \u_neuron.u_syn/_288_ ;
 wire \u_neuron.u_syn/_289_ ;
 wire \u_neuron.u_syn/_290_ ;
 wire \u_neuron.u_syn/_291_ ;
 wire \u_neuron.u_syn/_292_ ;
 wire \u_neuron.u_syn/_293_ ;
 wire \u_neuron.u_syn/_294_ ;
 wire \u_neuron.u_syn/_295_ ;
 wire \u_neuron.u_syn/_296_ ;
 wire \u_neuron.u_syn/_297_ ;
 wire \u_neuron.u_syn/_298_ ;
 wire \u_neuron.u_syn/_299_ ;
 wire \u_neuron.u_syn/_300_ ;
 wire \u_neuron.u_syn/_301_ ;
 wire \u_neuron.u_syn/_302_ ;
 wire \u_neuron.u_syn/_303_ ;
 wire \u_neuron.u_syn/_304_ ;
 wire \u_neuron.u_syn/_305_ ;
 wire \u_neuron.u_syn/_306_ ;
 wire \u_neuron.u_syn/_307_ ;
 wire \u_neuron.u_syn/_308_ ;
 wire \u_neuron.u_syn/_309_ ;
 wire \u_neuron.u_syn/_310_ ;
 wire \u_neuron.u_syn/_311_ ;
 wire \u_neuron.u_syn/_312_ ;
 wire \u_neuron.u_syn/_313_ ;
 wire \u_neuron.u_syn/_314_ ;
 wire \u_neuron.u_syn/_315_ ;
 wire \u_neuron.u_syn/_316_ ;
 wire \u_neuron.u_syn/_317_ ;
 wire \u_neuron.u_syn/_318_ ;
 wire \u_neuron.u_syn/_319_ ;
 wire \u_neuron.u_syn/_320_ ;
 wire \u_neuron.u_syn/_321_ ;
 wire \u_neuron.u_syn/_322_ ;
 wire \u_neuron.u_syn/_323_ ;
 wire \u_neuron.u_syn/_324_ ;
 wire \u_neuron.u_syn/_325_ ;
 wire \u_neuron.u_syn/_326_ ;
 wire \u_neuron.u_syn/_327_ ;
 wire \u_neuron.u_syn/_328_ ;
 wire \u_neuron.u_syn/_329_ ;
 wire \u_neuron.u_syn/_330_ ;
 wire \u_neuron.u_syn/_331_ ;
 wire \u_neuron.u_syn/_332_ ;
 wire \u_neuron.u_syn/_333_ ;
 wire \u_neuron.u_syn/_334_ ;
 wire \u_neuron.u_syn/_335_ ;
 wire \u_neuron.u_syn/_336_ ;
 wire \u_neuron.u_syn/_337_ ;
 wire \u_neuron.u_syn/_338_ ;
 wire \u_neuron.u_syn/_339_ ;
 wire \u_neuron.u_syn/_340_ ;
 wire \u_neuron.u_syn/_341_ ;
 wire \u_neuron.u_syn/_342_ ;
 wire \u_neuron.u_syn/_343_ ;
 wire \u_neuron.u_syn/_344_ ;
 wire \u_neuron.u_syn/_345_ ;
 wire \u_neuron.u_syn/_346_ ;
 wire \u_neuron.u_syn/_347_ ;
 wire \u_neuron.u_syn/_348_ ;
 wire \u_neuron.u_syn/_349_ ;
 wire \u_neuron.u_syn/_350_ ;
 wire \u_neuron.u_syn/_351_ ;
 wire \u_neuron.u_syn/_352_ ;
 wire \u_neuron.u_syn/_353_ ;
 wire \u_neuron.u_syn/_354_ ;
 wire \u_neuron.u_syn/_355_ ;
 wire \u_neuron.u_syn/_356_ ;
 wire \u_neuron.u_syn/_357_ ;
 wire \u_neuron.u_syn/_358_ ;
 wire \u_neuron.u_syn/_359_ ;
 wire \u_neuron.u_syn/_360_ ;
 wire \u_neuron.u_syn/_361_ ;
 wire \u_neuron.u_syn/_362_ ;
 wire \u_neuron.u_syn/_363_ ;
 wire \u_neuron.u_syn/_364_ ;
 wire \u_neuron.u_syn/_365_ ;
 wire \u_neuron.u_syn/_366_ ;
 wire \u_neuron.u_syn/_367_ ;
 wire \u_neuron.u_syn/_368_ ;
 wire \u_neuron.u_syn/_369_ ;
 wire \u_neuron.u_syn/_370_ ;
 wire \u_neuron.u_syn/_371_ ;
 wire \u_neuron.u_syn/_372_ ;
 wire \u_neuron.u_syn/_373_ ;
 wire \u_neuron.u_syn/_374_ ;
 wire \u_neuron.u_syn/_375_ ;
 wire \u_neuron.u_syn/_376_ ;
 wire \u_neuron.u_syn/_377_ ;
 wire \u_neuron.u_syn/_378_ ;
 wire \u_neuron.u_syn/_379_ ;
 wire \u_neuron.u_syn/_380_ ;
 wire \u_neuron.u_syn/_381_ ;
 wire \u_neuron.u_syn/_382_ ;
 wire \u_neuron.u_syn/_383_ ;
 wire \u_neuron.u_syn/_384_ ;
 wire \u_neuron.u_syn/_385_ ;
 wire \u_neuron.u_syn/_386_ ;
 wire \u_neuron.u_syn/_387_ ;
 wire \u_neuron.u_syn/_388_ ;
 wire \u_neuron.u_syn/_389_ ;
 wire \u_neuron.u_syn/_390_ ;
 wire \u_neuron.u_syn/_391_ ;
 wire \u_neuron.u_syn/_392_ ;
 wire \u_neuron.u_syn/_393_ ;
 wire \u_neuron.u_syn/_394_ ;
 wire \u_neuron.u_syn/_395_ ;
 wire \u_neuron.u_syn/_396_ ;
 wire \u_neuron.u_syn/_397_ ;
 wire \u_neuron.u_syn/_398_ ;
 wire \u_neuron.u_syn/_399_ ;
 wire \u_neuron.u_syn/_400_ ;
 wire \u_neuron.u_syn/_401_ ;
 wire \u_neuron.u_syn/_402_ ;
 wire \u_neuron.u_syn/_403_ ;
 wire \u_neuron.u_syn/_404_ ;
 wire \u_neuron.u_td/_000_ ;
 wire \u_neuron.u_td/_001_ ;
 wire \u_neuron.u_td/_002_ ;
 wire \u_neuron.u_td/_003_ ;
 wire \u_neuron.u_td/_004_ ;
 wire \u_neuron.u_td/_005_ ;
 wire \u_neuron.u_td/_006_ ;
 wire \u_neuron.u_td/_007_ ;
 wire \u_neuron.u_td/_008_ ;
 wire \u_neuron.u_td/_009_ ;
 wire \u_neuron.u_td/_010_ ;
 wire \u_neuron.u_td/_011_ ;
 wire \u_neuron.u_td/_012_ ;
 wire \u_neuron.u_td/_013_ ;
 wire \u_neuron.u_td/_014_ ;
 wire \u_neuron.u_td/_015_ ;
 wire \u_neuron.u_td/_016_ ;
 wire \u_neuron.u_td/_017_ ;
 wire \u_neuron.u_td/_018_ ;
 wire \u_neuron.u_td/_019_ ;
 wire \u_neuron.u_td/_020_ ;
 wire \u_neuron.u_td/_021_ ;
 wire \u_neuron.u_td/_022_ ;
 wire \u_neuron.u_td/_023_ ;
 wire \u_neuron.u_td/_024_ ;
 wire \u_neuron.u_td/_025_ ;
 wire \u_neuron.u_td/_026_ ;
 wire \u_neuron.u_td/_027_ ;
 wire \u_neuron.u_td/_028_ ;
 wire \u_neuron.u_td/_029_ ;
 wire \u_neuron.u_td/_030_ ;
 wire \u_neuron.u_td/_031_ ;
 wire \u_neuron.u_td/_032_ ;
 wire \u_neuron.u_td/_033_ ;
 wire \u_neuron.u_td/_034_ ;
 wire \u_neuron.u_td/_035_ ;
 wire \u_neuron.u_td/_036_ ;
 wire \u_neuron.u_td/_037_ ;
 wire \u_neuron.u_td/_038_ ;
 wire \u_neuron.u_td/_039_ ;
 wire \u_neuron.u_td/_040_ ;
 wire \u_neuron.u_td/_041_ ;
 wire \u_neuron.u_td/_042_ ;
 wire \u_neuron.u_td/_043_ ;
 wire \u_neuron.u_td/_044_ ;
 wire \u_neuron.u_td/_045_ ;
 wire \u_neuron.u_td/_046_ ;
 wire \u_neuron.u_td/_047_ ;
 wire \u_neuron.u_td/_048_ ;
 wire \u_neuron.u_td/_049_ ;
 wire \u_neuron.u_td/_050_ ;
 wire \u_neuron.u_td/_051_ ;
 wire \u_neuron.u_td/_052_ ;
 wire \u_neuron.u_td/_053_ ;
 wire \u_neuron.u_td/_054_ ;
 wire \u_neuron.u_td/_055_ ;
 wire \u_neuron.u_td/_056_ ;
 wire \u_neuron.u_td/_057_ ;
 wire \u_neuron.u_td/_058_ ;
 wire \u_neuron.u_td/_059_ ;
 wire \u_neuron.u_td/_060_ ;
 wire \u_neuron.u_td/_061_ ;
 wire \u_neuron.u_td/_062_ ;
 wire \u_neuron.u_td/_063_ ;
 wire \u_neuron.u_td/_064_ ;
 wire \u_neuron.u_td/_065_ ;
 wire \u_neuron.u_td/_066_ ;
 wire \u_neuron.u_td/_067_ ;
 wire \u_neuron.u_td/_068_ ;
 wire \u_neuron.u_td/_069_ ;
 wire \u_neuron.u_td/_070_ ;
 wire \u_neuron.u_td/_071_ ;
 wire \u_neuron.u_td/_072_ ;
 wire \u_neuron.u_td/_073_ ;
 wire \u_neuron.u_td/_074_ ;
 wire \u_neuron.u_td/_075_ ;
 wire \u_neuron.u_td/_076_ ;
 wire \u_neuron.u_td/_077_ ;
 wire \u_neuron.u_td/_078_ ;
 wire \u_neuron.u_td/_079_ ;
 wire \u_neuron.u_td/_080_ ;
 wire \u_neuron.u_td/_081_ ;
 wire \u_neuron.u_td/_082_ ;
 wire \u_neuron.u_td/_083_ ;
 wire \u_neuron.u_td/_084_ ;
 wire \u_neuron.u_td/_085_ ;
 wire \u_neuron.u_td/_086_ ;
 wire \u_neuron.u_td/_087_ ;
 wire \u_neuron.u_td/_088_ ;
 wire \u_neuron.u_td/_089_ ;
 wire \u_neuron.u_td/_090_ ;
 wire \u_neuron.u_td/_091_ ;
 wire \u_neuron.u_td/_092_ ;
 wire \u_neuron.u_td/_093_ ;
 wire \u_neuron.u_td/_094_ ;
 wire \u_neuron.u_td/_095_ ;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire clknet_5_0__leaf_clk;
 wire clknet_5_1__leaf_clk;
 wire clknet_5_2__leaf_clk;
 wire clknet_5_3__leaf_clk;
 wire clknet_5_4__leaf_clk;
 wire clknet_5_5__leaf_clk;
 wire clknet_5_6__leaf_clk;
 wire clknet_5_7__leaf_clk;
 wire clknet_5_8__leaf_clk;
 wire clknet_5_9__leaf_clk;
 wire clknet_5_10__leaf_clk;
 wire clknet_5_11__leaf_clk;
 wire clknet_5_12__leaf_clk;
 wire clknet_5_13__leaf_clk;
 wire clknet_5_14__leaf_clk;
 wire clknet_5_15__leaf_clk;
 wire clknet_5_16__leaf_clk;
 wire clknet_5_17__leaf_clk;
 wire clknet_5_18__leaf_clk;
 wire clknet_5_19__leaf_clk;
 wire clknet_5_20__leaf_clk;
 wire clknet_5_21__leaf_clk;
 wire clknet_5_22__leaf_clk;
 wire clknet_5_23__leaf_clk;
 wire clknet_5_24__leaf_clk;
 wire clknet_5_25__leaf_clk;
 wire clknet_5_26__leaf_clk;
 wire clknet_5_27__leaf_clk;
 wire clknet_5_28__leaf_clk;
 wire clknet_5_29__leaf_clk;
 wire clknet_5_30__leaf_clk;
 wire clknet_5_31__leaf_clk;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;

 sg13g2_inv_2 _248_ (.Y(\u_neuron.stream_act ),
    .A(_002_));
 sg13g2_inv_1 _249_ (.Y(_064_),
    .A(\u_neuron.cfg_op[0] ));
 sg13g2_inv_1 _250_ (.Y(_065_),
    .A(net433));
 sg13g2_nand2_1 _251_ (.Y(_066_),
    .A(\u_neuron.is_cfg_cmd ),
    .B(\u_neuron.in_fire ));
 sg13g2_nor3_1 _252_ (.A(\u_neuron.cfg_op[1] ),
    .B(_064_),
    .C(_066_),
    .Y(_001_));
 sg13g2_nor3_1 _253_ (.A(\u_neuron.cfg_op[1] ),
    .B(\u_neuron.cfg_op[0] ),
    .C(_066_),
    .Y(_000_));
 sg13g2_nand2b_2 _254_ (.Y(_067_),
    .B(\u_neuron.in_fire ),
    .A_N(\u_neuron.is_special_cmd ));
 sg13g2_inv_1 _255_ (.Y(\u_neuron.normal_event ),
    .A(_067_));
 sg13g2_and3_1 _256_ (.X(\u_neuron.mode_conv_evt ),
    .A(net431),
    .B(net433),
    .C(net356));
 sg13g2_and3_2 _257_ (.X(\u_neuron.mode_fst_evt ),
    .A(net431),
    .B(_065_),
    .C(\u_neuron.normal_event ));
 sg13g2_nor3_1 _258_ (.A(net431),
    .B(_065_),
    .C(_067_),
    .Y(\u_neuron.mode_td_evt ));
 sg13g2_nor3_1 _259_ (.A(net431),
    .B(net433),
    .C(_067_),
    .Y(\u_neuron.mode_lif_evt ));
 sg13g2_and2_1 _260_ (.A(net378),
    .B(\u_neuron.in_fire ),
    .X(\u_neuron.soft_reset_fire ));
 sg13g2_and2_1 _261_ (.A(\u_neuron.in_fire ),
    .B(\u_neuron.is_arm_cmd ),
    .X(\u_neuron.arm_event ));
 sg13g2_mux4_1 _262_ (.S0(net428),
    .A0(\u_neuron.wtab[16] ),
    .A1(\u_neuron.wtab[18] ),
    .A2(\u_neuron.wtab[20] ),
    .A3(\u_neuron.wtab[22] ),
    .S1(net425),
    .X(_068_));
 sg13g2_nor2_1 _263_ (.A(net423),
    .B(_068_),
    .Y(_069_));
 sg13g2_nand2_1 _264_ (.Y(_070_),
    .A(net430),
    .B(\u_neuron.wtab[26] ));
 sg13g2_nand2b_1 _265_ (.Y(_071_),
    .B(\u_neuron.wtab[24] ),
    .A_N(net430));
 sg13g2_a21oi_1 _266_ (.A1(_070_),
    .A2(_071_),
    .Y(_072_),
    .B1(net426));
 sg13g2_nor2b_1 _267_ (.A(\u_neuron.wtab[30] ),
    .B_N(net428),
    .Y(_073_));
 sg13g2_o21ai_1 _268_ (.B1(net426),
    .Y(_074_),
    .A1(net428),
    .A2(\u_neuron.wtab[28] ));
 sg13g2_o21ai_1 _269_ (.B1(net423),
    .Y(_075_),
    .A1(_073_),
    .A2(_074_));
 sg13g2_o21ai_1 _270_ (.B1(net420),
    .Y(_076_),
    .A1(_072_),
    .A2(_075_));
 sg13g2_mux2_1 _271_ (.A0(\u_neuron.wtab[8] ),
    .A1(\u_neuron.wtab[10] ),
    .S(net429),
    .X(_077_));
 sg13g2_mux2_1 _272_ (.A0(\u_neuron.wtab[12] ),
    .A1(\u_neuron.wtab[14] ),
    .S(net429),
    .X(_078_));
 sg13g2_mux2_1 _273_ (.A0(\u_neuron.wtab[4] ),
    .A1(\u_neuron.wtab[6] ),
    .S(net429),
    .X(_079_));
 sg13g2_mux2_1 _274_ (.A0(\u_neuron.wtab[0] ),
    .A1(\u_neuron.wtab[2] ),
    .S(net429),
    .X(_080_));
 sg13g2_mux4_1 _275_ (.S0(net426),
    .A0(_080_),
    .A1(_079_),
    .A2(_077_),
    .A3(_078_),
    .S1(net423),
    .X(_081_));
 sg13g2_nand2b_1 _276_ (.Y(_082_),
    .B(_081_),
    .A_N(net420));
 sg13g2_o21ai_1 _277_ (.B1(_082_),
    .Y(\u_neuron.w_ptr_curr[0] ),
    .A1(_069_),
    .A2(_076_));
 sg13g2_mux4_1 _278_ (.S0(net430),
    .A0(\u_neuron.wtab[17] ),
    .A1(\u_neuron.wtab[19] ),
    .A2(\u_neuron.wtab[21] ),
    .A3(\u_neuron.wtab[23] ),
    .S1(net426),
    .X(_083_));
 sg13g2_nor2_1 _279_ (.A(net423),
    .B(_083_),
    .Y(_084_));
 sg13g2_nand2_1 _280_ (.Y(_085_),
    .A(net430),
    .B(\u_neuron.wtab[27] ));
 sg13g2_nand2b_1 _281_ (.Y(_086_),
    .B(\u_neuron.wtab[25] ),
    .A_N(net430));
 sg13g2_a21oi_1 _282_ (.A1(_085_),
    .A2(_086_),
    .Y(_087_),
    .B1(net426));
 sg13g2_nor2b_1 _283_ (.A(\u_neuron.wtab[31] ),
    .B_N(net428),
    .Y(_088_));
 sg13g2_o21ai_1 _284_ (.B1(net426),
    .Y(_089_),
    .A1(\u_neuron.learn_ptr[0] ),
    .A2(\u_neuron.wtab[29] ));
 sg13g2_o21ai_1 _285_ (.B1(net423),
    .Y(_090_),
    .A1(_088_),
    .A2(_089_));
 sg13g2_o21ai_1 _286_ (.B1(net420),
    .Y(_091_),
    .A1(_087_),
    .A2(_090_));
 sg13g2_mux2_1 _287_ (.A0(\u_neuron.wtab[5] ),
    .A1(\u_neuron.wtab[7] ),
    .S(net429),
    .X(_092_));
 sg13g2_mux2_1 _288_ (.A0(\u_neuron.wtab[1] ),
    .A1(\u_neuron.wtab[3] ),
    .S(net430),
    .X(_093_));
 sg13g2_mux2_1 _289_ (.A0(\u_neuron.wtab[13] ),
    .A1(\u_neuron.wtab[15] ),
    .S(net429),
    .X(_094_));
 sg13g2_mux2_1 _290_ (.A0(\u_neuron.wtab[9] ),
    .A1(\u_neuron.wtab[11] ),
    .S(net429),
    .X(_095_));
 sg13g2_mux4_1 _291_ (.S0(net423),
    .A0(_093_),
    .A1(_095_),
    .A2(_092_),
    .A3(_094_),
    .S1(net426),
    .X(_096_));
 sg13g2_nand2b_1 _292_ (.Y(_097_),
    .B(_096_),
    .A_N(net420));
 sg13g2_o21ai_1 _293_ (.B1(_097_),
    .Y(\u_neuron.w_ptr_curr[1] ),
    .A1(_084_),
    .A2(_091_));
 sg13g2_mux4_1 _294_ (.S0(net398),
    .A0(\u_neuron.wtab[16] ),
    .A1(\u_neuron.wtab[18] ),
    .A2(\u_neuron.wtab[20] ),
    .A3(\u_neuron.wtab[22] ),
    .S1(net391),
    .X(_098_));
 sg13g2_nor2_1 _295_ (.A(net389),
    .B(_098_),
    .Y(_099_));
 sg13g2_nand2_1 _296_ (.Y(_100_),
    .A(\u_neuron.wtab[26] ),
    .B(net397));
 sg13g2_nand2b_1 _297_ (.Y(_101_),
    .B(\u_neuron.wtab[24] ),
    .A_N(net397));
 sg13g2_a21oi_1 _298_ (.A1(_100_),
    .A2(_101_),
    .Y(_102_),
    .B1(net391));
 sg13g2_nor2b_1 _299_ (.A(\u_neuron.wtab[30] ),
    .B_N(net396),
    .Y(_103_));
 sg13g2_o21ai_1 _300_ (.B1(net392),
    .Y(_104_),
    .A1(\u_neuron.wtab[28] ),
    .A2(net396));
 sg13g2_o21ai_1 _301_ (.B1(net389),
    .Y(_105_),
    .A1(_103_),
    .A2(_104_));
 sg13g2_o21ai_1 _302_ (.B1(net386),
    .Y(_106_),
    .A1(_102_),
    .A2(_105_));
 sg13g2_mux2_1 _303_ (.A0(\u_neuron.wtab[4] ),
    .A1(\u_neuron.wtab[6] ),
    .S(net400),
    .X(_107_));
 sg13g2_mux2_1 _304_ (.A0(\u_neuron.wtab[0] ),
    .A1(\u_neuron.wtab[2] ),
    .S(net401),
    .X(_108_));
 sg13g2_mux2_1 _305_ (.A0(\u_neuron.wtab[12] ),
    .A1(\u_neuron.wtab[14] ),
    .S(net400),
    .X(_109_));
 sg13g2_mux2_1 _306_ (.A0(\u_neuron.wtab[8] ),
    .A1(\u_neuron.wtab[10] ),
    .S(net402),
    .X(_110_));
 sg13g2_mux4_1 _307_ (.S0(net390),
    .A0(_108_),
    .A1(_110_),
    .A2(_107_),
    .A3(_109_),
    .S1(net394),
    .X(_111_));
 sg13g2_nand2b_1 _308_ (.Y(_112_),
    .B(_111_),
    .A_N(net386));
 sg13g2_o21ai_1 _309_ (.B1(_112_),
    .Y(\u_neuron.w_addr_curr[0] ),
    .A1(_099_),
    .A2(_106_));
 sg13g2_mux4_1 _310_ (.S0(net398),
    .A0(\u_neuron.wtab[17] ),
    .A1(\u_neuron.wtab[19] ),
    .A2(\u_neuron.wtab[21] ),
    .A3(\u_neuron.wtab[23] ),
    .S1(net391),
    .X(_113_));
 sg13g2_nor2_1 _311_ (.A(net389),
    .B(_113_),
    .Y(_114_));
 sg13g2_nand2_1 _312_ (.Y(_115_),
    .A(\u_neuron.wtab[27] ),
    .B(net397));
 sg13g2_nand2b_1 _313_ (.Y(_116_),
    .B(\u_neuron.wtab[25] ),
    .A_N(net397));
 sg13g2_a21oi_1 _314_ (.A1(_115_),
    .A2(_116_),
    .Y(_117_),
    .B1(net391));
 sg13g2_nor2b_1 _315_ (.A(\u_neuron.wtab[31] ),
    .B_N(net396),
    .Y(_118_));
 sg13g2_o21ai_1 _316_ (.B1(net392),
    .Y(_119_),
    .A1(\u_neuron.wtab[29] ),
    .A2(net396));
 sg13g2_o21ai_1 _317_ (.B1(net389),
    .Y(_120_),
    .A1(_118_),
    .A2(_119_));
 sg13g2_o21ai_1 _318_ (.B1(net387),
    .Y(_121_),
    .A1(_117_),
    .A2(_120_));
 sg13g2_mux2_1 _319_ (.A0(\u_neuron.wtab[5] ),
    .A1(\u_neuron.wtab[7] ),
    .S(net402),
    .X(_122_));
 sg13g2_mux2_1 _320_ (.A0(\u_neuron.wtab[1] ),
    .A1(\u_neuron.wtab[3] ),
    .S(net402),
    .X(_123_));
 sg13g2_mux2_1 _321_ (.A0(\u_neuron.wtab[13] ),
    .A1(\u_neuron.wtab[15] ),
    .S(net400),
    .X(_124_));
 sg13g2_mux2_1 _322_ (.A0(\u_neuron.wtab[9] ),
    .A1(\u_neuron.wtab[11] ),
    .S(net402),
    .X(_125_));
 sg13g2_mux4_1 _323_ (.S0(net390),
    .A0(_123_),
    .A1(_125_),
    .A2(_122_),
    .A3(_124_),
    .S1(net395),
    .X(_126_));
 sg13g2_nand2b_1 _324_ (.Y(_127_),
    .B(_126_),
    .A_N(net387));
 sg13g2_o21ai_1 _325_ (.B1(_127_),
    .Y(\u_neuron.w_addr_curr[1] ),
    .A1(_114_),
    .A2(_121_));
 sg13g2_nand2b_1 _326_ (.Y(_128_),
    .B(\u_neuron.is_cfg_cmd ),
    .A_N(net378));
 sg13g2_nand3_1 _327_ (.B(net469),
    .C(_128_),
    .A(\u_neuron.in_fire ),
    .Y(_129_));
 sg13g2_nand2b_1 _328_ (.Y(_130_),
    .B(\u_neuron.conv_last_sum_next[0] ),
    .A_N(net374));
 sg13g2_nand2_1 _329_ (.Y(_131_),
    .A(net76),
    .B(net344));
 sg13g2_o21ai_1 _330_ (.B1(_131_),
    .Y(_003_),
    .A1(net344),
    .A2(_130_));
 sg13g2_nand2b_1 _331_ (.Y(_132_),
    .B(\u_neuron.conv_last_sum_next[1] ),
    .A_N(net374));
 sg13g2_nand2_1 _332_ (.Y(_133_),
    .A(net83),
    .B(net346));
 sg13g2_o21ai_1 _333_ (.B1(_133_),
    .Y(_004_),
    .A1(net344),
    .A2(_132_));
 sg13g2_nand2b_1 _334_ (.Y(_134_),
    .B(\u_neuron.conv_last_sum_next[2] ),
    .A_N(net374));
 sg13g2_nand2_1 _335_ (.Y(_135_),
    .A(net72),
    .B(net345));
 sg13g2_o21ai_1 _336_ (.B1(_135_),
    .Y(_005_),
    .A1(net345),
    .A2(_134_));
 sg13g2_nand2b_1 _337_ (.Y(_136_),
    .B(\u_neuron.td_last_diff_next[0] ),
    .A_N(net373));
 sg13g2_nand2_1 _338_ (.Y(_137_),
    .A(net68),
    .B(net340));
 sg13g2_o21ai_1 _339_ (.B1(_137_),
    .Y(_006_),
    .A1(net340),
    .A2(_136_));
 sg13g2_nand2b_1 _340_ (.Y(_138_),
    .B(\u_neuron.td_last_diff_next[1] ),
    .A_N(net374));
 sg13g2_nand2_1 _341_ (.Y(_139_),
    .A(net75),
    .B(net344));
 sg13g2_o21ai_1 _342_ (.B1(_139_),
    .Y(_007_),
    .A1(net345),
    .A2(_138_));
 sg13g2_nand2b_1 _343_ (.Y(_140_),
    .B(\u_neuron.td_last_diff_next[2] ),
    .A_N(net374));
 sg13g2_nand2_1 _344_ (.Y(_141_),
    .A(net84),
    .B(net344));
 sg13g2_o21ai_1 _345_ (.B1(_141_),
    .Y(_008_),
    .A1(net344),
    .A2(_140_));
 sg13g2_nand2b_1 _346_ (.Y(_142_),
    .B(\u_neuron.td_last_diff_next[3] ),
    .A_N(net374));
 sg13g2_nand2_1 _347_ (.Y(_143_),
    .A(net79),
    .B(net344));
 sg13g2_o21ai_1 _348_ (.B1(_143_),
    .Y(_009_),
    .A1(net344),
    .A2(_142_));
 sg13g2_nand2b_1 _349_ (.Y(_144_),
    .B(\u_neuron.td_last_diff_next[4] ),
    .A_N(net372));
 sg13g2_nand2_1 _350_ (.Y(_145_),
    .A(net61),
    .B(net341));
 sg13g2_o21ai_1 _351_ (.B1(_145_),
    .Y(_010_),
    .A1(net341),
    .A2(_144_));
 sg13g2_nand2b_1 _352_ (.Y(_146_),
    .B(\u_neuron.td_last_diff_next[5] ),
    .A_N(net372));
 sg13g2_nand2_1 _353_ (.Y(_147_),
    .A(net80),
    .B(net340));
 sg13g2_o21ai_1 _354_ (.B1(_147_),
    .Y(_011_),
    .A1(net340),
    .A2(_146_));
 sg13g2_nand2b_1 _355_ (.Y(_148_),
    .B(\u_neuron.td_last_diff_next[6] ),
    .A_N(net372));
 sg13g2_nand2_1 _356_ (.Y(_149_),
    .A(net87),
    .B(net341));
 sg13g2_o21ai_1 _357_ (.B1(_149_),
    .Y(_012_),
    .A1(net341),
    .A2(_148_));
 sg13g2_nand2b_1 _358_ (.Y(_150_),
    .B(\u_neuron.td_last_diff_next[7] ),
    .A_N(net372));
 sg13g2_nand2_1 _359_ (.Y(_151_),
    .A(net64),
    .B(net341));
 sg13g2_o21ai_1 _360_ (.B1(_151_),
    .Y(_013_),
    .A1(net341),
    .A2(_150_));
 sg13g2_nand2b_1 _361_ (.Y(_152_),
    .B(\u_neuron.fst_t_next[0] ),
    .A_N(net376));
 sg13g2_nand2_1 _362_ (.Y(_153_),
    .A(net130),
    .B(net349));
 sg13g2_o21ai_1 _363_ (.B1(_153_),
    .Y(_014_),
    .A1(net349),
    .A2(_152_));
 sg13g2_nand2b_1 _364_ (.Y(_154_),
    .B(\u_neuron.fst_t_next[1] ),
    .A_N(net376));
 sg13g2_nand2_1 _365_ (.Y(_155_),
    .A(net192),
    .B(net349));
 sg13g2_o21ai_1 _366_ (.B1(_155_),
    .Y(_015_),
    .A1(net349),
    .A2(_154_));
 sg13g2_nand2b_1 _367_ (.Y(_156_),
    .B(\u_neuron.fst_t_next[2] ),
    .A_N(net377));
 sg13g2_nand2_1 _368_ (.Y(_157_),
    .A(net135),
    .B(net347));
 sg13g2_o21ai_1 _369_ (.B1(_157_),
    .Y(_016_),
    .A1(net349),
    .A2(_156_));
 sg13g2_nand2b_1 _370_ (.Y(_158_),
    .B(\u_neuron.fst_t_next[3] ),
    .A_N(net377));
 sg13g2_nand2_1 _371_ (.Y(_159_),
    .A(net123),
    .B(net350));
 sg13g2_o21ai_1 _372_ (.B1(_159_),
    .Y(_017_),
    .A1(net347),
    .A2(_158_));
 sg13g2_nand2b_1 _373_ (.Y(_160_),
    .B(\u_neuron.fst_t_next[4] ),
    .A_N(net377));
 sg13g2_nand2_1 _374_ (.Y(_161_),
    .A(net159),
    .B(net347));
 sg13g2_o21ai_1 _375_ (.B1(_161_),
    .Y(_018_),
    .A1(net347),
    .A2(_160_));
 sg13g2_nand2b_1 _376_ (.Y(_162_),
    .B(\u_neuron.fst_t_next[5] ),
    .A_N(net377));
 sg13g2_nand2_1 _377_ (.Y(_163_),
    .A(net116),
    .B(net347));
 sg13g2_o21ai_1 _378_ (.B1(_163_),
    .Y(_019_),
    .A1(net347),
    .A2(_162_));
 sg13g2_nand2b_1 _379_ (.Y(_164_),
    .B(\u_neuron.fst_t_next[6] ),
    .A_N(net376));
 sg13g2_nand2_1 _380_ (.Y(_165_),
    .A(net136),
    .B(net348));
 sg13g2_o21ai_1 _381_ (.B1(_165_),
    .Y(_020_),
    .A1(net348),
    .A2(_164_));
 sg13g2_nand2b_1 _382_ (.Y(_166_),
    .B(\u_neuron.fst_t_next[7] ),
    .A_N(net376));
 sg13g2_nand2_1 _383_ (.Y(_167_),
    .A(net133),
    .B(net348));
 sg13g2_o21ai_1 _384_ (.B1(_167_),
    .Y(_021_),
    .A1(net348),
    .A2(_166_));
 sg13g2_nand2b_1 _385_ (.Y(_168_),
    .B(\u_neuron.td_prev_next[0] ),
    .A_N(net372));
 sg13g2_nand2_1 _386_ (.Y(_169_),
    .A(net126),
    .B(net340));
 sg13g2_o21ai_1 _387_ (.B1(_169_),
    .Y(_022_),
    .A1(net340),
    .A2(_168_));
 sg13g2_nand2b_1 _388_ (.Y(_170_),
    .B(\u_neuron.td_prev_next[1] ),
    .A_N(net370));
 sg13g2_nand2_1 _389_ (.Y(_171_),
    .A(net114),
    .B(net337));
 sg13g2_o21ai_1 _390_ (.B1(_171_),
    .Y(_023_),
    .A1(net337),
    .A2(_170_));
 sg13g2_nand2b_1 _391_ (.Y(_172_),
    .B(\u_neuron.td_prev_next[2] ),
    .A_N(net369));
 sg13g2_nand2_1 _392_ (.Y(_173_),
    .A(net118),
    .B(net337));
 sg13g2_o21ai_1 _393_ (.B1(_173_),
    .Y(_024_),
    .A1(net337),
    .A2(_172_));
 sg13g2_nand2b_1 _394_ (.Y(_174_),
    .B(\u_neuron.td_prev_next[3] ),
    .A_N(net369));
 sg13g2_nand2_1 _395_ (.Y(_175_),
    .A(net140),
    .B(net335));
 sg13g2_o21ai_1 _396_ (.B1(_175_),
    .Y(_025_),
    .A1(net335),
    .A2(_174_));
 sg13g2_nand2b_1 _397_ (.Y(_176_),
    .B(\u_neuron.td_prev_next[4] ),
    .A_N(net369));
 sg13g2_nand2_1 _398_ (.Y(_177_),
    .A(net151),
    .B(net334));
 sg13g2_o21ai_1 _399_ (.B1(_177_),
    .Y(_026_),
    .A1(net334),
    .A2(_176_));
 sg13g2_nand2b_1 _400_ (.Y(_178_),
    .B(\u_neuron.td_prev_next[5] ),
    .A_N(net369));
 sg13g2_nand2_1 _401_ (.Y(_179_),
    .A(net144),
    .B(net334));
 sg13g2_o21ai_1 _402_ (.B1(_179_),
    .Y(_027_),
    .A1(net334),
    .A2(_178_));
 sg13g2_nand2b_1 _403_ (.Y(_180_),
    .B(\u_neuron.td_prev_next[6] ),
    .A_N(net370));
 sg13g2_nand2_1 _404_ (.Y(_181_),
    .A(net112),
    .B(net336));
 sg13g2_o21ai_1 _405_ (.B1(_181_),
    .Y(_028_),
    .A1(net336),
    .A2(_180_));
 sg13g2_nand2b_1 _406_ (.Y(_182_),
    .B(\u_neuron.td_prev_next[7] ),
    .A_N(net372));
 sg13g2_nand2_1 _407_ (.Y(_183_),
    .A(net131),
    .B(net340));
 sg13g2_o21ai_1 _408_ (.B1(_183_),
    .Y(_029_),
    .A1(net340),
    .A2(_182_));
 sg13g2_nand2b_1 _409_ (.Y(_184_),
    .B(\u_neuron.fst_last_t_next[0] ),
    .A_N(net376));
 sg13g2_nand2_1 _410_ (.Y(_185_),
    .A(net59),
    .B(net349));
 sg13g2_o21ai_1 _411_ (.B1(_185_),
    .Y(_030_),
    .A1(net349),
    .A2(_184_));
 sg13g2_nand2b_1 _412_ (.Y(_186_),
    .B(\u_neuron.fst_last_t_next[1] ),
    .A_N(net377));
 sg13g2_nand2_1 _413_ (.Y(_187_),
    .A(net109),
    .B(net351));
 sg13g2_o21ai_1 _414_ (.B1(_187_),
    .Y(_031_),
    .A1(net351),
    .A2(_186_));
 sg13g2_nand2b_1 _415_ (.Y(_188_),
    .B(\u_neuron.fst_last_t_next[2] ),
    .A_N(net377));
 sg13g2_nand2_1 _416_ (.Y(_189_),
    .A(net104),
    .B(net351));
 sg13g2_o21ai_1 _417_ (.B1(_189_),
    .Y(_032_),
    .A1(net351),
    .A2(_188_));
 sg13g2_nand2b_1 _418_ (.Y(_190_),
    .B(\u_neuron.fst_last_t_next[3] ),
    .A_N(net375));
 sg13g2_nand2_1 _419_ (.Y(_191_),
    .A(net88),
    .B(net345));
 sg13g2_o21ai_1 _420_ (.B1(_191_),
    .Y(_033_),
    .A1(net345),
    .A2(_190_));
 sg13g2_nand2b_1 _421_ (.Y(_192_),
    .B(\u_neuron.fst_last_t_next[4] ),
    .A_N(net375));
 sg13g2_nand2_1 _422_ (.Y(_193_),
    .A(net62),
    .B(net345));
 sg13g2_o21ai_1 _423_ (.B1(_193_),
    .Y(_034_),
    .A1(net345),
    .A2(_192_));
 sg13g2_nand2b_1 _424_ (.Y(_194_),
    .B(\u_neuron.fst_last_t_next[5] ),
    .A_N(net376));
 sg13g2_nand2_1 _425_ (.Y(_195_),
    .A(net66),
    .B(net347));
 sg13g2_o21ai_1 _426_ (.B1(_195_),
    .Y(_035_),
    .A1(net347),
    .A2(_194_));
 sg13g2_nand2b_1 _427_ (.Y(_196_),
    .B(\u_neuron.fst_last_t_next[6] ),
    .A_N(net376));
 sg13g2_nand2_1 _428_ (.Y(_197_),
    .A(net73),
    .B(net348));
 sg13g2_o21ai_1 _429_ (.B1(_197_),
    .Y(_036_),
    .A1(net348),
    .A2(_196_));
 sg13g2_nand2b_1 _430_ (.Y(_198_),
    .B(\u_neuron.fst_last_t_next[7] ),
    .A_N(net376));
 sg13g2_nand2_1 _431_ (.Y(_199_),
    .A(net81),
    .B(net348));
 sg13g2_o21ai_1 _432_ (.B1(_199_),
    .Y(_037_),
    .A1(net348),
    .A2(_198_));
 sg13g2_nand2b_1 _433_ (.Y(_200_),
    .B(\u_neuron.td_curr_next[0] ),
    .A_N(net370));
 sg13g2_nand2_1 _434_ (.Y(_201_),
    .A(net156),
    .B(net339));
 sg13g2_o21ai_1 _435_ (.B1(_201_),
    .Y(_038_),
    .A1(net339),
    .A2(_200_));
 sg13g2_nand2b_1 _436_ (.Y(_202_),
    .B(\u_neuron.td_curr_next[1] ),
    .A_N(net369));
 sg13g2_nand2_1 _437_ (.Y(_203_),
    .A(net170),
    .B(net337));
 sg13g2_o21ai_1 _438_ (.B1(_203_),
    .Y(_039_),
    .A1(net337),
    .A2(_202_));
 sg13g2_nand2b_1 _439_ (.Y(_204_),
    .B(\u_neuron.td_curr_next[2] ),
    .A_N(net370));
 sg13g2_nand2_1 _440_ (.Y(_205_),
    .A(net166),
    .B(net337));
 sg13g2_o21ai_1 _441_ (.B1(_205_),
    .Y(_040_),
    .A1(net335),
    .A2(_204_));
 sg13g2_nand2b_1 _442_ (.Y(_206_),
    .B(\u_neuron.td_curr_next[3] ),
    .A_N(net369));
 sg13g2_nand2_1 _443_ (.Y(_207_),
    .A(net182),
    .B(net335));
 sg13g2_o21ai_1 _444_ (.B1(_207_),
    .Y(_041_),
    .A1(net335),
    .A2(_206_));
 sg13g2_nand2b_1 _445_ (.Y(_208_),
    .B(\u_neuron.td_curr_next[4] ),
    .A_N(net369));
 sg13g2_nand2_1 _446_ (.Y(_209_),
    .A(net178),
    .B(net334));
 sg13g2_o21ai_1 _447_ (.B1(_209_),
    .Y(_042_),
    .A1(net334),
    .A2(_208_));
 sg13g2_nand2b_1 _448_ (.Y(_210_),
    .B(\u_neuron.td_curr_next[5] ),
    .A_N(net369));
 sg13g2_nand2_1 _449_ (.Y(_211_),
    .A(net162),
    .B(net334));
 sg13g2_o21ai_1 _450_ (.B1(_211_),
    .Y(_043_),
    .A1(net334),
    .A2(_210_));
 sg13g2_nand2b_1 _451_ (.Y(_212_),
    .B(\u_neuron.td_curr_next[6] ),
    .A_N(net370));
 sg13g2_nand2_1 _452_ (.Y(_213_),
    .A(net155),
    .B(net336));
 sg13g2_o21ai_1 _453_ (.B1(_213_),
    .Y(_044_),
    .A1(net336),
    .A2(_212_));
 sg13g2_nand2b_1 _454_ (.Y(_214_),
    .B(\u_neuron.td_curr_next[7] ),
    .A_N(net370));
 sg13g2_nand2_1 _455_ (.Y(_215_),
    .A(net153),
    .B(net336));
 sg13g2_o21ai_1 _456_ (.B1(_215_),
    .Y(_045_),
    .A1(net336),
    .A2(_214_));
 sg13g2_nand2b_1 _457_ (.Y(_216_),
    .B(\u_neuron.lif_V_next[0] ),
    .A_N(net373));
 sg13g2_nand2_1 _458_ (.Y(_217_),
    .A(net142),
    .B(net342));
 sg13g2_o21ai_1 _459_ (.B1(_217_),
    .Y(_046_),
    .A1(net343),
    .A2(_216_));
 sg13g2_nand2b_1 _460_ (.Y(_218_),
    .B(\u_neuron.lif_V_next[1] ),
    .A_N(net373));
 sg13g2_nand2_1 _461_ (.Y(_219_),
    .A(net173),
    .B(net343));
 sg13g2_o21ai_1 _462_ (.B1(_219_),
    .Y(_047_),
    .A1(net343),
    .A2(_218_));
 sg13g2_nand2b_1 _463_ (.Y(_220_),
    .B(\u_neuron.lif_V_next[2] ),
    .A_N(net373));
 sg13g2_nand2_1 _464_ (.Y(_221_),
    .A(net191),
    .B(net342));
 sg13g2_o21ai_1 _465_ (.B1(_221_),
    .Y(_048_),
    .A1(net342),
    .A2(_220_));
 sg13g2_nand2b_1 _466_ (.Y(_222_),
    .B(\u_neuron.lif_V_next[3] ),
    .A_N(net371));
 sg13g2_nand2_1 _467_ (.Y(_223_),
    .A(net161),
    .B(net342));
 sg13g2_o21ai_1 _468_ (.B1(_223_),
    .Y(_049_),
    .A1(net339),
    .A2(_222_));
 sg13g2_nand2b_1 _469_ (.Y(_224_),
    .B(\u_neuron.lif_V_next[4] ),
    .A_N(net371));
 sg13g2_nand2_1 _470_ (.Y(_225_),
    .A(net199),
    .B(net339));
 sg13g2_o21ai_1 _471_ (.B1(_225_),
    .Y(_050_),
    .A1(net339),
    .A2(_224_));
 sg13g2_nand2b_1 _472_ (.Y(_226_),
    .B(\u_neuron.lif_V_next[5] ),
    .A_N(net371));
 sg13g2_nand2_1 _473_ (.Y(_227_),
    .A(net195),
    .B(net338));
 sg13g2_o21ai_1 _474_ (.B1(_227_),
    .Y(_051_),
    .A1(net337),
    .A2(_226_));
 sg13g2_nand2b_1 _475_ (.Y(_228_),
    .B(\u_neuron.lif_V_next[6] ),
    .A_N(net371));
 sg13g2_nand2_1 _476_ (.Y(_229_),
    .A(net149),
    .B(net338));
 sg13g2_o21ai_1 _477_ (.B1(_229_),
    .Y(_052_),
    .A1(net338),
    .A2(_228_));
 sg13g2_nand2b_1 _478_ (.Y(_230_),
    .B(\u_neuron.lif_V_next[7] ),
    .A_N(net371));
 sg13g2_nand2_1 _479_ (.Y(_231_),
    .A(net120),
    .B(net338));
 sg13g2_o21ai_1 _480_ (.B1(_231_),
    .Y(_053_),
    .A1(net338),
    .A2(_230_));
 sg13g2_nand3_1 _481_ (.B(net469),
    .C(\u_neuron.cfg_op[1] ),
    .A(\u_neuron.in_fire ),
    .Y(_232_));
 sg13g2_nor3_2 _482_ (.A(\u_neuron.cfg_op[0] ),
    .B(_128_),
    .C(_232_),
    .Y(_233_));
 sg13g2_mux2_1 _483_ (.A0(net209),
    .A1(\u_neuron.cfg_arg[3] ),
    .S(_233_),
    .X(_054_));
 sg13g2_nand2b_1 _484_ (.Y(_234_),
    .B(\u_neuron.conv_shift_next[0] ),
    .A_N(net374));
 sg13g2_nand2_1 _485_ (.Y(_235_),
    .A(net124),
    .B(net346));
 sg13g2_o21ai_1 _486_ (.B1(_235_),
    .Y(_055_),
    .A1(net346),
    .A2(_234_));
 sg13g2_nand2b_1 _487_ (.Y(_236_),
    .B(\u_neuron.conv_shift_next[1] ),
    .A_N(net374));
 sg13g2_nand2_1 _488_ (.Y(_237_),
    .A(net181),
    .B(net346));
 sg13g2_o21ai_1 _489_ (.B1(_237_),
    .Y(_056_),
    .A1(net346),
    .A2(_236_));
 sg13g2_nand2b_1 _490_ (.Y(_238_),
    .B(\u_neuron.conv_shift_next[2] ),
    .A_N(net372));
 sg13g2_nand2_1 _491_ (.Y(_239_),
    .A(net98),
    .B(net342));
 sg13g2_o21ai_1 _492_ (.B1(_239_),
    .Y(_057_),
    .A1(net342),
    .A2(_238_));
 sg13g2_nand2b_1 _493_ (.Y(_240_),
    .B(\u_neuron.conv_shift_next[3] ),
    .A_N(net372));
 sg13g2_nand2_1 _494_ (.Y(_241_),
    .A(net77),
    .B(net342));
 sg13g2_o21ai_1 _495_ (.B1(_241_),
    .Y(_058_),
    .A1(net342),
    .A2(_240_));
 sg13g2_nor2_1 _496_ (.A(net137),
    .B(_233_),
    .Y(_242_));
 sg13g2_a21oi_1 _497_ (.A1(\u_neuron.cfg_arg[2] ),
    .A2(_233_),
    .Y(_059_),
    .B1(net138));
 sg13g2_nand2_1 _498_ (.Y(_243_),
    .A(\u_neuron.cfg_arg[0] ),
    .B(_233_));
 sg13g2_o21ai_1 _499_ (.B1(net222),
    .Y(_060_),
    .A1(_065_),
    .A2(_233_));
 sg13g2_mux2_1 _500_ (.A0(net432),
    .A1(\u_neuron.cfg_arg[1] ),
    .S(_233_),
    .X(_061_));
 sg13g2_nand2b_1 _501_ (.Y(_244_),
    .B(\u_neuron.fst_armed_next ),
    .A_N(net377));
 sg13g2_nand2_1 _502_ (.Y(_245_),
    .A(net158),
    .B(net350));
 sg13g2_o21ai_1 _503_ (.B1(_245_),
    .Y(_062_),
    .A1(net350),
    .A2(_244_));
 sg13g2_nand2b_1 _504_ (.Y(_246_),
    .B(\u_neuron.spike_seen_this_tick_next ),
    .A_N(net375));
 sg13g2_nand2_1 _505_ (.Y(_247_),
    .A(net165),
    .B(net346));
 sg13g2_o21ai_1 _506_ (.B1(_247_),
    .Y(_063_),
    .A1(net346),
    .A2(_246_));
 sg13g2_dfrbpq_1 _507_ (.RESET_B(net449),
    .D(_003_),
    .Q(\u_neuron.conv_last_sum[0] ),
    .CLK(clknet_5_16__leaf_clk));
 sg13g2_dfrbpq_1 _508_ (.RESET_B(net449),
    .D(_004_),
    .Q(\u_neuron.conv_last_sum[1] ),
    .CLK(clknet_5_0__leaf_clk));
 sg13g2_dfrbpq_1 _509_ (.RESET_B(net449),
    .D(_005_),
    .Q(\u_neuron.conv_last_sum[2] ),
    .CLK(clknet_5_16__leaf_clk));
 sg13g2_dfrbpq_1 _510_ (.RESET_B(net439),
    .D(_006_),
    .Q(\u_neuron.td_last_diff[0] ),
    .CLK(clknet_5_1__leaf_clk));
 sg13g2_dfrbpq_1 _511_ (.RESET_B(net449),
    .D(_007_),
    .Q(\u_neuron.td_last_diff[1] ),
    .CLK(clknet_5_0__leaf_clk));
 sg13g2_dfrbpq_1 _512_ (.RESET_B(net449),
    .D(_008_),
    .Q(\u_neuron.td_last_diff[2] ),
    .CLK(clknet_5_0__leaf_clk));
 sg13g2_dfrbpq_1 _513_ (.RESET_B(net449),
    .D(_009_),
    .Q(\u_neuron.td_last_diff[3] ),
    .CLK(clknet_5_1__leaf_clk));
 sg13g2_dfrbpq_1 _514_ (.RESET_B(net439),
    .D(_010_),
    .Q(\u_neuron.td_last_diff[4] ),
    .CLK(clknet_5_4__leaf_clk));
 sg13g2_dfrbpq_1 _515_ (.RESET_B(net438),
    .D(_011_),
    .Q(\u_neuron.td_last_diff[5] ),
    .CLK(clknet_5_1__leaf_clk));
 sg13g2_dfrbpq_1 _516_ (.RESET_B(net439),
    .D(_012_),
    .Q(\u_neuron.td_last_diff[6] ),
    .CLK(clknet_5_4__leaf_clk));
 sg13g2_dfrbpq_1 _517_ (.RESET_B(net439),
    .D(net65),
    .Q(\u_neuron.td_last_diff[7] ),
    .CLK(clknet_5_0__leaf_clk));
 sg13g2_dfrbpq_2 _518_ (.RESET_B(net452),
    .D(_014_),
    .Q(\u_neuron.fst_t[0] ),
    .CLK(clknet_5_20__leaf_clk));
 sg13g2_dfrbpq_2 _519_ (.RESET_B(net452),
    .D(_015_),
    .Q(\u_neuron.fst_t[1] ),
    .CLK(clknet_5_21__leaf_clk));
 sg13g2_dfrbpq_2 _520_ (.RESET_B(net451),
    .D(_016_),
    .Q(\u_neuron.fst_t[2] ),
    .CLK(clknet_5_19__leaf_clk));
 sg13g2_dfrbpq_2 _521_ (.RESET_B(net451),
    .D(_017_),
    .Q(\u_neuron.fst_t[3] ),
    .CLK(clknet_5_17__leaf_clk));
 sg13g2_dfrbpq_2 _522_ (.RESET_B(net449),
    .D(_018_),
    .Q(\u_neuron.fst_t[4] ),
    .CLK(clknet_5_17__leaf_clk));
 sg13g2_dfrbpq_2 _523_ (.RESET_B(net451),
    .D(net117),
    .Q(\u_neuron.fst_t[5] ),
    .CLK(clknet_5_17__leaf_clk));
 sg13g2_dfrbpq_1 _524_ (.RESET_B(net451),
    .D(_020_),
    .Q(\u_neuron.fst_t[6] ),
    .CLK(clknet_5_20__leaf_clk));
 sg13g2_dfrbpq_1 _525_ (.RESET_B(net451),
    .D(net134),
    .Q(\u_neuron.fst_t[7] ),
    .CLK(clknet_5_20__leaf_clk));
 sg13g2_dfrbpq_2 _526_ (.RESET_B(net438),
    .D(net127),
    .Q(\u_neuron.td_prev[0] ),
    .CLK(clknet_5_4__leaf_clk));
 sg13g2_dfrbpq_2 _527_ (.RESET_B(net437),
    .D(net115),
    .Q(\u_neuron.td_prev[1] ),
    .CLK(clknet_5_12__leaf_clk));
 sg13g2_dfrbpq_2 _528_ (.RESET_B(net437),
    .D(net119),
    .Q(\u_neuron.td_prev[2] ),
    .CLK(clknet_5_9__leaf_clk));
 sg13g2_dfrbpq_2 _529_ (.RESET_B(net436),
    .D(net141),
    .Q(\u_neuron.td_prev[3] ),
    .CLK(clknet_5_2__leaf_clk));
 sg13g2_dfrbpq_2 _530_ (.RESET_B(net436),
    .D(net152),
    .Q(\u_neuron.td_prev[4] ),
    .CLK(clknet_5_2__leaf_clk));
 sg13g2_dfrbpq_2 _531_ (.RESET_B(net436),
    .D(net145),
    .Q(\u_neuron.td_prev[5] ),
    .CLK(clknet_5_2__leaf_clk));
 sg13g2_dfrbpq_1 _532_ (.RESET_B(net438),
    .D(net113),
    .Q(\u_neuron.td_prev[6] ),
    .CLK(clknet_5_3__leaf_clk));
 sg13g2_dfrbpq_1 _533_ (.RESET_B(net438),
    .D(net132),
    .Q(\u_neuron.td_prev[7] ),
    .CLK(clknet_5_0__leaf_clk));
 sg13g2_dfrbpq_1 _534_ (.RESET_B(net452),
    .D(net60),
    .Q(\u_neuron.fst_last_t[0] ),
    .CLK(clknet_5_20__leaf_clk));
 sg13g2_dfrbpq_1 _535_ (.RESET_B(net451),
    .D(net110),
    .Q(\u_neuron.fst_last_t[1] ),
    .CLK(clknet_5_19__leaf_clk));
 sg13g2_dfrbpq_1 _536_ (.RESET_B(net451),
    .D(net105),
    .Q(\u_neuron.fst_last_t[2] ),
    .CLK(clknet_5_19__leaf_clk));
 sg13g2_dfrbpq_1 _537_ (.RESET_B(net449),
    .D(net89),
    .Q(\u_neuron.fst_last_t[3] ),
    .CLK(clknet_5_17__leaf_clk));
 sg13g2_dfrbpq_1 _538_ (.RESET_B(net450),
    .D(net63),
    .Q(\u_neuron.fst_last_t[4] ),
    .CLK(clknet_5_16__leaf_clk));
 sg13g2_dfrbpq_1 _539_ (.RESET_B(net451),
    .D(net67),
    .Q(\u_neuron.fst_last_t[5] ),
    .CLK(clknet_5_19__leaf_clk));
 sg13g2_dfrbpq_1 _540_ (.RESET_B(net452),
    .D(net74),
    .Q(\u_neuron.fst_last_t[6] ),
    .CLK(clknet_5_21__leaf_clk));
 sg13g2_dfrbpq_1 _541_ (.RESET_B(net452),
    .D(net82),
    .Q(\u_neuron.fst_last_t[7] ),
    .CLK(clknet_5_21__leaf_clk));
 sg13g2_dfrbpq_2 _542_ (.RESET_B(net438),
    .D(net157),
    .Q(\u_neuron.td_curr[0] ),
    .CLK(clknet_5_3__leaf_clk));
 sg13g2_dfrbpq_2 _543_ (.RESET_B(net437),
    .D(_039_),
    .Q(\u_neuron.td_curr[1] ),
    .CLK(clknet_5_12__leaf_clk));
 sg13g2_dfrbpq_2 _544_ (.RESET_B(net436),
    .D(_040_),
    .Q(\u_neuron.td_curr[2] ),
    .CLK(clknet_5_9__leaf_clk));
 sg13g2_dfrbpq_2 _545_ (.RESET_B(net436),
    .D(_041_),
    .Q(\u_neuron.td_curr[3] ),
    .CLK(clknet_5_2__leaf_clk));
 sg13g2_dfrbpq_2 _546_ (.RESET_B(net436),
    .D(_042_),
    .Q(\u_neuron.td_curr[4] ),
    .CLK(clknet_5_2__leaf_clk));
 sg13g2_dfrbpq_2 _547_ (.RESET_B(net436),
    .D(_043_),
    .Q(\u_neuron.td_curr[5] ),
    .CLK(clknet_5_3__leaf_clk));
 sg13g2_dfrbpq_2 _548_ (.RESET_B(net436),
    .D(_044_),
    .Q(\u_neuron.td_curr[6] ),
    .CLK(clknet_5_3__leaf_clk));
 sg13g2_dfrbpq_2 _549_ (.RESET_B(net438),
    .D(net154),
    .Q(\u_neuron.td_curr[7] ),
    .CLK(clknet_5_3__leaf_clk));
 sg13g2_dfrbpq_2 _550_ (.RESET_B(net440),
    .D(net143),
    .Q(\u_neuron.lif_V[0] ),
    .CLK(clknet_5_5__leaf_clk));
 sg13g2_dfrbpq_2 _551_ (.RESET_B(net450),
    .D(_047_),
    .Q(\u_neuron.lif_V[1] ),
    .CLK(clknet_5_5__leaf_clk));
 sg13g2_dfrbpq_2 _552_ (.RESET_B(net440),
    .D(_048_),
    .Q(\u_neuron.lif_V[2] ),
    .CLK(clknet_5_5__leaf_clk));
 sg13g2_dfrbpq_2 _553_ (.RESET_B(net440),
    .D(_049_),
    .Q(\u_neuron.lif_V[3] ),
    .CLK(clknet_5_5__leaf_clk));
 sg13g2_dfrbpq_2 _554_ (.RESET_B(net437),
    .D(_050_),
    .Q(\u_neuron.lif_V[4] ),
    .CLK(clknet_5_4__leaf_clk));
 sg13g2_dfrbpq_2 _555_ (.RESET_B(net437),
    .D(_051_),
    .Q(\u_neuron.lif_V[5] ),
    .CLK(clknet_5_7__leaf_clk));
 sg13g2_dfrbpq_2 _556_ (.RESET_B(net437),
    .D(net150),
    .Q(\u_neuron.lif_V[6] ),
    .CLK(clknet_5_13__leaf_clk));
 sg13g2_dfrbpq_2 _557_ (.RESET_B(net437),
    .D(net121),
    .Q(\u_neuron.lif_V[7] ),
    .CLK(clknet_5_6__leaf_clk));
 sg13g2_dfrbpq_2 _558_ (.RESET_B(net450),
    .D(net210),
    .Q(\u_neuron.learn_en ),
    .CLK(clknet_5_7__leaf_clk));
 sg13g2_dfrbpq_2 _559_ (.RESET_B(net450),
    .D(net125),
    .Q(\u_neuron.conv_shift[0] ),
    .CLK(clknet_5_0__leaf_clk));
 sg13g2_dfrbpq_2 _560_ (.RESET_B(net455),
    .D(_056_),
    .Q(\u_neuron.conv_shift[1] ),
    .CLK(clknet_5_16__leaf_clk));
 sg13g2_dfrbpq_1 _561_ (.RESET_B(net438),
    .D(net99),
    .Q(\u_neuron.conv_shift[2] ),
    .CLK(clknet_5_1__leaf_clk));
 sg13g2_dfrbpq_1 _562_ (.RESET_B(net438),
    .D(net78),
    .Q(\u_neuron.conv_shift[3] ),
    .CLK(clknet_5_1__leaf_clk));
 sg13g2_dfrbpq_1 _563_ (.RESET_B(net450),
    .D(net139),
    .Q(_002_),
    .CLK(clknet_5_7__leaf_clk));
 sg13g2_dfrbpq_1 _564_ (.RESET_B(net450),
    .D(net223),
    .Q(\u_neuron.mode[0] ),
    .CLK(clknet_5_7__leaf_clk));
 sg13g2_dfrbpq_2 _565_ (.RESET_B(net454),
    .D(net232),
    .Q(\u_neuron.mode[1] ),
    .CLK(clknet_5_7__leaf_clk));
 sg13g2_dfrbpq_2 _566_ (.RESET_B(net450),
    .D(_062_),
    .Q(\u_neuron.fst_armed ),
    .CLK(clknet_5_17__leaf_clk));
 sg13g2_dfrbpq_2 _567_ (.RESET_B(net455),
    .D(_063_),
    .Q(\u_neuron.spike_seen_this_tick ),
    .CLK(clknet_5_16__leaf_clk));
 sg13g2_inv_2 \u_neuron.u_conv/_08_  (.Y(\u_neuron.u_conv/_00_ ),
    .A(net124));
 sg13g2_and3_2 \u_neuron.u_conv/_09_  (.X(\u_neuron.conv_emit_data[2] ),
    .A(\u_neuron.conv_shift[1] ),
    .B(\u_neuron.spike_seen_this_tick ),
    .C(net236));
 sg13g2_nor2_1 \u_neuron.u_conv/_10_  (.A(\u_neuron.conv_shift[1] ),
    .B(\u_neuron.spike_seen_this_tick ),
    .Y(\u_neuron.u_conv/_01_ ));
 sg13g2_xor2_1 \u_neuron.u_conv/_11_  (.B(net237),
    .A(\u_neuron.conv_shift[1] ),
    .X(\u_neuron.conv_emit_data[0] ));
 sg13g2_a21oi_1 \u_neuron.u_conv/_12_  (.A1(\u_neuron.conv_shift[1] ),
    .A2(\u_neuron.spike_seen_this_tick ),
    .Y(\u_neuron.u_conv/_02_ ),
    .B1(net236));
 sg13g2_nor2_1 \u_neuron.u_conv/_13_  (.A(\u_neuron.conv_emit_data[2] ),
    .B(\u_neuron.u_conv/_02_ ),
    .Y(\u_neuron.conv_emit_data[1] ));
 sg13g2_nand2_1 \u_neuron.u_conv/_14_  (.Y(\u_neuron.u_conv/_03_ ),
    .A(net385),
    .B(\u_neuron.mode_conv_evt ));
 sg13g2_nor4_1 \u_neuron.u_conv/_15_  (.A(\u_neuron.u_conv/_00_ ),
    .B(net417),
    .C(\u_neuron.u_conv/_01_ ),
    .D(net325),
    .Y(\u_neuron.conv_post_spike ));
 sg13g2_inv_1 \u_neuron.u_conv/_16_  (.Y(\u_neuron.conv_emit_data[6] ),
    .A(\u_neuron.conv_post_spike ));
 sg13g2_nor2_1 \u_neuron.u_conv/_17_  (.A(net417),
    .B(net325),
    .Y(\u_neuron.u_conv/_04_ ));
 sg13g2_a21o_1 \u_neuron.u_conv/_18_  (.A2(\u_neuron.u_conv/_04_ ),
    .A1(\u_neuron.stream_act ),
    .B1(\u_neuron.conv_post_spike ),
    .X(\u_neuron.conv_emit_valid ));
 sg13g2_nor2_1 \u_neuron.u_conv/_19_  (.A(\u_neuron.spike_seen_this_tick ),
    .B(net324),
    .Y(\u_neuron.u_conv/_05_ ));
 sg13g2_a21oi_1 \u_neuron.u_conv/_20_  (.A1(\u_neuron.u_conv/_00_ ),
    .A2(net324),
    .Y(\u_neuron.conv_shift_next[0] ),
    .B1(\u_neuron.u_conv/_05_ ));
 sg13g2_nand2_1 \u_neuron.u_conv/_21_  (.Y(\u_neuron.u_conv/_06_ ),
    .A(net181),
    .B(net324));
 sg13g2_o21ai_1 \u_neuron.u_conv/_22_  (.B1(\u_neuron.u_conv/_06_ ),
    .Y(\u_neuron.conv_shift_next[1] ),
    .A1(\u_neuron.u_conv/_00_ ),
    .A2(net324));
 sg13g2_mux2_1 \u_neuron.u_conv/_23_  (.A0(\u_neuron.conv_shift[1] ),
    .A1(net98),
    .S(net324),
    .X(\u_neuron.conv_shift_next[2] ));
 sg13g2_mux2_1 \u_neuron.u_conv/_24_  (.A0(\u_neuron.conv_shift[2] ),
    .A1(net77),
    .S(net324),
    .X(\u_neuron.conv_shift_next[3] ));
 sg13g2_mux2_1 \u_neuron.u_conv/_25_  (.A0(\u_neuron.conv_emit_data[0] ),
    .A1(net76),
    .S(net324),
    .X(\u_neuron.conv_last_sum_next[0] ));
 sg13g2_mux2_1 \u_neuron.u_conv/_26_  (.A0(\u_neuron.conv_emit_data[1] ),
    .A1(net83),
    .S(net325),
    .X(\u_neuron.conv_last_sum_next[1] ));
 sg13g2_mux2_1 \u_neuron.u_conv/_27_  (.A0(\u_neuron.conv_emit_data[2] ),
    .A1(net72),
    .S(net324),
    .X(\u_neuron.conv_last_sum_next[2] ));
 sg13g2_o21ai_1 \u_neuron.u_conv/_28_  (.B1(net325),
    .Y(\u_neuron.u_conv/_07_ ),
    .A1(net165),
    .A2(\u_neuron.mode_conv_evt ));
 sg13g2_inv_1 \u_neuron.u_conv/_29_  (.Y(\u_neuron.spike_seen_this_tick_next ),
    .A(\u_neuron.u_conv/_07_ ));
 sg13g2_tiehi tt_um_crockpotveggies_neuron_38 (.L_HI(net38));
 sg13g2_tielo \u_neuron.u_mode_sel/_07__18  (.L_LO(net18));
 sg13g2_tielo \u_neuron.u_mode_sel/_00__19  (.L_LO(net19));
 sg13g2_tielo tt_um_crockpotveggies_neuron_20 (.L_LO(net20));
 sg13g2_buf_1 \u_neuron.u_conv/_34_  (.A(\u_neuron.conv_emit_data[6] ),
    .X(\u_neuron.conv_emit_data[4] ));
 sg13g2_inv_1 \u_neuron.u_decode/_04_  (.Y(\u_neuron.u_decode/_00_ ),
    .A(\u_neuron.in_data[0] ));
 sg13g2_nand4_1 \u_neuron.u_decode/_05_  (.B(\u_neuron.in_data[2] ),
    .C(\u_neuron.in_data[5] ),
    .A(\u_neuron.in_data[3] ),
    .Y(\u_neuron.u_decode/_01_ ),
    .D(\u_neuron.in_data[4] ));
 sg13g2_nor4_1 \u_neuron.u_decode/_06_  (.A(\u_neuron.in_data[7] ),
    .B(\u_neuron.in_data[1] ),
    .C(\u_neuron.u_decode/_00_ ),
    .D(\u_neuron.u_decode/_01_ ),
    .Y(\u_neuron.is_reset_cmd ));
 sg13g2_nor2b_1 \u_neuron.u_decode/_07_  (.A(\u_neuron.in_data[7] ),
    .B_N(\u_neuron.in_data[1] ),
    .Y(\u_neuron.u_decode/_02_ ));
 sg13g2_nand2b_1 \u_neuron.u_decode/_08_  (.Y(\u_neuron.u_decode/_03_ ),
    .B(\u_neuron.u_decode/_02_ ),
    .A_N(\u_neuron.u_decode/_01_ ));
 sg13g2_nor2_1 \u_neuron.u_decode/_09_  (.A(\u_neuron.in_data[0] ),
    .B(\u_neuron.u_decode/_03_ ),
    .Y(\u_neuron.is_arm_cmd ));
 sg13g2_nor2_1 \u_neuron.u_decode/_10_  (.A(\u_neuron.u_decode/_00_ ),
    .B(\u_neuron.u_decode/_03_ ),
    .Y(\u_neuron.is_cfg_cmd ));
 sg13g2_nand2b_1 \u_neuron.u_decode/_11_  (.Y(\u_neuron.is_special_cmd ),
    .B(\u_neuron.u_decode/_03_ ),
    .A_N(net378));
 sg13g2_buf_8 \u_neuron.u_decode/_12_  (.A(\u_neuron.in_data[0] ),
    .X(\u_neuron.addr[0] ));
 sg13g2_buf_1 \u_neuron.u_decode/_13_  (.A(\u_neuron.in_data[1] ),
    .X(\u_neuron.addr[1] ));
 sg13g2_buf_1 \u_neuron.u_decode/_14_  (.A(\u_neuron.in_data[2] ),
    .X(\u_neuron.addr[2] ));
 sg13g2_buf_1 \u_neuron.u_decode/_15_  (.A(\u_neuron.in_data[3] ),
    .X(\u_neuron.addr[3] ));
 sg13g2_buf_1 \u_neuron.u_decode/_16_  (.A(\u_neuron.in_data[4] ),
    .X(\u_neuron.addr[4] ));
 sg13g2_buf_1 \u_neuron.u_decode/_17_  (.A(\u_neuron.in_data[5] ),
    .X(\u_neuron.addr[5] ));
 sg13g2_buf_8 \u_neuron.u_decode/_18_  (.A(net221),
    .X(\u_neuron.cfg_arg[0] ));
 sg13g2_buf_8 \u_neuron.u_decode/_19_  (.A(net228),
    .X(\u_neuron.cfg_arg[1] ));
 sg13g2_buf_1 \u_neuron.u_decode/_20_  (.A(net219),
    .X(\u_neuron.cfg_arg[2] ));
 sg13g2_buf_1 \u_neuron.u_decode/_21_  (.A(\u_neuron.uio_in_sync[7] ),
    .X(\u_neuron.cfg_arg[3] ));
 sg13g2_buf_1 \u_neuron.u_decode/_22_  (.A(\u_neuron.uio_in_sync[2] ),
    .X(\u_neuron.cfg_op[0] ));
 sg13g2_buf_1 \u_neuron.u_decode/_23_  (.A(\u_neuron.uio_in_sync[3] ),
    .X(\u_neuron.cfg_op[1] ));
 sg13g2_buf_2 \u_neuron.u_decode/_24_  (.A(\u_neuron.in_data[7] ),
    .X(\u_neuron.is_tick ));
 sg13g2_buf_1 \u_neuron.u_decode/_25_  (.A(\u_neuron.in_data[6] ),
    .X(\u_neuron.polarity ));
 sg13g2_nand2b_2 \u_neuron.u_frontend/_04_  (.Y(\u_neuron.u_frontend/_01_ ),
    .B(\u_neuron.u_frontend/in_req ),
    .A_N(net417));
 sg13g2_nand3b_1 \u_neuron.u_frontend/_05_  (.B(net469),
    .C(net458),
    .Y(\u_neuron.u_frontend/_02_ ),
    .A_N(net69));
 sg13g2_nor2_2 \u_neuron.u_frontend/_06_  (.A(\u_neuron.u_frontend/_01_ ),
    .B(\u_neuron.u_frontend/_02_ ),
    .Y(\u_neuron.in_fire ));
 sg13g2_and2_1 \u_neuron.u_frontend/_07_  (.A(net417),
    .B(\u_neuron.u_frontend/out_ack ),
    .X(\u_neuron.out_fire ));
 sg13g2_nand2_1 \u_neuron.u_frontend/_08_  (.Y(\u_neuron.u_frontend/_03_ ),
    .A(\u_neuron.u_frontend/in_req ),
    .B(net69));
 sg13g2_o21ai_1 \u_neuron.u_frontend/_09_  (.B1(net70),
    .Y(\u_neuron.u_frontend/_00_ ),
    .A1(\u_neuron.u_frontend/_01_ ),
    .A2(\u_neuron.u_frontend/_02_ ));
 sg13g2_nor2_1 \u_neuron.u_frontend/_10_  (.A(\u_neuron.u_frontend/_01_ ),
    .B(\u_neuron.u_frontend/_02_ ),
    .Y(\u_neuron.in_ack ));
 sg13g2_dfrbpq_2 \u_neuron.u_frontend/_11_  (.RESET_B(net462),
    .D(net53),
    .Q(\u_neuron.in_data[0] ),
    .CLK(clknet_5_25__leaf_clk));
 sg13g2_dfrbpq_2 \u_neuron.u_frontend/_12_  (.RESET_B(net462),
    .D(net54),
    .Q(\u_neuron.in_data[1] ),
    .CLK(clknet_5_31__leaf_clk));
 sg13g2_dfrbpq_1 \u_neuron.u_frontend/_13_  (.RESET_B(net461),
    .D(net46),
    .Q(\u_neuron.in_data[2] ),
    .CLK(clknet_5_24__leaf_clk));
 sg13g2_dfrbpq_1 \u_neuron.u_frontend/_14_  (.RESET_B(net461),
    .D(net49),
    .Q(\u_neuron.in_data[3] ),
    .CLK(clknet_5_24__leaf_clk));
 sg13g2_dfrbpq_1 \u_neuron.u_frontend/_15_  (.RESET_B(net461),
    .D(net51),
    .Q(\u_neuron.in_data[4] ),
    .CLK(clknet_5_24__leaf_clk));
 sg13g2_dfrbpq_1 \u_neuron.u_frontend/_16_  (.RESET_B(net462),
    .D(net52),
    .Q(\u_neuron.in_data[5] ),
    .CLK(clknet_5_24__leaf_clk));
 sg13g2_dfrbpq_1 \u_neuron.u_frontend/_17_  (.RESET_B(net461),
    .D(net48),
    .Q(\u_neuron.in_data[6] ),
    .CLK(clknet_5_25__leaf_clk));
 sg13g2_dfrbpq_2 \u_neuron.u_frontend/_18_  (.RESET_B(net462),
    .D(net55),
    .Q(\u_neuron.in_data[7] ),
    .CLK(clknet_5_31__leaf_clk));
 sg13g2_dfrbpq_2 \u_neuron.u_frontend/_19_  (.RESET_B(net458),
    .D(net56),
    .Q(\u_neuron.u_frontend/in_req ),
    .CLK(clknet_5_23__leaf_clk));
 sg13g2_dfrbpq_1 \u_neuron.u_frontend/_20_  (.RESET_B(net458),
    .D(net57),
    .Q(\u_neuron.u_frontend/out_ack ),
    .CLK(clknet_5_23__leaf_clk));
 sg13g2_dfrbpq_1 \u_neuron.u_frontend/_21_  (.RESET_B(net459),
    .D(net47),
    .Q(\u_neuron.uio_in_sync[2] ),
    .CLK(clknet_5_29__leaf_clk));
 sg13g2_dfrbpq_1 \u_neuron.u_frontend/_22_  (.RESET_B(net459),
    .D(net50),
    .Q(\u_neuron.uio_in_sync[3] ),
    .CLK(clknet_5_29__leaf_clk));
 sg13g2_dfrbpq_1 \u_neuron.u_frontend/_23_  (.RESET_B(net459),
    .D(net58),
    .Q(\u_neuron.uio_in_sync[4] ),
    .CLK(clknet_5_31__leaf_clk));
 sg13g2_dfrbpq_1 \u_neuron.u_frontend/_24_  (.RESET_B(net459),
    .D(net45),
    .Q(\u_neuron.uio_in_sync[5] ),
    .CLK(clknet_5_29__leaf_clk));
 sg13g2_dfrbpq_1 \u_neuron.u_frontend/_25_  (.RESET_B(net460),
    .D(net43),
    .Q(\u_neuron.uio_in_sync[6] ),
    .CLK(clknet_5_28__leaf_clk));
 sg13g2_dfrbpq_1 \u_neuron.u_frontend/_26_  (.RESET_B(net460),
    .D(net44),
    .Q(\u_neuron.uio_in_sync[7] ),
    .CLK(clknet_5_28__leaf_clk));
 sg13g2_dfrbpq_1 \u_neuron.u_frontend/_27_  (.RESET_B(net461),
    .D(net1),
    .Q(\u_neuron.u_frontend/ui_in_meta[0] ),
    .CLK(clknet_5_25__leaf_clk));
 sg13g2_dfrbpq_1 \u_neuron.u_frontend/_28_  (.RESET_B(net462),
    .D(net2),
    .Q(\u_neuron.u_frontend/ui_in_meta[1] ),
    .CLK(clknet_5_31__leaf_clk));
 sg13g2_dfrbpq_1 \u_neuron.u_frontend/_29_  (.RESET_B(net461),
    .D(net3),
    .Q(\u_neuron.u_frontend/ui_in_meta[2] ),
    .CLK(clknet_5_25__leaf_clk));
 sg13g2_dfrbpq_1 \u_neuron.u_frontend/_30_  (.RESET_B(net461),
    .D(net4),
    .Q(\u_neuron.u_frontend/ui_in_meta[3] ),
    .CLK(clknet_5_27__leaf_clk));
 sg13g2_dfrbpq_1 \u_neuron.u_frontend/_31_  (.RESET_B(net461),
    .D(net5),
    .Q(\u_neuron.u_frontend/ui_in_meta[4] ),
    .CLK(clknet_5_27__leaf_clk));
 sg13g2_dfrbpq_1 \u_neuron.u_frontend/_32_  (.RESET_B(net462),
    .D(net6),
    .Q(\u_neuron.u_frontend/ui_in_meta[5] ),
    .CLK(clknet_5_31__leaf_clk));
 sg13g2_dfrbpq_1 \u_neuron.u_frontend/_33_  (.RESET_B(net462),
    .D(net7),
    .Q(\u_neuron.u_frontend/ui_in_meta[6] ),
    .CLK(clknet_5_25__leaf_clk));
 sg13g2_dfrbpq_1 \u_neuron.u_frontend/_34_  (.RESET_B(net459),
    .D(net8),
    .Q(\u_neuron.u_frontend/ui_in_meta[7] ),
    .CLK(clknet_5_29__leaf_clk));
 sg13g2_dfrbpq_1 \u_neuron.u_frontend/_35_  (.RESET_B(net453),
    .D(net9),
    .Q(\u_neuron.u_frontend/uio_in_meta[0] ),
    .CLK(clknet_5_21__leaf_clk));
 sg13g2_dfrbpq_1 \u_neuron.u_frontend/_36_  (.RESET_B(net458),
    .D(net10),
    .Q(\u_neuron.u_frontend/uio_in_meta[1] ),
    .CLK(clknet_5_23__leaf_clk));
 sg13g2_dfrbpq_1 \u_neuron.u_frontend/_37_  (.RESET_B(net459),
    .D(net11),
    .Q(\u_neuron.u_frontend/uio_in_meta[2] ),
    .CLK(clknet_5_22__leaf_clk));
 sg13g2_dfrbpq_1 \u_neuron.u_frontend/_38_  (.RESET_B(net458),
    .D(net12),
    .Q(\u_neuron.u_frontend/uio_in_meta[3] ),
    .CLK(clknet_5_22__leaf_clk));
 sg13g2_dfrbpq_1 \u_neuron.u_frontend/_39_  (.RESET_B(net459),
    .D(net13),
    .Q(\u_neuron.u_frontend/uio_in_meta[4] ),
    .CLK(clknet_5_29__leaf_clk));
 sg13g2_dfrbpq_1 \u_neuron.u_frontend/_40_  (.RESET_B(net458),
    .D(net14),
    .Q(\u_neuron.u_frontend/uio_in_meta[5] ),
    .CLK(clknet_5_23__leaf_clk));
 sg13g2_dfrbpq_1 \u_neuron.u_frontend/_41_  (.RESET_B(net458),
    .D(net15),
    .Q(\u_neuron.u_frontend/uio_in_meta[6] ),
    .CLK(clknet_5_22__leaf_clk));
 sg13g2_dfrbpq_1 \u_neuron.u_frontend/_42_  (.RESET_B(net458),
    .D(net16),
    .Q(\u_neuron.u_frontend/uio_in_meta[7] ),
    .CLK(clknet_5_22__leaf_clk));
 sg13g2_dfrbpq_1 \u_neuron.u_frontend/_43_  (.RESET_B(net454),
    .D(net71),
    .Q(\u_neuron.in_req_seen ),
    .CLK(clknet_5_18__leaf_clk));
 sg13g2_tiehi tt_um_crockpotveggies_neuron_39 (.L_HI(net39));
 sg13g2_tiehi \u_neuron.u_mode_sel/_09__40  (.L_HI(net40));
 sg13g2_tielo tt_um_crockpotveggies_neuron_21 (.L_LO(net21));
 sg13g2_tielo tt_um_crockpotveggies_neuron_22 (.L_LO(net22));
 sg13g2_tielo tt_um_crockpotveggies_neuron_23 (.L_LO(net23));
 sg13g2_tielo tt_um_crockpotveggies_neuron_24 (.L_LO(net24));
 sg13g2_tielo tt_um_crockpotveggies_neuron_25 (.L_LO(net25));
 sg13g2_tielo tt_um_crockpotveggies_neuron_26 (.L_LO(net26));
 sg13g2_tielo tt_um_crockpotveggies_neuron_27 (.L_LO(net27));
 sg13g2_tielo tt_um_crockpotveggies_neuron_28 (.L_LO(net28));
 sg13g2_tielo tt_um_crockpotveggies_neuron_29 (.L_LO(net29));
 sg13g2_tielo tt_um_crockpotveggies_neuron_30 (.L_LO(net30));
 sg13g2_tielo tt_um_crockpotveggies_neuron_31 (.L_LO(net31));
 sg13g2_tielo \u_neuron.u_mode_sel/_07__32  (.L_LO(net32));
 sg13g2_buf_1 \u_neuron.u_frontend/_58_  (.A(net418),
    .X(\u_neuron.out_req ));
 sg13g2_buf_1 \u_neuron.u_frontend/_59_  (.A(\u_neuron.u_frontend/in_req ),
    .X(\u_neuron.uio_in_sync[0] ));
 sg13g2_buf_1 \u_neuron.u_frontend/_60_  (.A(\u_neuron.u_frontend/out_ack ),
    .X(\u_neuron.uio_in_sync[1] ));
 sg13g2_buf_1 \u_neuron.u_frontend/_61_  (.A(\u_neuron.in_ack ),
    .X(uio_out[0]));
 sg13g2_buf_1 \u_neuron.u_frontend/_62_  (.A(net418),
    .X(uio_out[1]));
 sg13g2_inv_2 \u_neuron.u_fst/_048_  (.Y(\u_neuron.u_fst/_010_ ),
    .A(net158));
 sg13g2_inv_1 \u_neuron.u_fst/_049_  (.Y(\u_neuron.u_fst/_011_ ),
    .A(net192));
 sg13g2_inv_2 \u_neuron.u_fst/_050_  (.Y(\u_neuron.u_fst/_012_ ),
    .A(net123));
 sg13g2_inv_1 \u_neuron.u_fst/_051_  (.Y(\u_neuron.u_fst/_013_ ),
    .A(net135));
 sg13g2_inv_1 \u_neuron.u_fst/_052_  (.Y(\u_neuron.u_fst/_014_ ),
    .A(\u_neuron.fst_t[6] ));
 sg13g2_inv_1 \u_neuron.u_fst/_053_  (.Y(\u_neuron.u_fst/_015_ ),
    .A(net133));
 sg13g2_inv_2 \u_neuron.u_fst/_054_  (.Y(\u_neuron.u_fst/_016_ ),
    .A(\u_neuron.arm_event ));
 sg13g2_inv_1 \u_neuron.u_fst/_055_  (.Y(\u_neuron.u_fst/_017_ ),
    .A(net59));
 sg13g2_nor2b_1 \u_neuron.u_fst/_056_  (.A(net385),
    .B_N(\u_neuron.mode_fst_evt ),
    .Y(\u_neuron.u_fst/_018_ ));
 sg13g2_nand3b_1 \u_neuron.u_fst/_057_  (.B(\u_neuron.mode_fst_evt ),
    .C(\u_neuron.fst_armed ),
    .Y(\u_neuron.u_fst/_019_ ),
    .A_N(net385));
 sg13g2_or2_1 \u_neuron.u_fst/_058_  (.X(\u_neuron.fst_emit_data[6] ),
    .B(net323),
    .A(net417));
 sg13g2_inv_4 \u_neuron.u_fst/_059_  (.A(\u_neuron.fst_emit_data[6] ),
    .Y(\u_neuron.fst_post_spike ));
 sg13g2_and2_1 \u_neuron.u_fst/_060_  (.A(net385),
    .B(\u_neuron.mode_fst_evt ),
    .X(\u_neuron.u_fst/_020_ ));
 sg13g2_nand2_1 \u_neuron.u_fst/_061_  (.Y(\u_neuron.u_fst/_021_ ),
    .A(\u_neuron.stream_act ),
    .B(\u_neuron.u_fst/_020_ ));
 sg13g2_a21oi_1 \u_neuron.u_fst/_062_  (.A1(net323),
    .A2(\u_neuron.u_fst/_021_ ),
    .Y(\u_neuron.fst_emit_valid ),
    .B1(net417));
 sg13g2_nand2_1 \u_neuron.u_fst/_063_  (.Y(\u_neuron.u_fst/_022_ ),
    .A(net116),
    .B(\u_neuron.fst_t[4] ));
 sg13g2_and4_1 \u_neuron.u_fst/_064_  (.A(\u_neuron.fst_t[5] ),
    .B(\u_neuron.fst_t[4] ),
    .C(\u_neuron.fst_t[6] ),
    .D(\u_neuron.fst_t[7] ),
    .X(\u_neuron.u_fst/_023_ ));
 sg13g2_nand2_1 \u_neuron.u_fst/_065_  (.Y(\u_neuron.u_fst/_024_ ),
    .A(\u_neuron.fst_t[1] ),
    .B(net435));
 sg13g2_nand3_1 \u_neuron.u_fst/_066_  (.B(net435),
    .C(\u_neuron.fst_t[2] ),
    .A(\u_neuron.fst_t[1] ),
    .Y(\u_neuron.u_fst/_025_ ));
 sg13g2_and4_1 \u_neuron.u_fst/_067_  (.A(\u_neuron.fst_t[1] ),
    .B(net435),
    .C(\u_neuron.fst_t[3] ),
    .D(\u_neuron.fst_t[2] ),
    .X(\u_neuron.u_fst/_026_ ));
 sg13g2_nand4_1 \u_neuron.u_fst/_068_  (.B(net435),
    .C(\u_neuron.fst_t[3] ),
    .A(\u_neuron.fst_t[1] ),
    .Y(\u_neuron.u_fst/_027_ ),
    .D(\u_neuron.fst_t[2] ));
 sg13g2_a21oi_1 \u_neuron.u_fst/_069_  (.A1(\u_neuron.u_fst/_023_ ),
    .A2(\u_neuron.u_fst/_026_ ),
    .Y(\u_neuron.u_fst/_028_ ),
    .B1(\u_neuron.u_fst/_010_ ));
 sg13g2_nand3_1 \u_neuron.u_fst/_070_  (.B(\u_neuron.mode_fst_evt ),
    .C(\u_neuron.fst_armed ),
    .A(net385),
    .Y(\u_neuron.u_fst/_029_ ));
 sg13g2_a21oi_1 \u_neuron.u_fst/_071_  (.A1(\u_neuron.u_fst/_023_ ),
    .A2(\u_neuron.u_fst/_026_ ),
    .Y(\u_neuron.u_fst/_030_ ),
    .B1(\u_neuron.u_fst/_029_ ));
 sg13g2_mux2_1 \u_neuron.u_fst/_072_  (.A0(\u_neuron.u_fst/_029_ ),
    .A1(\u_neuron.u_fst/_030_ ),
    .S(net130),
    .X(\u_neuron.u_fst/_031_ ));
 sg13g2_nor2_1 \u_neuron.u_fst/_073_  (.A(\u_neuron.arm_event ),
    .B(\u_neuron.u_fst/_031_ ),
    .Y(\u_neuron.fst_t_next[0] ));
 sg13g2_or2_1 \u_neuron.u_fst/_074_  (.X(\u_neuron.u_fst/_032_ ),
    .B(net435),
    .A(\u_neuron.fst_t[1] ));
 sg13g2_a221oi_1 \u_neuron.u_fst/_075_  (.B2(\u_neuron.u_fst/_024_ ),
    .C1(\u_neuron.u_fst/_010_ ),
    .B1(\u_neuron.u_fst/_032_ ),
    .A1(\u_neuron.u_fst/_023_ ),
    .Y(\u_neuron.u_fst/_033_ ),
    .A2(\u_neuron.u_fst/_026_ ));
 sg13g2_a221oi_1 \u_neuron.u_fst/_076_  (.B2(\u_neuron.u_fst/_020_ ),
    .C1(\u_neuron.arm_event ),
    .B1(\u_neuron.u_fst/_033_ ),
    .A1(\u_neuron.u_fst/_011_ ),
    .Y(\u_neuron.fst_t_next[1] ),
    .A2(\u_neuron.u_fst/_029_ ));
 sg13g2_nand2_1 \u_neuron.u_fst/_077_  (.Y(\u_neuron.u_fst/_034_ ),
    .A(\u_neuron.u_fst/_013_ ),
    .B(\u_neuron.u_fst/_024_ ));
 sg13g2_a221oi_1 \u_neuron.u_fst/_078_  (.B2(\u_neuron.u_fst/_025_ ),
    .C1(\u_neuron.u_fst/_010_ ),
    .B1(\u_neuron.u_fst/_034_ ),
    .A1(\u_neuron.u_fst/_023_ ),
    .Y(\u_neuron.u_fst/_035_ ),
    .A2(\u_neuron.u_fst/_026_ ));
 sg13g2_a221oi_1 \u_neuron.u_fst/_079_  (.B2(\u_neuron.u_fst/_020_ ),
    .C1(\u_neuron.arm_event ),
    .B1(\u_neuron.u_fst/_035_ ),
    .A1(\u_neuron.u_fst/_013_ ),
    .Y(\u_neuron.fst_t_next[2] ),
    .A2(\u_neuron.u_fst/_029_ ));
 sg13g2_nor3_1 \u_neuron.u_fst/_080_  (.A(\u_neuron.u_fst/_023_ ),
    .B(\u_neuron.u_fst/_027_ ),
    .C(\u_neuron.u_fst/_029_ ),
    .Y(\u_neuron.u_fst/_036_ ));
 sg13g2_or2_1 \u_neuron.u_fst/_081_  (.X(\u_neuron.u_fst/_037_ ),
    .B(\u_neuron.u_fst/_029_ ),
    .A(\u_neuron.u_fst/_025_ ));
 sg13g2_a221oi_1 \u_neuron.u_fst/_082_  (.B2(\u_neuron.u_fst/_012_ ),
    .C1(\u_neuron.arm_event ),
    .B1(\u_neuron.u_fst/_037_ ),
    .A1(\u_neuron.u_fst/_026_ ),
    .Y(\u_neuron.fst_t_next[3] ),
    .A2(\u_neuron.u_fst/_030_ ));
 sg13g2_o21ai_1 \u_neuron.u_fst/_083_  (.B1(\u_neuron.u_fst/_016_ ),
    .Y(\u_neuron.u_fst/_038_ ),
    .A1(net159),
    .A2(\u_neuron.u_fst/_036_ ));
 sg13g2_a21oi_1 \u_neuron.u_fst/_084_  (.A1(net159),
    .A2(\u_neuron.u_fst/_036_ ),
    .Y(\u_neuron.fst_t_next[4] ),
    .B1(\u_neuron.u_fst/_038_ ));
 sg13g2_a21oi_1 \u_neuron.u_fst/_085_  (.A1(\u_neuron.fst_t[4] ),
    .A2(\u_neuron.u_fst/_036_ ),
    .Y(\u_neuron.u_fst/_039_ ),
    .B1(net116));
 sg13g2_nor4_1 \u_neuron.u_fst/_086_  (.A(\u_neuron.u_fst/_022_ ),
    .B(\u_neuron.u_fst/_023_ ),
    .C(\u_neuron.u_fst/_027_ ),
    .D(\u_neuron.u_fst/_029_ ),
    .Y(\u_neuron.u_fst/_040_ ));
 sg13g2_nor3_1 \u_neuron.u_fst/_087_  (.A(\u_neuron.arm_event ),
    .B(\u_neuron.u_fst/_039_ ),
    .C(\u_neuron.u_fst/_040_ ),
    .Y(\u_neuron.fst_t_next[5] ));
 sg13g2_nor4_1 \u_neuron.u_fst/_088_  (.A(\u_neuron.u_fst/_014_ ),
    .B(\u_neuron.u_fst/_022_ ),
    .C(\u_neuron.u_fst/_027_ ),
    .D(\u_neuron.u_fst/_029_ ),
    .Y(\u_neuron.u_fst/_041_ ));
 sg13g2_o21ai_1 \u_neuron.u_fst/_089_  (.B1(\u_neuron.u_fst/_016_ ),
    .Y(\u_neuron.u_fst/_042_ ),
    .A1(net136),
    .A2(\u_neuron.u_fst/_040_ ));
 sg13g2_a21oi_1 \u_neuron.u_fst/_090_  (.A1(\u_neuron.u_fst/_015_ ),
    .A2(\u_neuron.u_fst/_041_ ),
    .Y(\u_neuron.fst_t_next[6] ),
    .B1(\u_neuron.u_fst/_042_ ));
 sg13g2_nor2_1 \u_neuron.u_fst/_091_  (.A(net133),
    .B(\u_neuron.u_fst/_041_ ),
    .Y(\u_neuron.u_fst/_043_ ));
 sg13g2_nor2_1 \u_neuron.u_fst/_092_  (.A(\u_neuron.arm_event ),
    .B(\u_neuron.u_fst/_043_ ),
    .Y(\u_neuron.fst_t_next[7] ));
 sg13g2_nor2_1 \u_neuron.u_fst/_093_  (.A(net435),
    .B(net323),
    .Y(\u_neuron.u_fst/_044_ ));
 sg13g2_a21oi_1 \u_neuron.u_fst/_094_  (.A1(\u_neuron.u_fst/_017_ ),
    .A2(net323),
    .Y(\u_neuron.fst_last_t_next[0] ),
    .B1(\u_neuron.u_fst/_044_ ));
 sg13g2_nand2_1 \u_neuron.u_fst/_095_  (.Y(\u_neuron.u_fst/_045_ ),
    .A(net109),
    .B(net323));
 sg13g2_o21ai_1 \u_neuron.u_fst/_096_  (.B1(\u_neuron.u_fst/_045_ ),
    .Y(\u_neuron.fst_last_t_next[1] ),
    .A1(\u_neuron.u_fst/_011_ ),
    .A2(net323));
 sg13g2_nand2_1 \u_neuron.u_fst/_097_  (.Y(\u_neuron.u_fst/_046_ ),
    .A(net104),
    .B(net323));
 sg13g2_o21ai_1 \u_neuron.u_fst/_098_  (.B1(\u_neuron.u_fst/_046_ ),
    .Y(\u_neuron.fst_last_t_next[2] ),
    .A1(\u_neuron.u_fst/_013_ ),
    .A2(net323));
 sg13g2_nand2_1 \u_neuron.u_fst/_099_  (.Y(\u_neuron.u_fst/_047_ ),
    .A(net88),
    .B(net322));
 sg13g2_o21ai_1 \u_neuron.u_fst/_100_  (.B1(\u_neuron.u_fst/_047_ ),
    .Y(\u_neuron.fst_last_t_next[3] ),
    .A1(\u_neuron.u_fst/_012_ ),
    .A2(net322));
 sg13g2_mux2_1 \u_neuron.u_fst/_101_  (.A0(\u_neuron.fst_t[4] ),
    .A1(net62),
    .S(net322),
    .X(\u_neuron.fst_last_t_next[4] ));
 sg13g2_mux2_1 \u_neuron.u_fst/_102_  (.A0(\u_neuron.fst_t[5] ),
    .A1(net66),
    .S(net322),
    .X(\u_neuron.fst_last_t_next[5] ));
 sg13g2_nand2_1 \u_neuron.u_fst/_103_  (.Y(\u_neuron.u_fst/_000_ ),
    .A(net73),
    .B(net322));
 sg13g2_o21ai_1 \u_neuron.u_fst/_104_  (.B1(\u_neuron.u_fst/_000_ ),
    .Y(\u_neuron.fst_last_t_next[6] ),
    .A1(\u_neuron.u_fst/_014_ ),
    .A2(net322));
 sg13g2_nand2_1 \u_neuron.u_fst/_105_  (.Y(\u_neuron.u_fst/_001_ ),
    .A(net81),
    .B(net322));
 sg13g2_o21ai_1 \u_neuron.u_fst/_106_  (.B1(\u_neuron.u_fst/_001_ ),
    .Y(\u_neuron.fst_last_t_next[7] ),
    .A1(\u_neuron.u_fst/_015_ ),
    .A2(net322));
 sg13g2_a221oi_1 \u_neuron.u_fst/_107_  (.B2(net435),
    .C1(\u_neuron.fst_post_spike ),
    .B1(\u_neuron.u_fst/_028_ ),
    .A1(\u_neuron.u_fst/_010_ ),
    .Y(\u_neuron.u_fst/_002_ ),
    .A2(\u_neuron.u_fst/_017_ ));
 sg13g2_a21o_1 \u_neuron.u_fst/_108_  (.A2(\u_neuron.fst_post_spike ),
    .A1(net435),
    .B1(\u_neuron.u_fst/_002_ ),
    .X(\u_neuron.fst_emit_data[0] ));
 sg13g2_nand2_1 \u_neuron.u_fst/_109_  (.Y(\u_neuron.u_fst/_003_ ),
    .A(\u_neuron.fst_t[1] ),
    .B(\u_neuron.fst_post_spike ));
 sg13g2_o21ai_1 \u_neuron.u_fst/_110_  (.B1(\u_neuron.fst_emit_data[6] ),
    .Y(\u_neuron.u_fst/_004_ ),
    .A1(\u_neuron.fst_armed ),
    .A2(\u_neuron.fst_last_t[1] ));
 sg13g2_o21ai_1 \u_neuron.u_fst/_111_  (.B1(\u_neuron.u_fst/_003_ ),
    .Y(\u_neuron.fst_emit_data[1] ),
    .A1(\u_neuron.u_fst/_033_ ),
    .A2(\u_neuron.u_fst/_004_ ));
 sg13g2_o21ai_1 \u_neuron.u_fst/_112_  (.B1(\u_neuron.fst_emit_data[6] ),
    .Y(\u_neuron.u_fst/_005_ ),
    .A1(\u_neuron.fst_armed ),
    .A2(\u_neuron.fst_last_t[2] ));
 sg13g2_nand2_1 \u_neuron.u_fst/_113_  (.Y(\u_neuron.u_fst/_006_ ),
    .A(\u_neuron.fst_t[2] ),
    .B(\u_neuron.fst_post_spike ));
 sg13g2_o21ai_1 \u_neuron.u_fst/_114_  (.B1(\u_neuron.u_fst/_006_ ),
    .Y(\u_neuron.fst_emit_data[2] ),
    .A1(\u_neuron.u_fst/_035_ ),
    .A2(\u_neuron.u_fst/_005_ ));
 sg13g2_a21oi_1 \u_neuron.u_fst/_115_  (.A1(\u_neuron.u_fst/_012_ ),
    .A2(\u_neuron.u_fst/_025_ ),
    .Y(\u_neuron.u_fst/_007_ ),
    .B1(\u_neuron.u_fst/_010_ ));
 sg13g2_o21ai_1 \u_neuron.u_fst/_116_  (.B1(\u_neuron.u_fst/_007_ ),
    .Y(\u_neuron.u_fst/_008_ ),
    .A1(\u_neuron.u_fst/_023_ ),
    .A2(\u_neuron.u_fst/_027_ ));
 sg13g2_a21oi_1 \u_neuron.u_fst/_117_  (.A1(\u_neuron.u_fst/_010_ ),
    .A2(\u_neuron.fst_last_t[3] ),
    .Y(\u_neuron.u_fst/_009_ ),
    .B1(\u_neuron.fst_post_spike ));
 sg13g2_a22oi_1 \u_neuron.u_fst/_118_  (.Y(\u_neuron.fst_emit_data[3] ),
    .B1(\u_neuron.u_fst/_008_ ),
    .B2(\u_neuron.u_fst/_009_ ),
    .A2(\u_neuron.fst_post_spike ),
    .A1(\u_neuron.u_fst/_012_ ));
 sg13g2_o21ai_1 \u_neuron.u_fst/_119_  (.B1(\u_neuron.u_fst/_016_ ),
    .Y(\u_neuron.fst_armed_next ),
    .A1(\u_neuron.u_fst/_010_ ),
    .A2(\u_neuron.u_fst/_018_ ));
 sg13g2_tiehi \u_neuron.u_mode_sel/_09__41  (.L_HI(net41));
 sg13g2_tielo \u_neuron.u_mode_sel/_00__33  (.L_LO(net33));
 sg13g2_tielo \u_neuron.u_mode_sel/_07__34  (.L_LO(net34));
 sg13g2_buf_1 \u_neuron.u_fst/_123_  (.A(\u_neuron.fst_emit_data[6] ),
    .X(\u_neuron.fst_emit_data[4] ));
 sg13g2_inv_1 \u_neuron.u_learning/_151_  (.Y(\u_neuron.u_learning/_118_ ),
    .A(\u_neuron.soft_reset_fire ));
 sg13g2_inv_1 \u_neuron.u_learning/_152_  (.Y(\u_neuron.u_learning/_119_ ),
    .A(net235));
 sg13g2_inv_1 \u_neuron.u_learning/_153_  (.Y(\u_neuron.u_learning/_120_ ),
    .A(net421));
 sg13g2_inv_1 \u_neuron.u_learning/_154_  (.Y(\u_neuron.u_learning/_121_ ),
    .A(\u_neuron.pre_trace[1] ));
 sg13g2_inv_1 \u_neuron.u_learning/_155_  (.Y(\u_neuron.u_learning/_122_ ),
    .A(net427));
 sg13g2_inv_1 \u_neuron.u_learning/_156_  (.Y(\u_neuron.u_learning/_123_ ),
    .A(\u_neuron.pre_trace[2] ));
 sg13g2_inv_1 \u_neuron.u_learning/_157_  (.Y(\u_neuron.u_learning/_124_ ),
    .A(\u_neuron.pre_trace[3] ));
 sg13g2_inv_1 \u_neuron.u_learning/_158_  (.Y(\u_neuron.u_learning/_125_ ),
    .A(net424));
 sg13g2_inv_1 \u_neuron.u_learning/_159_  (.Y(\u_neuron.u_learning/_126_ ),
    .A(\u_neuron.pre_trace[6] ));
 sg13g2_inv_1 \u_neuron.u_learning/_160_  (.Y(\u_neuron.u_learning/_127_ ),
    .A(\u_neuron.pre_trace[7] ));
 sg13g2_inv_1 \u_neuron.u_learning/_161_  (.Y(\u_neuron.u_learning/_128_ ),
    .A(\u_neuron.pre_trace[9] ));
 sg13g2_inv_1 \u_neuron.u_learning/_162_  (.Y(\u_neuron.u_learning/_129_ ),
    .A(\u_neuron.pre_trace[10] ));
 sg13g2_inv_1 \u_neuron.u_learning/_163_  (.Y(\u_neuron.u_learning/_130_ ),
    .A(\u_neuron.pre_trace[11] ));
 sg13g2_inv_1 \u_neuron.u_learning/_164_  (.Y(\u_neuron.u_learning/_131_ ),
    .A(\u_neuron.pre_trace[13] ));
 sg13g2_inv_1 \u_neuron.u_learning/_165_  (.Y(\u_neuron.u_learning/_132_ ),
    .A(\u_neuron.pre_trace[14] ));
 sg13g2_inv_1 \u_neuron.u_learning/_166_  (.Y(\u_neuron.u_learning/_133_ ),
    .A(net212));
 sg13g2_inv_2 \u_neuron.u_learning/_167_  (.Y(\u_neuron.u_learning/_134_ ),
    .A(net388));
 sg13g2_nor2b_2 \u_neuron.u_learning/_168_  (.A(net424),
    .B_N(net427),
    .Y(\u_neuron.u_learning/_135_ ));
 sg13g2_nand2b_1 \u_neuron.u_learning/_169_  (.Y(\u_neuron.u_learning/_136_ ),
    .B(\u_neuron.u_learning/_135_ ),
    .A_N(\u_neuron.pre_trace[5] ));
 sg13g2_nor3_1 \u_neuron.u_learning/_170_  (.A(net427),
    .B(net424),
    .C(\u_neuron.pre_trace[4] ),
    .Y(\u_neuron.u_learning/_137_ ));
 sg13g2_and2_1 \u_neuron.u_learning/_171_  (.A(net427),
    .B(net424),
    .X(\u_neuron.u_learning/_138_ ));
 sg13g2_nor2b_2 \u_neuron.u_learning/_172_  (.A(net428),
    .B_N(net424),
    .Y(\u_neuron.u_learning/_139_ ));
 sg13g2_a221oi_1 \u_neuron.u_learning/_173_  (.B2(\u_neuron.u_learning/_126_ ),
    .C1(\u_neuron.u_learning/_137_ ),
    .B1(\u_neuron.u_learning/_139_ ),
    .A1(\u_neuron.u_learning/_127_ ),
    .Y(\u_neuron.u_learning/_140_ ),
    .A2(\u_neuron.u_learning/_138_ ));
 sg13g2_nand3_1 \u_neuron.u_learning/_174_  (.B(\u_neuron.u_learning/_136_ ),
    .C(\u_neuron.u_learning/_140_ ),
    .A(net421),
    .Y(\u_neuron.u_learning/_141_ ));
 sg13g2_nor3_1 \u_neuron.u_learning/_175_  (.A(\u_neuron.pre_trace[0] ),
    .B(net428),
    .C(net425),
    .Y(\u_neuron.u_learning/_142_ ));
 sg13g2_a21oi_1 \u_neuron.u_learning/_176_  (.A1(\u_neuron.u_learning/_124_ ),
    .A2(\u_neuron.u_learning/_138_ ),
    .Y(\u_neuron.u_learning/_143_ ),
    .B1(net422));
 sg13g2_a221oi_1 \u_neuron.u_learning/_177_  (.B2(\u_neuron.u_learning/_123_ ),
    .C1(\u_neuron.u_learning/_142_ ),
    .B1(\u_neuron.u_learning/_139_ ),
    .A1(\u_neuron.u_learning/_121_ ),
    .Y(\u_neuron.u_learning/_144_ ),
    .A2(\u_neuron.u_learning/_135_ ));
 sg13g2_a21oi_1 \u_neuron.u_learning/_178_  (.A1(\u_neuron.u_learning/_143_ ),
    .A2(\u_neuron.u_learning/_144_ ),
    .Y(\u_neuron.u_learning/_145_ ),
    .B1(net419));
 sg13g2_a21oi_1 \u_neuron.u_learning/_179_  (.A1(\u_neuron.u_learning/_130_ ),
    .A2(\u_neuron.u_learning/_138_ ),
    .Y(\u_neuron.u_learning/_146_ ),
    .B1(net422));
 sg13g2_nor3_1 \u_neuron.u_learning/_180_  (.A(net428),
    .B(net425),
    .C(\u_neuron.pre_trace[8] ),
    .Y(\u_neuron.u_learning/_147_ ));
 sg13g2_a221oi_1 \u_neuron.u_learning/_181_  (.B2(\u_neuron.u_learning/_129_ ),
    .C1(\u_neuron.u_learning/_147_ ),
    .B1(\u_neuron.u_learning/_139_ ),
    .A1(\u_neuron.u_learning/_128_ ),
    .Y(\u_neuron.u_learning/_148_ ),
    .A2(\u_neuron.u_learning/_135_ ));
 sg13g2_a21oi_1 \u_neuron.u_learning/_182_  (.A1(\u_neuron.u_learning/_132_ ),
    .A2(\u_neuron.u_learning/_139_ ),
    .Y(\u_neuron.u_learning/_149_ ),
    .B1(\u_neuron.u_learning/_120_ ));
 sg13g2_nor3_1 \u_neuron.u_learning/_183_  (.A(net427),
    .B(net424),
    .C(\u_neuron.pre_trace[12] ),
    .Y(\u_neuron.u_learning/_150_ ));
 sg13g2_a221oi_1 \u_neuron.u_learning/_184_  (.B2(\u_neuron.u_learning/_133_ ),
    .C1(\u_neuron.u_learning/_150_ ),
    .B1(\u_neuron.u_learning/_138_ ),
    .A1(\u_neuron.u_learning/_131_ ),
    .Y(\u_neuron.u_learning/_022_ ),
    .A2(\u_neuron.u_learning/_135_ ));
 sg13g2_a22oi_1 \u_neuron.u_learning/_185_  (.Y(\u_neuron.u_learning/_023_ ),
    .B1(\u_neuron.u_learning/_149_ ),
    .B2(\u_neuron.u_learning/_022_ ),
    .A2(\u_neuron.u_learning/_148_ ),
    .A1(\u_neuron.u_learning/_146_ ));
 sg13g2_nand2_1 \u_neuron.u_learning/_186_  (.Y(\u_neuron.u_learning/_024_ ),
    .A(net356),
    .B(\u_neuron.learn_pending ));
 sg13g2_a221oi_1 \u_neuron.u_learning/_187_  (.B2(net419),
    .C1(\u_neuron.u_learning/_024_ ),
    .B1(\u_neuron.u_learning/_023_ ),
    .A1(\u_neuron.u_learning/_141_ ),
    .Y(\u_neuron.ltp_we ),
    .A2(\u_neuron.u_learning/_145_ ));
 sg13g2_nor2b_1 \u_neuron.u_learning/_188_  (.A(net384),
    .B_N(\u_neuron.is_prog_addr ),
    .Y(\u_neuron.u_learning/_025_ ));
 sg13g2_and4_1 \u_neuron.u_learning/_189_  (.A(net356),
    .B(\u_neuron.learn_en ),
    .C(\u_neuron.post_trace ),
    .D(net366),
    .X(\u_neuron.ltd_we ));
 sg13g2_nand2b_2 \u_neuron.u_learning/_190_  (.Y(\u_neuron.ltp_wdata[0] ),
    .B(\u_neuron.w_ptr_curr[0] ),
    .A_N(\u_neuron.w_ptr_curr[1] ));
 sg13g2_or2_1 \u_neuron.u_learning/_191_  (.X(\u_neuron.ltp_wdata[1] ),
    .B(\u_neuron.w_ptr_curr[0] ),
    .A(\u_neuron.w_ptr_curr[1] ));
 sg13g2_nor2b_2 \u_neuron.u_learning/_192_  (.A(\u_neuron.w_addr_curr[0] ),
    .B_N(\u_neuron.w_addr_curr[1] ),
    .Y(\u_neuron.ltd_wdata[0] ));
 sg13g2_and2_1 \u_neuron.u_learning/_193_  (.A(\u_neuron.w_addr_curr[1] ),
    .B(\u_neuron.w_addr_curr[0] ),
    .X(\u_neuron.ltd_wdata[1] ));
 sg13g2_nor3_2 \u_neuron.u_learning/_194_  (.A(net421),
    .B(net427),
    .C(net424),
    .Y(\u_neuron.u_learning/_026_ ));
 sg13g2_and2_1 \u_neuron.u_learning/_195_  (.A(net465),
    .B(net356),
    .X(\u_neuron.u_learning/_027_ ));
 sg13g2_nand2_1 \u_neuron.u_learning/_196_  (.Y(\u_neuron.u_learning/_028_ ),
    .A(net465),
    .B(net356));
 sg13g2_and3_2 \u_neuron.u_learning/_197_  (.X(\u_neuron.u_learning/_029_ ),
    .A(net465),
    .B(net356),
    .C(net200));
 sg13g2_nand2_1 \u_neuron.u_learning/_198_  (.Y(\u_neuron.u_learning/_030_ ),
    .A(net200),
    .B(net330));
 sg13g2_xnor2_1 \u_neuron.u_learning/_199_  (.Y(\u_neuron.u_learning/_031_ ),
    .A(net419),
    .B(\u_neuron.u_learning/_026_ ));
 sg13g2_xor2_1 \u_neuron.u_learning/_200_  (.B(\u_neuron.u_learning/_026_ ),
    .A(net419),
    .X(\u_neuron.u_learning/_032_ ));
 sg13g2_nand3b_1 \u_neuron.u_learning/_201_  (.B(\u_neuron.u_learning/_026_ ),
    .C(\u_neuron.u_learning/_029_ ),
    .Y(\u_neuron.u_learning/_033_ ),
    .A_N(net419));
 sg13g2_nand3_1 \u_neuron.u_learning/_202_  (.B(net85),
    .C(\u_neuron.u_learning/_033_ ),
    .A(net362),
    .Y(\u_neuron.u_learning/_034_ ));
 sg13g2_nor3_2 \u_neuron.u_learning/_203_  (.A(net388),
    .B(net393),
    .C(net399),
    .Y(\u_neuron.u_learning/_035_ ));
 sg13g2_nor2_1 \u_neuron.u_learning/_204_  (.A(\u_neuron.soft_reset_fire ),
    .B(\u_neuron.u_learning/_028_ ),
    .Y(\u_neuron.u_learning/_036_ ));
 sg13g2_nand3b_1 \u_neuron.u_learning/_205_  (.B(net356),
    .C(net465),
    .Y(\u_neuron.u_learning/_037_ ),
    .A_N(\u_neuron.soft_reset_fire ));
 sg13g2_nand3b_1 \u_neuron.u_learning/_206_  (.B(net366),
    .C(\u_neuron.u_learning/_035_ ),
    .Y(\u_neuron.u_learning/_038_ ),
    .A_N(net386));
 sg13g2_o21ai_1 \u_neuron.u_learning/_207_  (.B1(net86),
    .Y(\u_neuron.u_learning/_000_ ),
    .A1(\u_neuron.u_learning/_037_ ),
    .A2(\u_neuron.u_learning/_038_ ));
 sg13g2_xnor2_1 \u_neuron.u_learning/_208_  (.Y(\u_neuron.u_learning/_039_ ),
    .A(net386),
    .B(\u_neuron.u_learning/_035_ ));
 sg13g2_xor2_1 \u_neuron.u_learning/_209_  (.B(\u_neuron.u_learning/_035_ ),
    .A(net386),
    .X(\u_neuron.u_learning/_040_ ));
 sg13g2_nand2b_1 \u_neuron.u_learning/_210_  (.Y(\u_neuron.u_learning/_041_ ),
    .B(net399),
    .A_N(net393));
 sg13g2_nor3_1 \u_neuron.u_learning/_211_  (.A(net388),
    .B(\u_neuron.u_learning/_037_ ),
    .C(\u_neuron.u_learning/_041_ ),
    .Y(\u_neuron.u_learning/_042_ ));
 sg13g2_nand3_1 \u_neuron.u_learning/_212_  (.B(\u_neuron.u_learning/_039_ ),
    .C(\u_neuron.u_learning/_042_ ),
    .A(net364),
    .Y(\u_neuron.u_learning/_043_ ));
 sg13g2_nand3_1 \u_neuron.u_learning/_213_  (.B(\u_neuron.u_learning/_135_ ),
    .C(net330),
    .A(\u_neuron.u_learning/_120_ ),
    .Y(\u_neuron.u_learning/_044_ ));
 sg13g2_nor3_1 \u_neuron.u_learning/_214_  (.A(net381),
    .B(\u_neuron.u_learning/_032_ ),
    .C(\u_neuron.u_learning/_044_ ),
    .Y(\u_neuron.u_learning/_045_ ));
 sg13g2_nand2_1 \u_neuron.u_learning/_215_  (.Y(\u_neuron.u_learning/_046_ ),
    .A(net362),
    .B(net91));
 sg13g2_o21ai_1 \u_neuron.u_learning/_216_  (.B1(\u_neuron.u_learning/_043_ ),
    .Y(\u_neuron.u_learning/_001_ ),
    .A1(\u_neuron.u_learning/_045_ ),
    .A2(\u_neuron.u_learning/_046_ ));
 sg13g2_nand2b_1 \u_neuron.u_learning/_217_  (.Y(\u_neuron.u_learning/_047_ ),
    .B(net393),
    .A_N(net399));
 sg13g2_nor3_1 \u_neuron.u_learning/_218_  (.A(net388),
    .B(\u_neuron.u_learning/_037_ ),
    .C(\u_neuron.u_learning/_047_ ),
    .Y(\u_neuron.u_learning/_048_ ));
 sg13g2_nand3_1 \u_neuron.u_learning/_219_  (.B(\u_neuron.u_learning/_039_ ),
    .C(\u_neuron.u_learning/_048_ ),
    .A(net364),
    .Y(\u_neuron.u_learning/_049_ ));
 sg13g2_nand3_1 \u_neuron.u_learning/_220_  (.B(\u_neuron.u_learning/_139_ ),
    .C(net330),
    .A(\u_neuron.u_learning/_120_ ),
    .Y(\u_neuron.u_learning/_050_ ));
 sg13g2_nor3_1 \u_neuron.u_learning/_221_  (.A(net381),
    .B(\u_neuron.u_learning/_032_ ),
    .C(\u_neuron.u_learning/_050_ ),
    .Y(\u_neuron.u_learning/_051_ ));
 sg13g2_nand2_1 \u_neuron.u_learning/_222_  (.Y(\u_neuron.u_learning/_052_ ),
    .A(net361),
    .B(net90));
 sg13g2_o21ai_1 \u_neuron.u_learning/_223_  (.B1(\u_neuron.u_learning/_049_ ),
    .Y(\u_neuron.u_learning/_002_ ),
    .A1(\u_neuron.u_learning/_051_ ),
    .A2(\u_neuron.u_learning/_052_ ));
 sg13g2_nand2_1 \u_neuron.u_learning/_224_  (.Y(\u_neuron.u_learning/_053_ ),
    .A(net393),
    .B(net399));
 sg13g2_nor3_1 \u_neuron.u_learning/_225_  (.A(net388),
    .B(\u_neuron.u_learning/_037_ ),
    .C(\u_neuron.u_learning/_053_ ),
    .Y(\u_neuron.u_learning/_054_ ));
 sg13g2_nand3_1 \u_neuron.u_learning/_226_  (.B(\u_neuron.u_learning/_039_ ),
    .C(\u_neuron.u_learning/_054_ ),
    .A(net364),
    .Y(\u_neuron.u_learning/_055_ ));
 sg13g2_nand3_1 \u_neuron.u_learning/_227_  (.B(\u_neuron.u_learning/_138_ ),
    .C(net330),
    .A(\u_neuron.u_learning/_120_ ),
    .Y(\u_neuron.u_learning/_056_ ));
 sg13g2_nor3_1 \u_neuron.u_learning/_228_  (.A(net381),
    .B(\u_neuron.u_learning/_032_ ),
    .C(\u_neuron.u_learning/_056_ ),
    .Y(\u_neuron.u_learning/_057_ ));
 sg13g2_nand2_1 \u_neuron.u_learning/_229_  (.Y(\u_neuron.u_learning/_058_ ),
    .A(net361),
    .B(net94));
 sg13g2_o21ai_1 \u_neuron.u_learning/_230_  (.B1(\u_neuron.u_learning/_055_ ),
    .Y(\u_neuron.u_learning/_003_ ),
    .A1(\u_neuron.u_learning/_057_ ),
    .A2(\u_neuron.u_learning/_058_ ));
 sg13g2_nor4_1 \u_neuron.u_learning/_231_  (.A(\u_neuron.u_learning/_134_ ),
    .B(net393),
    .C(net399),
    .D(\u_neuron.u_learning/_037_ ),
    .Y(\u_neuron.u_learning/_059_ ));
 sg13g2_nand3_1 \u_neuron.u_learning/_232_  (.B(\u_neuron.u_learning/_039_ ),
    .C(\u_neuron.u_learning/_059_ ),
    .A(net364),
    .Y(\u_neuron.u_learning/_060_ ));
 sg13g2_nand4_1 \u_neuron.u_learning/_233_  (.B(\u_neuron.u_learning/_122_ ),
    .C(\u_neuron.u_learning/_125_ ),
    .A(net421),
    .Y(\u_neuron.u_learning/_061_ ),
    .D(net330));
 sg13g2_nor3_1 \u_neuron.u_learning/_234_  (.A(net380),
    .B(\u_neuron.u_learning/_032_ ),
    .C(\u_neuron.u_learning/_061_ ),
    .Y(\u_neuron.u_learning/_062_ ));
 sg13g2_nand2_1 \u_neuron.u_learning/_235_  (.Y(\u_neuron.u_learning/_063_ ),
    .A(net363),
    .B(net101));
 sg13g2_o21ai_1 \u_neuron.u_learning/_236_  (.B1(\u_neuron.u_learning/_060_ ),
    .Y(\u_neuron.u_learning/_004_ ),
    .A1(\u_neuron.u_learning/_062_ ),
    .A2(\u_neuron.u_learning/_063_ ));
 sg13g2_nor3_1 \u_neuron.u_learning/_237_  (.A(\u_neuron.u_learning/_134_ ),
    .B(\u_neuron.u_learning/_037_ ),
    .C(\u_neuron.u_learning/_041_ ),
    .Y(\u_neuron.u_learning/_064_ ));
 sg13g2_nand3_1 \u_neuron.u_learning/_238_  (.B(\u_neuron.u_learning/_039_ ),
    .C(\u_neuron.u_learning/_064_ ),
    .A(net364),
    .Y(\u_neuron.u_learning/_065_ ));
 sg13g2_nand3_1 \u_neuron.u_learning/_239_  (.B(\u_neuron.u_learning/_135_ ),
    .C(net330),
    .A(net421),
    .Y(\u_neuron.u_learning/_066_ ));
 sg13g2_nor3_1 \u_neuron.u_learning/_240_  (.A(net380),
    .B(\u_neuron.u_learning/_032_ ),
    .C(\u_neuron.u_learning/_066_ ),
    .Y(\u_neuron.u_learning/_067_ ));
 sg13g2_nand2_1 \u_neuron.u_learning/_241_  (.Y(\u_neuron.u_learning/_068_ ),
    .A(net361),
    .B(net106));
 sg13g2_o21ai_1 \u_neuron.u_learning/_242_  (.B1(\u_neuron.u_learning/_065_ ),
    .Y(\u_neuron.u_learning/_005_ ),
    .A1(\u_neuron.u_learning/_067_ ),
    .A2(\u_neuron.u_learning/_068_ ));
 sg13g2_nor3_1 \u_neuron.u_learning/_243_  (.A(\u_neuron.u_learning/_134_ ),
    .B(\u_neuron.u_learning/_037_ ),
    .C(\u_neuron.u_learning/_047_ ),
    .Y(\u_neuron.u_learning/_069_ ));
 sg13g2_nand3_1 \u_neuron.u_learning/_244_  (.B(\u_neuron.u_learning/_039_ ),
    .C(\u_neuron.u_learning/_069_ ),
    .A(net365),
    .Y(\u_neuron.u_learning/_070_ ));
 sg13g2_nand3_1 \u_neuron.u_learning/_245_  (.B(\u_neuron.u_learning/_139_ ),
    .C(\u_neuron.u_learning/_027_ ),
    .A(net422),
    .Y(\u_neuron.u_learning/_071_ ));
 sg13g2_nor3_1 \u_neuron.u_learning/_246_  (.A(net381),
    .B(\u_neuron.u_learning/_032_ ),
    .C(\u_neuron.u_learning/_071_ ),
    .Y(\u_neuron.u_learning/_072_ ));
 sg13g2_nand2_1 \u_neuron.u_learning/_247_  (.Y(\u_neuron.u_learning/_073_ ),
    .A(net361),
    .B(net102));
 sg13g2_o21ai_1 \u_neuron.u_learning/_248_  (.B1(\u_neuron.u_learning/_070_ ),
    .Y(\u_neuron.u_learning/_006_ ),
    .A1(\u_neuron.u_learning/_072_ ),
    .A2(\u_neuron.u_learning/_073_ ));
 sg13g2_nor3_1 \u_neuron.u_learning/_249_  (.A(\u_neuron.u_learning/_134_ ),
    .B(\u_neuron.u_learning/_037_ ),
    .C(\u_neuron.u_learning/_053_ ),
    .Y(\u_neuron.u_learning/_074_ ));
 sg13g2_nand4_1 \u_neuron.u_learning/_250_  (.B(net393),
    .C(net399),
    .A(net388),
    .Y(\u_neuron.u_learning/_075_ ),
    .D(\u_neuron.u_learning/_036_ ));
 sg13g2_nand3_1 \u_neuron.u_learning/_251_  (.B(\u_neuron.u_learning/_039_ ),
    .C(\u_neuron.u_learning/_074_ ),
    .A(net364),
    .Y(\u_neuron.u_learning/_076_ ));
 sg13g2_and3_1 \u_neuron.u_learning/_252_  (.X(\u_neuron.u_learning/_077_ ),
    .A(net421),
    .B(net427),
    .C(net424));
 sg13g2_and4_1 \u_neuron.u_learning/_253_  (.A(\u_neuron.learn_pending ),
    .B(net330),
    .C(\u_neuron.u_learning/_031_ ),
    .D(\u_neuron.u_learning/_077_ ),
    .X(\u_neuron.u_learning/_078_ ));
 sg13g2_nand2_1 \u_neuron.u_learning/_254_  (.Y(\u_neuron.u_learning/_079_ ),
    .A(net361),
    .B(net96));
 sg13g2_o21ai_1 \u_neuron.u_learning/_255_  (.B1(\u_neuron.u_learning/_076_ ),
    .Y(\u_neuron.u_learning/_007_ ),
    .A1(\u_neuron.u_learning/_078_ ),
    .A2(\u_neuron.u_learning/_079_ ));
 sg13g2_nand3_1 \u_neuron.u_learning/_256_  (.B(\u_neuron.u_learning/_026_ ),
    .C(\u_neuron.u_learning/_029_ ),
    .A(net419),
    .Y(\u_neuron.u_learning/_080_ ));
 sg13g2_nand3_1 \u_neuron.u_learning/_257_  (.B(net107),
    .C(\u_neuron.u_learning/_080_ ),
    .A(net362),
    .Y(\u_neuron.u_learning/_081_ ));
 sg13g2_nand4_1 \u_neuron.u_learning/_258_  (.B(net366),
    .C(\u_neuron.u_learning/_036_ ),
    .A(net386),
    .Y(\u_neuron.u_learning/_082_ ),
    .D(\u_neuron.u_learning/_039_ ));
 sg13g2_nand2_1 \u_neuron.u_learning/_259_  (.Y(\u_neuron.u_learning/_008_ ),
    .A(net108),
    .B(\u_neuron.u_learning/_082_ ));
 sg13g2_nand2_1 \u_neuron.u_learning/_260_  (.Y(\u_neuron.u_learning/_083_ ),
    .A(net366),
    .B(\u_neuron.u_learning/_040_ ));
 sg13g2_nand3_1 \u_neuron.u_learning/_261_  (.B(\u_neuron.u_learning/_040_ ),
    .C(\u_neuron.u_learning/_042_ ),
    .A(net365),
    .Y(\u_neuron.u_learning/_084_ ));
 sg13g2_nor3_1 \u_neuron.u_learning/_262_  (.A(net380),
    .B(\u_neuron.u_learning/_031_ ),
    .C(\u_neuron.u_learning/_044_ ),
    .Y(\u_neuron.u_learning/_085_ ));
 sg13g2_nand2_1 \u_neuron.u_learning/_263_  (.Y(\u_neuron.u_learning/_086_ ),
    .A(net361),
    .B(net92));
 sg13g2_o21ai_1 \u_neuron.u_learning/_264_  (.B1(\u_neuron.u_learning/_084_ ),
    .Y(\u_neuron.u_learning/_009_ ),
    .A1(\u_neuron.u_learning/_085_ ),
    .A2(\u_neuron.u_learning/_086_ ));
 sg13g2_nand3_1 \u_neuron.u_learning/_265_  (.B(\u_neuron.u_learning/_040_ ),
    .C(\u_neuron.u_learning/_048_ ),
    .A(net365),
    .Y(\u_neuron.u_learning/_087_ ));
 sg13g2_nor3_1 \u_neuron.u_learning/_266_  (.A(net380),
    .B(\u_neuron.u_learning/_031_ ),
    .C(\u_neuron.u_learning/_050_ ),
    .Y(\u_neuron.u_learning/_088_ ));
 sg13g2_nand2_1 \u_neuron.u_learning/_267_  (.Y(\u_neuron.u_learning/_089_ ),
    .A(net361),
    .B(net100));
 sg13g2_o21ai_1 \u_neuron.u_learning/_268_  (.B1(\u_neuron.u_learning/_087_ ),
    .Y(\u_neuron.u_learning/_010_ ),
    .A1(\u_neuron.u_learning/_088_ ),
    .A2(\u_neuron.u_learning/_089_ ));
 sg13g2_nand3_1 \u_neuron.u_learning/_269_  (.B(\u_neuron.u_learning/_040_ ),
    .C(\u_neuron.u_learning/_054_ ),
    .A(net365),
    .Y(\u_neuron.u_learning/_090_ ));
 sg13g2_nor3_1 \u_neuron.u_learning/_270_  (.A(net380),
    .B(\u_neuron.u_learning/_031_ ),
    .C(\u_neuron.u_learning/_056_ ),
    .Y(\u_neuron.u_learning/_091_ ));
 sg13g2_nand2_1 \u_neuron.u_learning/_271_  (.Y(\u_neuron.u_learning/_092_ ),
    .A(net361),
    .B(net122));
 sg13g2_o21ai_1 \u_neuron.u_learning/_272_  (.B1(\u_neuron.u_learning/_090_ ),
    .Y(\u_neuron.u_learning/_011_ ),
    .A1(\u_neuron.u_learning/_091_ ),
    .A2(\u_neuron.u_learning/_092_ ));
 sg13g2_nand3_1 \u_neuron.u_learning/_273_  (.B(\u_neuron.u_learning/_040_ ),
    .C(\u_neuron.u_learning/_059_ ),
    .A(net364),
    .Y(\u_neuron.u_learning/_093_ ));
 sg13g2_nor3_1 \u_neuron.u_learning/_274_  (.A(net380),
    .B(\u_neuron.u_learning/_031_ ),
    .C(\u_neuron.u_learning/_061_ ),
    .Y(\u_neuron.u_learning/_094_ ));
 sg13g2_nand2_1 \u_neuron.u_learning/_275_  (.Y(\u_neuron.u_learning/_095_ ),
    .A(net363),
    .B(net93));
 sg13g2_o21ai_1 \u_neuron.u_learning/_276_  (.B1(\u_neuron.u_learning/_093_ ),
    .Y(\u_neuron.u_learning/_012_ ),
    .A1(\u_neuron.u_learning/_094_ ),
    .A2(\u_neuron.u_learning/_095_ ));
 sg13g2_nand3_1 \u_neuron.u_learning/_277_  (.B(\u_neuron.u_learning/_040_ ),
    .C(\u_neuron.u_learning/_064_ ),
    .A(net364),
    .Y(\u_neuron.u_learning/_096_ ));
 sg13g2_nor3_1 \u_neuron.u_learning/_278_  (.A(net380),
    .B(\u_neuron.u_learning/_031_ ),
    .C(\u_neuron.u_learning/_066_ ),
    .Y(\u_neuron.u_learning/_097_ ));
 sg13g2_nand2_1 \u_neuron.u_learning/_279_  (.Y(\u_neuron.u_learning/_098_ ),
    .A(net363),
    .B(net95));
 sg13g2_o21ai_1 \u_neuron.u_learning/_280_  (.B1(\u_neuron.u_learning/_096_ ),
    .Y(\u_neuron.u_learning/_013_ ),
    .A1(\u_neuron.u_learning/_097_ ),
    .A2(\u_neuron.u_learning/_098_ ));
 sg13g2_nand3_1 \u_neuron.u_learning/_281_  (.B(\u_neuron.u_learning/_040_ ),
    .C(\u_neuron.u_learning/_069_ ),
    .A(net365),
    .Y(\u_neuron.u_learning/_099_ ));
 sg13g2_nor3_1 \u_neuron.u_learning/_282_  (.A(net380),
    .B(\u_neuron.u_learning/_031_ ),
    .C(\u_neuron.u_learning/_071_ ),
    .Y(\u_neuron.u_learning/_100_ ));
 sg13g2_nand2_1 \u_neuron.u_learning/_283_  (.Y(\u_neuron.u_learning/_101_ ),
    .A(net362),
    .B(net103));
 sg13g2_o21ai_1 \u_neuron.u_learning/_284_  (.B1(\u_neuron.u_learning/_099_ ),
    .Y(\u_neuron.u_learning/_014_ ),
    .A1(\u_neuron.u_learning/_100_ ),
    .A2(\u_neuron.u_learning/_101_ ));
 sg13g2_nand2_1 \u_neuron.u_learning/_285_  (.Y(\u_neuron.u_learning/_102_ ),
    .A(net419),
    .B(\u_neuron.u_learning/_077_ ));
 sg13g2_nor2_1 \u_neuron.u_learning/_286_  (.A(\u_neuron.u_learning/_030_ ),
    .B(\u_neuron.u_learning/_102_ ),
    .Y(\u_neuron.u_learning/_103_ ));
 sg13g2_nor2_1 \u_neuron.u_learning/_287_  (.A(\u_neuron.soft_reset_fire ),
    .B(\u_neuron.u_learning/_133_ ),
    .Y(\u_neuron.u_learning/_104_ ));
 sg13g2_o21ai_1 \u_neuron.u_learning/_288_  (.B1(\u_neuron.u_learning/_104_ ),
    .Y(\u_neuron.u_learning/_105_ ),
    .A1(\u_neuron.u_learning/_030_ ),
    .A2(\u_neuron.u_learning/_102_ ));
 sg13g2_o21ai_1 \u_neuron.u_learning/_289_  (.B1(net213),
    .Y(\u_neuron.u_learning/_015_ ),
    .A1(\u_neuron.u_learning/_075_ ),
    .A2(\u_neuron.u_learning/_083_ ));
 sg13g2_nand2_1 \u_neuron.u_learning/_290_  (.Y(\u_neuron.u_learning/_106_ ),
    .A(net363),
    .B(net206));
 sg13g2_a21oi_1 \u_neuron.u_learning/_291_  (.A1(net384),
    .A2(net330),
    .Y(\u_neuron.u_learning/_107_ ),
    .B1(\u_neuron.u_learning/_106_ ));
 sg13g2_a21o_1 \u_neuron.u_learning/_292_  (.A2(\u_neuron.u_learning/_036_ ),
    .A1(\u_neuron.mode_post_spike ),
    .B1(\u_neuron.u_learning/_107_ ),
    .X(\u_neuron.u_learning/_016_ ));
 sg13g2_nand4_1 \u_neuron.u_learning/_293_  (.B(net356),
    .C(\u_neuron.mode_learn_start ),
    .A(net465),
    .Y(\u_neuron.u_learning/_108_ ),
    .D(net209));
 sg13g2_o21ai_1 \u_neuron.u_learning/_294_  (.B1(net200),
    .Y(\u_neuron.u_learning/_109_ ),
    .A1(\u_neuron.u_learning/_028_ ),
    .A2(\u_neuron.u_learning/_102_ ));
 sg13g2_a21oi_1 \u_neuron.u_learning/_295_  (.A1(\u_neuron.u_learning/_108_ ),
    .A2(\u_neuron.u_learning/_109_ ),
    .Y(\u_neuron.u_learning/_017_ ),
    .B1(\u_neuron.soft_reset_fire ));
 sg13g2_nand2_1 \u_neuron.u_learning/_296_  (.Y(\u_neuron.u_learning/_110_ ),
    .A(net363),
    .B(\u_neuron.u_learning/_108_ ));
 sg13g2_a21oi_1 \u_neuron.u_learning/_297_  (.A1(\u_neuron.mode_learn_start ),
    .A2(net209),
    .Y(\u_neuron.u_learning/_111_ ),
    .B1(\u_neuron.soft_reset_fire ));
 sg13g2_a21o_1 \u_neuron.u_learning/_298_  (.A2(\u_neuron.u_learning/_029_ ),
    .A1(net427),
    .B1(\u_neuron.u_learning/_110_ ),
    .X(\u_neuron.u_learning/_112_ ));
 sg13g2_a21oi_1 \u_neuron.u_learning/_299_  (.A1(\u_neuron.u_learning/_122_ ),
    .A2(\u_neuron.u_learning/_030_ ),
    .Y(\u_neuron.u_learning/_018_ ),
    .B1(\u_neuron.u_learning/_112_ ));
 sg13g2_nand2_1 \u_neuron.u_learning/_300_  (.Y(\u_neuron.u_learning/_113_ ),
    .A(\u_neuron.u_learning/_029_ ),
    .B(\u_neuron.u_learning/_111_ ));
 sg13g2_nand3_1 \u_neuron.u_learning/_301_  (.B(\u_neuron.u_learning/_029_ ),
    .C(\u_neuron.u_learning/_111_ ),
    .A(\u_neuron.u_learning/_135_ ),
    .Y(\u_neuron.u_learning/_114_ ));
 sg13g2_o21ai_1 \u_neuron.u_learning/_302_  (.B1(\u_neuron.u_learning/_114_ ),
    .Y(\u_neuron.u_learning/_019_ ),
    .A1(\u_neuron.u_learning/_125_ ),
    .A2(\u_neuron.u_learning/_112_ ));
 sg13g2_nand4_1 \u_neuron.u_learning/_303_  (.B(net421),
    .C(\u_neuron.u_learning/_030_ ),
    .A(net363),
    .Y(\u_neuron.u_learning/_115_ ),
    .D(\u_neuron.u_learning/_108_ ));
 sg13g2_xnor2_1 \u_neuron.u_learning/_304_  (.Y(\u_neuron.u_learning/_116_ ),
    .A(net421),
    .B(\u_neuron.u_learning/_138_ ));
 sg13g2_o21ai_1 \u_neuron.u_learning/_305_  (.B1(\u_neuron.u_learning/_115_ ),
    .Y(\u_neuron.u_learning/_020_ ),
    .A1(\u_neuron.u_learning/_113_ ),
    .A2(\u_neuron.u_learning/_116_ ));
 sg13g2_a21oi_1 \u_neuron.u_learning/_306_  (.A1(\u_neuron.u_learning/_029_ ),
    .A2(\u_neuron.u_learning/_077_ ),
    .Y(\u_neuron.u_learning/_117_ ),
    .B1(net419));
 sg13g2_nor3_1 \u_neuron.u_learning/_307_  (.A(\u_neuron.u_learning/_103_ ),
    .B(\u_neuron.u_learning/_110_ ),
    .C(\u_neuron.u_learning/_117_ ),
    .Y(\u_neuron.u_learning/_021_ ));
 sg13g2_dfrbpq_1 \u_neuron.u_learning/_308_  (.RESET_B(net443),
    .D(\u_neuron.u_learning/_000_ ),
    .Q(\u_neuron.pre_trace[0] ),
    .CLK(clknet_5_9__leaf_clk));
 sg13g2_dfrbpq_1 \u_neuron.u_learning/_309_  (.RESET_B(net442),
    .D(\u_neuron.u_learning/_001_ ),
    .Q(\u_neuron.pre_trace[1] ),
    .CLK(clknet_5_11__leaf_clk));
 sg13g2_dfrbpq_1 \u_neuron.u_learning/_310_  (.RESET_B(net442),
    .D(\u_neuron.u_learning/_002_ ),
    .Q(\u_neuron.pre_trace[2] ),
    .CLK(clknet_5_10__leaf_clk));
 sg13g2_dfrbpq_1 \u_neuron.u_learning/_311_  (.RESET_B(net442),
    .D(\u_neuron.u_learning/_003_ ),
    .Q(\u_neuron.pre_trace[3] ),
    .CLK(clknet_5_10__leaf_clk));
 sg13g2_dfrbpq_1 \u_neuron.u_learning/_312_  (.RESET_B(net441),
    .D(\u_neuron.u_learning/_004_ ),
    .Q(\u_neuron.pre_trace[4] ),
    .CLK(clknet_5_8__leaf_clk));
 sg13g2_dfrbpq_1 \u_neuron.u_learning/_313_  (.RESET_B(net442),
    .D(\u_neuron.u_learning/_005_ ),
    .Q(\u_neuron.pre_trace[5] ),
    .CLK(clknet_5_10__leaf_clk));
 sg13g2_dfrbpq_1 \u_neuron.u_learning/_314_  (.RESET_B(net442),
    .D(\u_neuron.u_learning/_006_ ),
    .Q(\u_neuron.pre_trace[6] ),
    .CLK(clknet_5_11__leaf_clk));
 sg13g2_dfrbpq_1 \u_neuron.u_learning/_315_  (.RESET_B(net442),
    .D(net97),
    .Q(\u_neuron.pre_trace[7] ),
    .CLK(clknet_5_10__leaf_clk));
 sg13g2_dfrbpq_1 \u_neuron.u_learning/_316_  (.RESET_B(net443),
    .D(\u_neuron.u_learning/_008_ ),
    .Q(\u_neuron.pre_trace[8] ),
    .CLK(clknet_5_9__leaf_clk));
 sg13g2_dfrbpq_1 \u_neuron.u_learning/_317_  (.RESET_B(net442),
    .D(\u_neuron.u_learning/_009_ ),
    .Q(\u_neuron.pre_trace[9] ),
    .CLK(clknet_5_11__leaf_clk));
 sg13g2_dfrbpq_1 \u_neuron.u_learning/_318_  (.RESET_B(net442),
    .D(\u_neuron.u_learning/_010_ ),
    .Q(\u_neuron.pre_trace[10] ),
    .CLK(clknet_5_11__leaf_clk));
 sg13g2_dfrbpq_1 \u_neuron.u_learning/_319_  (.RESET_B(net443),
    .D(\u_neuron.u_learning/_011_ ),
    .Q(\u_neuron.pre_trace[11] ),
    .CLK(clknet_5_10__leaf_clk));
 sg13g2_dfrbpq_1 \u_neuron.u_learning/_320_  (.RESET_B(net441),
    .D(\u_neuron.u_learning/_012_ ),
    .Q(\u_neuron.pre_trace[12] ),
    .CLK(clknet_5_8__leaf_clk));
 sg13g2_dfrbpq_1 \u_neuron.u_learning/_321_  (.RESET_B(net441),
    .D(\u_neuron.u_learning/_013_ ),
    .Q(\u_neuron.pre_trace[13] ),
    .CLK(clknet_5_11__leaf_clk));
 sg13g2_dfrbpq_1 \u_neuron.u_learning/_322_  (.RESET_B(net443),
    .D(\u_neuron.u_learning/_014_ ),
    .Q(\u_neuron.pre_trace[14] ),
    .CLK(clknet_5_8__leaf_clk));
 sg13g2_dfrbpq_1 \u_neuron.u_learning/_323_  (.RESET_B(net444),
    .D(net214),
    .Q(\u_neuron.pre_trace[15] ),
    .CLK(clknet_5_8__leaf_clk));
 sg13g2_dfrbpq_1 \u_neuron.u_learning/_324_  (.RESET_B(net444),
    .D(\u_neuron.u_learning/_016_ ),
    .Q(\u_neuron.post_trace ),
    .CLK(clknet_5_13__leaf_clk));
 sg13g2_dfrbpq_2 \u_neuron.u_learning/_325_  (.RESET_B(net441),
    .D(net201),
    .Q(\u_neuron.learn_pending ),
    .CLK(clknet_5_8__leaf_clk));
 sg13g2_dfrbpq_2 \u_neuron.u_learning/_326_  (.RESET_B(net441),
    .D(\u_neuron.u_learning/_018_ ),
    .Q(\u_neuron.learn_ptr[0] ),
    .CLK(clknet_5_12__leaf_clk));
 sg13g2_dfrbpq_2 \u_neuron.u_learning/_327_  (.RESET_B(net441),
    .D(\u_neuron.u_learning/_019_ ),
    .Q(\u_neuron.learn_ptr[1] ),
    .CLK(clknet_5_12__leaf_clk));
 sg13g2_dfrbpq_1 \u_neuron.u_learning/_328_  (.RESET_B(net441),
    .D(\u_neuron.u_learning/_020_ ),
    .Q(\u_neuron.learn_ptr[2] ),
    .CLK(clknet_5_9__leaf_clk));
 sg13g2_dfrbpq_1 \u_neuron.u_learning/_329_  (.RESET_B(net441),
    .D(\u_neuron.u_learning/_021_ ),
    .Q(\u_neuron.learn_ptr[3] ),
    .CLK(clknet_5_12__leaf_clk));
 sg13g2_buf_8 \u_neuron.u_learning/_330_  (.A(net398),
    .X(\u_neuron.ltd_idx[0] ));
 sg13g2_buf_1 \u_neuron.u_learning/_331_  (.A(net391),
    .X(\u_neuron.ltd_idx[1] ));
 sg13g2_buf_1 \u_neuron.u_learning/_332_  (.A(net389),
    .X(\u_neuron.ltd_idx[2] ));
 sg13g2_buf_1 \u_neuron.u_learning/_333_  (.A(net386),
    .X(\u_neuron.ltd_idx[3] ));
 sg13g2_buf_2 \u_neuron.u_learning/_334_  (.A(net429),
    .X(\u_neuron.ltp_idx[0] ));
 sg13g2_buf_8 \u_neuron.u_learning/_335_  (.A(\u_neuron.learn_ptr[1] ),
    .X(\u_neuron.ltp_idx[1] ));
 sg13g2_buf_8 \u_neuron.u_learning/_336_  (.A(net423),
    .X(\u_neuron.ltp_idx[2] ));
 sg13g2_buf_8 \u_neuron.u_learning/_337_  (.A(net420),
    .X(\u_neuron.ltp_idx[3] ));
 sg13g2_inv_2 \u_neuron.u_lif/_061_  (.Y(\u_neuron.u_lif/_003_ ),
    .A(net353));
 sg13g2_inv_2 \u_neuron.u_lif/_062_  (.Y(\u_neuron.u_lif/_004_ ),
    .A(net161));
 sg13g2_inv_1 \u_neuron.u_lif/_063_  (.Y(\u_neuron.u_lif/_005_ ),
    .A(net195));
 sg13g2_inv_1 \u_neuron.u_lif/_064_  (.Y(\u_neuron.u_lif/_006_ ),
    .A(net120));
 sg13g2_inv_1 \u_neuron.u_lif/_065_  (.Y(\u_neuron.u_lif/_007_ ),
    .A(net149));
 sg13g2_nor3_1 \u_neuron.u_lif/_066_  (.A(\u_neuron.lif_V[5] ),
    .B(\u_neuron.lif_V[7] ),
    .C(\u_neuron.lif_V[6] ),
    .Y(\u_neuron.u_lif/_008_ ));
 sg13g2_inv_1 \u_neuron.u_lif/_067_  (.Y(\u_neuron.u_lif/_009_ ),
    .A(\u_neuron.u_lif/_008_ ));
 sg13g2_nand2_1 \u_neuron.u_lif/_068_  (.Y(\u_neuron.u_lif/_010_ ),
    .A(\u_neuron.w_eff[1] ),
    .B(\u_neuron.lif_V[1] ));
 sg13g2_nand2_1 \u_neuron.u_lif/_069_  (.Y(\u_neuron.u_lif/_011_ ),
    .A(\u_neuron.w_eff[0] ),
    .B(\u_neuron.lif_V[0] ));
 sg13g2_xnor2_1 \u_neuron.u_lif/_070_  (.Y(\u_neuron.u_lif/_012_ ),
    .A(\u_neuron.w_eff[1] ),
    .B(\u_neuron.lif_V[1] ));
 sg13g2_o21ai_1 \u_neuron.u_lif/_071_  (.B1(\u_neuron.u_lif/_010_ ),
    .Y(\u_neuron.u_lif/_013_ ),
    .A1(\u_neuron.u_lif/_011_ ),
    .A2(\u_neuron.u_lif/_012_ ));
 sg13g2_and3_1 \u_neuron.u_lif/_072_  (.X(\u_neuron.u_lif/_014_ ),
    .A(\u_neuron.lif_V[3] ),
    .B(\u_neuron.lif_V[2] ),
    .C(\u_neuron.u_lif/_013_ ));
 sg13g2_a21o_2 \u_neuron.u_lif/_073_  (.A2(\u_neuron.u_lif/_014_ ),
    .A1(\u_neuron.lif_V[4] ),
    .B1(\u_neuron.u_lif/_009_ ),
    .X(\u_neuron.u_lif/_015_ ));
 sg13g2_nor2_1 \u_neuron.u_lif/_074_  (.A(net417),
    .B(\u_neuron.u_lif/_003_ ),
    .Y(\u_neuron.u_lif/_016_ ));
 sg13g2_nand2_1 \u_neuron.u_lif/_075_  (.Y(\u_neuron.u_lif/_017_ ),
    .A(\u_neuron.u_lif/_015_ ),
    .B(\u_neuron.u_lif/_016_ ));
 sg13g2_nor2_2 \u_neuron.u_lif/_076_  (.A(net385),
    .B(\u_neuron.u_lif/_017_ ),
    .Y(\u_neuron.lif_post_spike ));
 sg13g2_inv_1 \u_neuron.u_lif/_077_  (.Y(\u_neuron.lif_emit_data[6] ),
    .A(\u_neuron.lif_post_spike ));
 sg13g2_nand2_1 \u_neuron.u_lif/_078_  (.Y(\u_neuron.u_lif/_018_ ),
    .A(net383),
    .B(net353));
 sg13g2_nand3_1 \u_neuron.u_lif/_079_  (.B(\u_neuron.stream_act ),
    .C(\u_neuron.u_lif/_016_ ),
    .A(net385),
    .Y(\u_neuron.u_lif/_019_ ));
 sg13g2_o21ai_1 \u_neuron.u_lif/_080_  (.B1(\u_neuron.u_lif/_019_ ),
    .Y(\u_neuron.lif_emit_valid ),
    .A1(\u_neuron.is_tick ),
    .A2(\u_neuron.u_lif/_017_ ));
 sg13g2_and2_1 \u_neuron.u_lif/_081_  (.A(\u_neuron.learn_en ),
    .B(\u_neuron.lif_post_spike ),
    .X(\u_neuron.lif_learn_start ));
 sg13g2_nor2_1 \u_neuron.u_lif/_082_  (.A(net382),
    .B(\u_neuron.u_lif/_015_ ),
    .Y(\u_neuron.u_lif/_020_ ));
 sg13g2_or2_1 \u_neuron.u_lif/_083_  (.X(\u_neuron.u_lif/_021_ ),
    .B(net142),
    .A(\u_neuron.w_eff[0] ));
 sg13g2_nand4_1 \u_neuron.u_lif/_084_  (.B(\u_neuron.u_lif/_011_ ),
    .C(\u_neuron.u_lif/_020_ ),
    .A(net353),
    .Y(\u_neuron.u_lif/_022_ ),
    .D(\u_neuron.u_lif/_021_ ));
 sg13g2_nor2b_1 \u_neuron.u_lif/_085_  (.A(\u_neuron.lif_V[3] ),
    .B_N(net383),
    .Y(\u_neuron.u_lif/_023_ ));
 sg13g2_o21ai_1 \u_neuron.u_lif/_086_  (.B1(net142),
    .Y(\u_neuron.u_lif/_024_ ),
    .A1(\u_neuron.u_lif/_003_ ),
    .A2(\u_neuron.u_lif/_023_ ));
 sg13g2_nand2b_2 \u_neuron.u_lif/_087_  (.Y(\u_neuron.u_lif/_025_ ),
    .B(\u_neuron.lif_V[3] ),
    .A_N(\u_neuron.lif_V[0] ));
 sg13g2_o21ai_1 \u_neuron.u_lif/_088_  (.B1(\u_neuron.u_lif/_024_ ),
    .Y(\u_neuron.u_lif/_026_ ),
    .A1(\u_neuron.u_lif/_018_ ),
    .A2(\u_neuron.u_lif/_025_ ));
 sg13g2_nand2b_1 \u_neuron.u_lif/_089_  (.Y(\u_neuron.lif_V_next[0] ),
    .B(\u_neuron.u_lif/_022_ ),
    .A_N(\u_neuron.u_lif/_026_ ));
 sg13g2_nor2_1 \u_neuron.u_lif/_090_  (.A(\u_neuron.mode_lif_evt ),
    .B(net173),
    .Y(\u_neuron.u_lif/_027_ ));
 sg13g2_xor2_1 \u_neuron.u_lif/_091_  (.B(\u_neuron.u_lif/_012_ ),
    .A(\u_neuron.u_lif/_011_ ),
    .X(\u_neuron.u_lif/_028_ ));
 sg13g2_nor2b_1 \u_neuron.u_lif/_092_  (.A(\u_neuron.lif_V[4] ),
    .B_N(\u_neuron.lif_V[1] ),
    .Y(\u_neuron.u_lif/_029_ ));
 sg13g2_xnor2_1 \u_neuron.u_lif/_093_  (.Y(\u_neuron.u_lif/_030_ ),
    .A(\u_neuron.lif_V[1] ),
    .B(\u_neuron.lif_V[4] ));
 sg13g2_o21ai_1 \u_neuron.u_lif/_094_  (.B1(net383),
    .Y(\u_neuron.u_lif/_031_ ),
    .A1(\u_neuron.u_lif/_025_ ),
    .A2(\u_neuron.u_lif/_030_ ));
 sg13g2_a21oi_1 \u_neuron.u_lif/_095_  (.A1(\u_neuron.u_lif/_025_ ),
    .A2(\u_neuron.u_lif/_030_ ),
    .Y(\u_neuron.u_lif/_032_ ),
    .B1(\u_neuron.u_lif/_031_ ));
 sg13g2_a21oi_1 \u_neuron.u_lif/_096_  (.A1(\u_neuron.u_lif/_020_ ),
    .A2(\u_neuron.u_lif/_028_ ),
    .Y(\u_neuron.u_lif/_033_ ),
    .B1(\u_neuron.u_lif/_032_ ));
 sg13g2_a21oi_1 \u_neuron.u_lif/_097_  (.A1(net353),
    .A2(\u_neuron.u_lif/_033_ ),
    .Y(\u_neuron.lif_V_next[1] ),
    .B1(\u_neuron.u_lif/_027_ ));
 sg13g2_nor2_1 \u_neuron.u_lif/_098_  (.A(net353),
    .B(net191),
    .Y(\u_neuron.u_lif/_034_ ));
 sg13g2_xor2_1 \u_neuron.u_lif/_099_  (.B(\u_neuron.u_lif/_013_ ),
    .A(\u_neuron.lif_V[2] ),
    .X(\u_neuron.u_lif/_035_ ));
 sg13g2_nand2_1 \u_neuron.u_lif/_100_  (.Y(\u_neuron.u_lif/_036_ ),
    .A(\u_neuron.lif_V[2] ),
    .B(\u_neuron.u_lif/_005_ ));
 sg13g2_xor2_1 \u_neuron.u_lif/_101_  (.B(\u_neuron.lif_V[5] ),
    .A(\u_neuron.lif_V[2] ),
    .X(\u_neuron.u_lif/_037_ ));
 sg13g2_a21oi_1 \u_neuron.u_lif/_102_  (.A1(\u_neuron.u_lif/_025_ ),
    .A2(\u_neuron.u_lif/_030_ ),
    .Y(\u_neuron.u_lif/_038_ ),
    .B1(\u_neuron.u_lif/_029_ ));
 sg13g2_o21ai_1 \u_neuron.u_lif/_103_  (.B1(net383),
    .Y(\u_neuron.u_lif/_039_ ),
    .A1(\u_neuron.u_lif/_037_ ),
    .A2(\u_neuron.u_lif/_038_ ));
 sg13g2_a21oi_1 \u_neuron.u_lif/_104_  (.A1(\u_neuron.u_lif/_037_ ),
    .A2(\u_neuron.u_lif/_038_ ),
    .Y(\u_neuron.u_lif/_040_ ),
    .B1(\u_neuron.u_lif/_039_ ));
 sg13g2_a21oi_1 \u_neuron.u_lif/_105_  (.A1(\u_neuron.u_lif/_020_ ),
    .A2(\u_neuron.u_lif/_035_ ),
    .Y(\u_neuron.u_lif/_041_ ),
    .B1(\u_neuron.u_lif/_040_ ));
 sg13g2_a21oi_1 \u_neuron.u_lif/_106_  (.A1(net353),
    .A2(\u_neuron.u_lif/_041_ ),
    .Y(\u_neuron.lif_V_next[2] ),
    .B1(\u_neuron.u_lif/_034_ ));
 sg13g2_o21ai_1 \u_neuron.u_lif/_107_  (.B1(\u_neuron.u_lif/_036_ ),
    .Y(\u_neuron.u_lif/_042_ ),
    .A1(\u_neuron.u_lif/_037_ ),
    .A2(\u_neuron.u_lif/_038_ ));
 sg13g2_nor2_1 \u_neuron.u_lif/_108_  (.A(\u_neuron.u_lif/_004_ ),
    .B(\u_neuron.lif_V[6] ),
    .Y(\u_neuron.u_lif/_043_ ));
 sg13g2_nand2_1 \u_neuron.u_lif/_109_  (.Y(\u_neuron.u_lif/_044_ ),
    .A(\u_neuron.u_lif/_004_ ),
    .B(\u_neuron.lif_V[6] ));
 sg13g2_nand2b_1 \u_neuron.u_lif/_110_  (.Y(\u_neuron.u_lif/_045_ ),
    .B(\u_neuron.u_lif/_044_ ),
    .A_N(\u_neuron.u_lif/_043_ ));
 sg13g2_xnor2_1 \u_neuron.u_lif/_111_  (.Y(\u_neuron.u_lif/_046_ ),
    .A(\u_neuron.u_lif/_042_ ),
    .B(\u_neuron.u_lif/_045_ ));
 sg13g2_a21oi_1 \u_neuron.u_lif/_112_  (.A1(\u_neuron.lif_V[2] ),
    .A2(\u_neuron.u_lif/_013_ ),
    .Y(\u_neuron.u_lif/_047_ ),
    .B1(\u_neuron.lif_V[3] ));
 sg13g2_or3_1 \u_neuron.u_lif/_113_  (.A(net383),
    .B(\u_neuron.u_lif/_009_ ),
    .C(\u_neuron.u_lif/_047_ ),
    .X(\u_neuron.u_lif/_048_ ));
 sg13g2_o21ai_1 \u_neuron.u_lif/_114_  (.B1(net353),
    .Y(\u_neuron.u_lif/_049_ ),
    .A1(\u_neuron.u_lif/_014_ ),
    .A2(\u_neuron.u_lif/_048_ ));
 sg13g2_a21oi_1 \u_neuron.u_lif/_115_  (.A1(net382),
    .A2(\u_neuron.u_lif/_046_ ),
    .Y(\u_neuron.u_lif/_050_ ),
    .B1(\u_neuron.u_lif/_049_ ));
 sg13g2_a21oi_1 \u_neuron.u_lif/_116_  (.A1(\u_neuron.u_lif/_003_ ),
    .A2(\u_neuron.u_lif/_004_ ),
    .Y(\u_neuron.lif_V_next[3] ),
    .B1(\u_neuron.u_lif/_050_ ));
 sg13g2_nand2_1 \u_neuron.u_lif/_117_  (.Y(\u_neuron.u_lif/_051_ ),
    .A(\u_neuron.lif_V[4] ),
    .B(\u_neuron.u_lif/_006_ ));
 sg13g2_xor2_1 \u_neuron.u_lif/_118_  (.B(\u_neuron.lif_V[7] ),
    .A(\u_neuron.lif_V[4] ),
    .X(\u_neuron.u_lif/_052_ ));
 sg13g2_a21oi_1 \u_neuron.u_lif/_119_  (.A1(\u_neuron.u_lif/_042_ ),
    .A2(\u_neuron.u_lif/_044_ ),
    .Y(\u_neuron.u_lif/_053_ ),
    .B1(\u_neuron.u_lif/_043_ ));
 sg13g2_xnor2_1 \u_neuron.u_lif/_120_  (.Y(\u_neuron.u_lif/_054_ ),
    .A(\u_neuron.u_lif/_052_ ),
    .B(\u_neuron.u_lif/_053_ ));
 sg13g2_o21ai_1 \u_neuron.u_lif/_121_  (.B1(net353),
    .Y(\u_neuron.u_lif/_055_ ),
    .A1(\u_neuron.lif_V[4] ),
    .A2(\u_neuron.u_lif/_014_ ));
 sg13g2_or2_1 \u_neuron.u_lif/_122_  (.X(\u_neuron.u_lif/_056_ ),
    .B(\u_neuron.u_lif/_055_ ),
    .A(\u_neuron.u_lif/_015_ ));
 sg13g2_a22oi_1 \u_neuron.u_lif/_123_  (.Y(\u_neuron.u_lif/_057_ ),
    .B1(\u_neuron.u_lif/_056_ ),
    .B2(\u_neuron.u_lif/_018_ ),
    .A2(\u_neuron.u_lif/_054_ ),
    .A1(net382));
 sg13g2_a21o_1 \u_neuron.u_lif/_124_  (.A2(net199),
    .A1(\u_neuron.u_lif/_003_ ),
    .B1(\u_neuron.u_lif/_057_ ),
    .X(\u_neuron.lif_V_next[4] ));
 sg13g2_o21ai_1 \u_neuron.u_lif/_125_  (.B1(\u_neuron.u_lif/_051_ ),
    .Y(\u_neuron.u_lif/_058_ ),
    .A1(\u_neuron.u_lif/_052_ ),
    .A2(\u_neuron.u_lif/_053_ ));
 sg13g2_a21oi_1 \u_neuron.u_lif/_126_  (.A1(net382),
    .A2(\u_neuron.u_lif/_058_ ),
    .Y(\u_neuron.u_lif/_059_ ),
    .B1(\u_neuron.u_lif/_003_ ));
 sg13g2_or3_1 \u_neuron.u_lif/_127_  (.A(net195),
    .B(\u_neuron.u_lif/_018_ ),
    .C(\u_neuron.u_lif/_058_ ),
    .X(\u_neuron.u_lif/_060_ ));
 sg13g2_o21ai_1 \u_neuron.u_lif/_128_  (.B1(\u_neuron.u_lif/_060_ ),
    .Y(\u_neuron.lif_V_next[5] ),
    .A1(\u_neuron.u_lif/_005_ ),
    .A2(\u_neuron.u_lif/_059_ ));
 sg13g2_o21ai_1 \u_neuron.u_lif/_129_  (.B1(net382),
    .Y(\u_neuron.u_lif/_000_ ),
    .A1(\u_neuron.lif_V[5] ),
    .A2(\u_neuron.u_lif/_058_ ));
 sg13g2_nor2_1 \u_neuron.u_lif/_130_  (.A(\u_neuron.u_lif/_003_ ),
    .B(\u_neuron.u_lif/_007_ ),
    .Y(\u_neuron.u_lif/_001_ ));
 sg13g2_a22oi_1 \u_neuron.u_lif/_131_  (.Y(\u_neuron.lif_V_next[6] ),
    .B1(\u_neuron.u_lif/_000_ ),
    .B2(\u_neuron.u_lif/_001_ ),
    .A2(\u_neuron.u_lif/_060_ ),
    .A1(\u_neuron.u_lif/_007_ ));
 sg13g2_o21ai_1 \u_neuron.u_lif/_132_  (.B1(net382),
    .Y(\u_neuron.u_lif/_002_ ),
    .A1(\u_neuron.lif_V[5] ),
    .A2(\u_neuron.lif_V[6] ));
 sg13g2_a21oi_1 \u_neuron.u_lif/_133_  (.A1(\u_neuron.u_lif/_059_ ),
    .A2(\u_neuron.u_lif/_002_ ),
    .Y(\u_neuron.lif_V_next[7] ),
    .B1(\u_neuron.u_lif/_006_ ));
 sg13g2_nor2b_1 \u_neuron.u_lif/_134_  (.A(\u_neuron.lif_post_spike ),
    .B_N(\u_neuron.lif_V[0] ),
    .Y(\u_neuron.lif_emit_data[0] ));
 sg13g2_nor2b_1 \u_neuron.u_lif/_135_  (.A(\u_neuron.lif_post_spike ),
    .B_N(\u_neuron.lif_V[1] ),
    .Y(\u_neuron.lif_emit_data[1] ));
 sg13g2_nor2b_1 \u_neuron.u_lif/_136_  (.A(\u_neuron.lif_post_spike ),
    .B_N(\u_neuron.lif_V[2] ),
    .Y(\u_neuron.lif_emit_data[2] ));
 sg13g2_nor2_1 \u_neuron.u_lif/_137_  (.A(\u_neuron.u_lif/_004_ ),
    .B(\u_neuron.lif_post_spike ),
    .Y(\u_neuron.lif_emit_data[3] ));
 sg13g2_tiehi \u_neuron.u_mode_sel/_09__42  (.L_HI(net42));
 sg13g2_tielo \u_neuron.u_mode_sel/_07__35  (.L_LO(net35));
 sg13g2_buf_1 \u_neuron.u_lif/_140_  (.A(\u_neuron.lif_emit_data[6] ),
    .X(\u_neuron.lif_emit_data[4] ));
 sg13g2_mux4_1 \u_neuron.u_mode_sel/_00_  (.S0(net433),
    .A0(\u_neuron.lif_learn_start ),
    .A1(net36),
    .A2(net33),
    .A3(net19),
    .S1(net432),
    .X(\u_neuron.mode_learn_start ));
 sg13g2_mux4_1 \u_neuron.u_mode_sel/_01_  (.S0(net433),
    .A0(\u_neuron.lif_post_spike ),
    .A1(\u_neuron.td_post_spike ),
    .A2(\u_neuron.fst_post_spike ),
    .A3(\u_neuron.conv_post_spike ),
    .S1(net431),
    .X(\u_neuron.mode_post_spike ));
 sg13g2_mux4_1 \u_neuron.u_mode_sel/_02_  (.S0(net433),
    .A0(\u_neuron.lif_emit_data[0] ),
    .A1(\u_neuron.td_emit_data[0] ),
    .A2(\u_neuron.fst_emit_data[0] ),
    .A3(\u_neuron.conv_emit_data[0] ),
    .S1(net431),
    .X(\u_neuron.mode_emit_data[0] ));
 sg13g2_mux4_1 \u_neuron.u_mode_sel/_03_  (.S0(net433),
    .A0(\u_neuron.lif_emit_data[1] ),
    .A1(\u_neuron.td_emit_data[1] ),
    .A2(\u_neuron.fst_emit_data[1] ),
    .A3(\u_neuron.conv_emit_data[1] ),
    .S1(net431),
    .X(\u_neuron.mode_emit_data[1] ));
 sg13g2_mux4_1 \u_neuron.u_mode_sel/_04_  (.S0(net433),
    .A0(\u_neuron.lif_emit_data[2] ),
    .A1(\u_neuron.td_emit_data[2] ),
    .A2(\u_neuron.fst_emit_data[2] ),
    .A3(\u_neuron.conv_emit_data[2] ),
    .S1(net431),
    .X(\u_neuron.mode_emit_data[2] ));
 sg13g2_mux4_1 \u_neuron.u_mode_sel/_05_  (.S0(net434),
    .A0(\u_neuron.lif_emit_data[3] ),
    .A1(\u_neuron.td_emit_data[3] ),
    .A2(\u_neuron.fst_emit_data[3] ),
    .A3(net17),
    .S1(\u_neuron.mode[1] ),
    .X(\u_neuron.mode_emit_data[3] ));
 sg13g2_mux4_1 \u_neuron.u_mode_sel/_06_  (.S0(net434),
    .A0(\u_neuron.lif_emit_data[4] ),
    .A1(\u_neuron.td_emit_data[4] ),
    .A2(\u_neuron.fst_emit_data[4] ),
    .A3(\u_neuron.conv_emit_data[4] ),
    .S1(net432),
    .X(\u_neuron.mode_emit_data[4] ));
 sg13g2_mux4_1 \u_neuron.u_mode_sel/_07_  (.S0(net434),
    .A0(net34),
    .A1(net35),
    .A2(net32),
    .A3(net18),
    .S1(net432),
    .X(\u_neuron.mode_emit_data[5] ));
 sg13g2_mux4_1 \u_neuron.u_mode_sel/_08_  (.S0(net434),
    .A0(\u_neuron.lif_emit_data[6] ),
    .A1(\u_neuron.td_emit_data[6] ),
    .A2(\u_neuron.fst_emit_data[6] ),
    .A3(\u_neuron.conv_emit_data[6] ),
    .S1(net432),
    .X(\u_neuron.mode_emit_data[6] ));
 sg13g2_mux4_1 \u_neuron.u_mode_sel/_09_  (.S0(net434),
    .A0(net41),
    .A1(net42),
    .A2(net40),
    .A3(net37),
    .S1(net432),
    .X(\u_neuron.mode_emit_data[7] ));
 sg13g2_mux4_1 \u_neuron.u_mode_sel/_10_  (.S0(net434),
    .A0(\u_neuron.lif_emit_valid ),
    .A1(\u_neuron.td_emit_valid ),
    .A2(\u_neuron.fst_emit_valid ),
    .A3(\u_neuron.conv_emit_valid ),
    .S1(net432),
    .X(\u_neuron.mode_emit_valid ));
 sg13g2_inv_1 \u_neuron.u_outq/_29_  (.Y(\u_neuron.u_outq/_09_ ),
    .A(net418));
 sg13g2_inv_1 \u_neuron.u_outq/_30_  (.Y(\u_neuron.u_outq/_10_ ),
    .A(\u_neuron.mode_emit_data[0] ));
 sg13g2_inv_1 \u_neuron.u_outq/_31_  (.Y(\u_neuron.u_outq/_11_ ),
    .A(\u_neuron.mode_emit_data[1] ));
 sg13g2_inv_1 \u_neuron.u_outq/_32_  (.Y(\u_neuron.u_outq/_12_ ),
    .A(\u_neuron.mode_emit_data[2] ));
 sg13g2_inv_1 \u_neuron.u_outq/_33_  (.Y(\u_neuron.u_outq/_13_ ),
    .A(\u_neuron.mode_emit_data[3] ));
 sg13g2_inv_1 \u_neuron.u_outq/_34_  (.Y(\u_neuron.u_outq/_14_ ),
    .A(\u_neuron.mode_emit_data[4] ));
 sg13g2_inv_1 \u_neuron.u_outq/_35_  (.Y(\u_neuron.u_outq/_15_ ),
    .A(\u_neuron.mode_emit_data[5] ));
 sg13g2_inv_1 \u_neuron.u_outq/_36_  (.Y(\u_neuron.u_outq/_16_ ),
    .A(\u_neuron.mode_emit_data[6] ));
 sg13g2_inv_1 \u_neuron.u_outq/_37_  (.Y(\u_neuron.u_outq/_17_ ),
    .A(\u_neuron.mode_emit_data[7] ));
 sg13g2_nand2b_1 \u_neuron.u_outq/_38_  (.Y(\u_neuron.u_outq/_18_ ),
    .B(net469),
    .A_N(\u_neuron.out_fire ));
 sg13g2_a21oi_2 \u_neuron.u_outq/_39_  (.B1(\u_neuron.u_outq/_18_ ),
    .Y(\u_neuron.u_outq/_19_ ),
    .A2(\u_neuron.mode_emit_valid ),
    .A1(\u_neuron.u_outq/_09_ ));
 sg13g2_nand3b_1 \u_neuron.u_outq/_40_  (.B(\u_neuron.mode_emit_valid ),
    .C(net469),
    .Y(\u_neuron.u_outq/_20_ ),
    .A_N(net418));
 sg13g2_nor2_1 \u_neuron.u_outq/_41_  (.A(\u_neuron.u_outq/_10_ ),
    .B(net314),
    .Y(\u_neuron.u_outq/_21_ ));
 sg13g2_a21o_1 \u_neuron.u_outq/_42_  (.A2(\u_neuron.u_outq/_19_ ),
    .A1(net180),
    .B1(\u_neuron.u_outq/_21_ ),
    .X(\u_neuron.u_outq/_00_ ));
 sg13g2_nor2_1 \u_neuron.u_outq/_43_  (.A(\u_neuron.u_outq/_11_ ),
    .B(net314),
    .Y(\u_neuron.u_outq/_22_ ));
 sg13g2_a21o_1 \u_neuron.u_outq/_44_  (.A2(\u_neuron.u_outq/_19_ ),
    .A1(net175),
    .B1(\u_neuron.u_outq/_22_ ),
    .X(\u_neuron.u_outq/_01_ ));
 sg13g2_nor2_1 \u_neuron.u_outq/_45_  (.A(\u_neuron.u_outq/_12_ ),
    .B(net314),
    .Y(\u_neuron.u_outq/_23_ ));
 sg13g2_a21o_1 \u_neuron.u_outq/_46_  (.A2(\u_neuron.u_outq/_19_ ),
    .A1(net168),
    .B1(\u_neuron.u_outq/_23_ ),
    .X(\u_neuron.u_outq/_02_ ));
 sg13g2_nor2_1 \u_neuron.u_outq/_47_  (.A(\u_neuron.u_outq/_13_ ),
    .B(\u_neuron.u_outq/_20_ ),
    .Y(\u_neuron.u_outq/_24_ ));
 sg13g2_a21o_1 \u_neuron.u_outq/_48_  (.A2(\u_neuron.u_outq/_19_ ),
    .A1(net176),
    .B1(\u_neuron.u_outq/_24_ ),
    .X(\u_neuron.u_outq/_03_ ));
 sg13g2_nor2_1 \u_neuron.u_outq/_49_  (.A(\u_neuron.u_outq/_14_ ),
    .B(net314),
    .Y(\u_neuron.u_outq/_25_ ));
 sg13g2_a21o_1 \u_neuron.u_outq/_50_  (.A2(\u_neuron.u_outq/_19_ ),
    .A1(net171),
    .B1(\u_neuron.u_outq/_25_ ),
    .X(\u_neuron.u_outq/_04_ ));
 sg13g2_nor2_1 \u_neuron.u_outq/_51_  (.A(\u_neuron.u_outq/_15_ ),
    .B(net314),
    .Y(\u_neuron.u_outq/_26_ ));
 sg13g2_a21o_1 \u_neuron.u_outq/_52_  (.A2(\u_neuron.u_outq/_19_ ),
    .A1(net167),
    .B1(\u_neuron.u_outq/_26_ ),
    .X(\u_neuron.u_outq/_05_ ));
 sg13g2_nor2_1 \u_neuron.u_outq/_53_  (.A(\u_neuron.u_outq/_16_ ),
    .B(net314),
    .Y(\u_neuron.u_outq/_27_ ));
 sg13g2_a21o_1 \u_neuron.u_outq/_54_  (.A2(\u_neuron.u_outq/_19_ ),
    .A1(net164),
    .B1(\u_neuron.u_outq/_27_ ),
    .X(\u_neuron.u_outq/_06_ ));
 sg13g2_nor2_1 \u_neuron.u_outq/_55_  (.A(\u_neuron.u_outq/_17_ ),
    .B(net314),
    .Y(\u_neuron.u_outq/_28_ ));
 sg13g2_a21o_1 \u_neuron.u_outq/_56_  (.A2(\u_neuron.u_outq/_19_ ),
    .A1(net160),
    .B1(\u_neuron.u_outq/_28_ ),
    .X(\u_neuron.u_outq/_07_ ));
 sg13g2_o21ai_1 \u_neuron.u_outq/_57_  (.B1(net314),
    .Y(\u_neuron.u_outq/_08_ ),
    .A1(\u_neuron.u_outq/_09_ ),
    .A2(\u_neuron.u_outq/_18_ ));
 sg13g2_dfrbpq_2 \u_neuron.u_outq/_58_  (.RESET_B(net454),
    .D(\u_neuron.u_outq/_00_ ),
    .Q(uo_out[0]),
    .CLK(clknet_5_18__leaf_clk));
 sg13g2_dfrbpq_1 \u_neuron.u_outq/_59_  (.RESET_B(net453),
    .D(\u_neuron.u_outq/_01_ ),
    .Q(uo_out[1]),
    .CLK(clknet_5_21__leaf_clk));
 sg13g2_dfrbpq_1 \u_neuron.u_outq/_60_  (.RESET_B(net453),
    .D(\u_neuron.u_outq/_02_ ),
    .Q(uo_out[2]),
    .CLK(clknet_5_20__leaf_clk));
 sg13g2_dfrbpq_2 \u_neuron.u_outq/_61_  (.RESET_B(net453),
    .D(net177),
    .Q(uo_out[3]),
    .CLK(clknet_5_18__leaf_clk));
 sg13g2_dfrbpq_2 \u_neuron.u_outq/_62_  (.RESET_B(net453),
    .D(\u_neuron.u_outq/_04_ ),
    .Q(uo_out[4]),
    .CLK(clknet_5_18__leaf_clk));
 sg13g2_dfrbpq_1 \u_neuron.u_outq/_63_  (.RESET_B(net453),
    .D(\u_neuron.u_outq/_05_ ),
    .Q(uo_out[5]),
    .CLK(clknet_5_23__leaf_clk));
 sg13g2_dfrbpq_2 \u_neuron.u_outq/_64_  (.RESET_B(net453),
    .D(\u_neuron.u_outq/_06_ ),
    .Q(uo_out[6]),
    .CLK(clknet_5_19__leaf_clk));
 sg13g2_dfrbpq_2 \u_neuron.u_outq/_65_  (.RESET_B(net453),
    .D(\u_neuron.u_outq/_07_ ),
    .Q(uo_out[7]),
    .CLK(clknet_5_22__leaf_clk));
 sg13g2_dfrbpq_1 \u_neuron.u_outq/_66_  (.RESET_B(net454),
    .D(net234),
    .Q(\u_neuron.have_out ),
    .CLK(clknet_5_18__leaf_clk));
 sg13g2_inv_2 \u_neuron.u_syn/_405_  (.Y(\u_neuron.u_syn/_036_ ),
    .A(net468));
 sg13g2_inv_4 \u_neuron.u_syn/_406_  (.A(net215),
    .Y(\u_neuron.u_syn/_037_ ));
 sg13g2_inv_1 \u_neuron.u_syn/_407_  (.Y(\u_neuron.u_syn/_038_ ),
    .A(net408));
 sg13g2_inv_1 \u_neuron.u_syn/_408_  (.Y(\u_neuron.u_syn/_039_ ),
    .A(net409));
 sg13g2_inv_1 \u_neuron.u_syn/_409_  (.Y(\u_neuron.u_syn/_040_ ),
    .A(net196));
 sg13g2_inv_4 \u_neuron.u_syn/_410_  (.A(\u_neuron.cfg_arg[0] ),
    .Y(\u_neuron.u_syn/_041_ ));
 sg13g2_inv_2 \u_neuron.u_syn/_411_  (.Y(\u_neuron.u_syn/_042_ ),
    .A(\u_neuron.ltp_idx[3] ));
 sg13g2_inv_4 \u_neuron.u_syn/_412_  (.A(\u_neuron.ltp_idx[2] ),
    .Y(\u_neuron.u_syn/_043_ ));
 sg13g2_inv_4 \u_neuron.u_syn/_413_  (.A(\u_neuron.ltp_wdata[0] ),
    .Y(\u_neuron.u_syn/_044_ ));
 sg13g2_inv_1 \u_neuron.u_syn/_414_  (.Y(\u_neuron.u_syn/_045_ ),
    .A(net321));
 sg13g2_inv_4 \u_neuron.u_syn/_415_  (.A(\u_neuron.ltd_idx[1] ),
    .Y(\u_neuron.u_syn/_046_ ));
 sg13g2_inv_1 \u_neuron.u_syn/_416_  (.Y(\u_neuron.u_syn/_047_ ),
    .A(\u_neuron.ltd_idx[0] ));
 sg13g2_inv_1 \u_neuron.u_syn/_417_  (.Y(\u_neuron.u_syn/_048_ ),
    .A(\u_neuron.ltd_idx[3] ));
 sg13g2_inv_1 \u_neuron.u_syn/_418_  (.Y(\u_neuron.u_syn/_049_ ),
    .A(net332));
 sg13g2_inv_1 \u_neuron.u_syn/_419_  (.Y(\u_neuron.u_syn/_050_ ),
    .A(net188));
 sg13g2_inv_4 \u_neuron.u_syn/_420_  (.A(\u_neuron.cfg_arg[1] ),
    .Y(\u_neuron.u_syn/_051_ ));
 sg13g2_inv_2 \u_neuron.u_syn/_421_  (.Y(\u_neuron.u_syn/_052_ ),
    .A(\u_neuron.ltp_wdata[1] ));
 sg13g2_inv_1 \u_neuron.u_syn/_422_  (.Y(\u_neuron.u_syn/_053_ ),
    .A(net331));
 sg13g2_inv_1 \u_neuron.u_syn/_423_  (.Y(\u_neuron.u_syn/_054_ ),
    .A(net225));
 sg13g2_inv_1 \u_neuron.u_syn/_424_  (.Y(\u_neuron.u_syn/_055_ ),
    .A(net169));
 sg13g2_inv_2 \u_neuron.u_syn/_425_  (.Y(\u_neuron.u_syn/_056_ ),
    .A(net217));
 sg13g2_inv_1 \u_neuron.u_syn/_426_  (.Y(\u_neuron.u_syn/_057_ ),
    .A(net202));
 sg13g2_inv_1 \u_neuron.u_syn/_427_  (.Y(\u_neuron.u_syn/_058_ ),
    .A(\u_neuron.wtab[6] ));
 sg13g2_inv_1 \u_neuron.u_syn/_428_  (.Y(\u_neuron.u_syn/_059_ ),
    .A(net179));
 sg13g2_inv_1 \u_neuron.u_syn/_429_  (.Y(\u_neuron.u_syn/_060_ ),
    .A(net184));
 sg13g2_inv_1 \u_neuron.u_syn/_430_  (.Y(\u_neuron.u_syn/_061_ ),
    .A(net207));
 sg13g2_inv_1 \u_neuron.u_syn/_431_  (.Y(\u_neuron.u_syn/_062_ ),
    .A(net172));
 sg13g2_inv_1 \u_neuron.u_syn/_432_  (.Y(\u_neuron.u_syn/_063_ ),
    .A(net186));
 sg13g2_inv_1 \u_neuron.u_syn/_433_  (.Y(\u_neuron.u_syn/_064_ ),
    .A(net111));
 sg13g2_inv_1 \u_neuron.u_syn/_434_  (.Y(\u_neuron.u_syn/_065_ ),
    .A(net205));
 sg13g2_inv_1 \u_neuron.u_syn/_435_  (.Y(\u_neuron.u_syn/_066_ ),
    .A(net204));
 sg13g2_inv_1 \u_neuron.u_syn/_436_  (.Y(\u_neuron.u_syn/_067_ ),
    .A(\u_neuron.wtab[19] ));
 sg13g2_inv_1 \u_neuron.u_syn/_437_  (.Y(\u_neuron.u_syn/_068_ ),
    .A(net185));
 sg13g2_inv_1 \u_neuron.u_syn/_438_  (.Y(\u_neuron.u_syn/_069_ ),
    .A(net208));
 sg13g2_inv_1 \u_neuron.u_syn/_439_  (.Y(\u_neuron.u_syn/_070_ ),
    .A(net148));
 sg13g2_inv_1 \u_neuron.u_syn/_440_  (.Y(\u_neuron.u_syn/_071_ ),
    .A(net147));
 sg13g2_inv_1 \u_neuron.u_syn/_441_  (.Y(\u_neuron.u_syn/_072_ ),
    .A(net197));
 sg13g2_inv_1 \u_neuron.u_syn/_442_  (.Y(\u_neuron.u_syn/_073_ ),
    .A(net198));
 sg13g2_inv_1 \u_neuron.u_syn/_443_  (.Y(\u_neuron.u_syn/_074_ ),
    .A(net189));
 sg13g2_inv_1 \u_neuron.u_syn/_444_  (.Y(\u_neuron.u_syn/_075_ ),
    .A(net211));
 sg13g2_inv_1 \u_neuron.u_syn/_445_  (.Y(\u_neuron.u_syn/_076_ ),
    .A(net194));
 sg13g2_inv_2 \u_neuron.u_syn/_446_  (.Y(\u_neuron.u_syn/_077_ ),
    .A(net391));
 sg13g2_inv_4 \u_neuron.u_syn/_447_  (.A(net390),
    .Y(\u_neuron.u_syn/_078_ ));
 sg13g2_nor2_2 \u_neuron.u_syn/_448_  (.A(\u_neuron.addr[5] ),
    .B(\u_neuron.addr[4] ),
    .Y(\u_neuron.is_prog_addr ));
 sg13g2_nand2_1 \u_neuron.u_syn/_449_  (.Y(\u_neuron.u_syn/_079_ ),
    .A(\u_neuron.wtab[6] ),
    .B(net400));
 sg13g2_o21ai_1 \u_neuron.u_syn/_450_  (.B1(\u_neuron.u_syn/_079_ ),
    .Y(\u_neuron.u_syn/_080_ ),
    .A1(\u_neuron.u_syn/_056_ ),
    .A2(net400));
 sg13g2_mux2_1 \u_neuron.u_syn/_451_  (.A0(\u_neuron.u_syn/_040_ ),
    .A1(\u_neuron.u_syn/_054_ ),
    .S(net401),
    .X(\u_neuron.u_syn/_081_ ));
 sg13g2_o21ai_1 \u_neuron.u_syn/_452_  (.B1(\u_neuron.u_syn/_078_ ),
    .Y(\u_neuron.u_syn/_082_ ),
    .A1(net394),
    .A2(\u_neuron.u_syn/_081_ ));
 sg13g2_a21oi_1 \u_neuron.u_syn/_453_  (.A1(net394),
    .A2(\u_neuron.u_syn/_080_ ),
    .Y(\u_neuron.u_syn/_083_ ),
    .B1(\u_neuron.u_syn/_082_ ));
 sg13g2_nand2_1 \u_neuron.u_syn/_454_  (.Y(\u_neuron.u_syn/_084_ ),
    .A(\u_neuron.wtab[14] ),
    .B(net400));
 sg13g2_o21ai_1 \u_neuron.u_syn/_455_  (.B1(\u_neuron.u_syn/_084_ ),
    .Y(\u_neuron.u_syn/_085_ ),
    .A1(\u_neuron.u_syn/_061_ ),
    .A2(net400));
 sg13g2_nor2b_1 \u_neuron.u_syn/_456_  (.A(net402),
    .B_N(\u_neuron.wtab[8] ),
    .Y(\u_neuron.u_syn/_086_ ));
 sg13g2_a21oi_1 \u_neuron.u_syn/_457_  (.A1(\u_neuron.wtab[10] ),
    .A2(net402),
    .Y(\u_neuron.u_syn/_087_ ),
    .B1(\u_neuron.u_syn/_086_ ));
 sg13g2_o21ai_1 \u_neuron.u_syn/_458_  (.B1(net390),
    .Y(\u_neuron.u_syn/_088_ ),
    .A1(net394),
    .A2(\u_neuron.u_syn/_087_ ));
 sg13g2_a21oi_1 \u_neuron.u_syn/_459_  (.A1(net394),
    .A2(\u_neuron.u_syn/_085_ ),
    .Y(\u_neuron.u_syn/_089_ ),
    .B1(\u_neuron.u_syn/_088_ ));
 sg13g2_or3_1 \u_neuron.u_syn/_460_  (.A(net387),
    .B(\u_neuron.u_syn/_083_ ),
    .C(\u_neuron.u_syn/_089_ ),
    .X(\u_neuron.u_syn/_090_ ));
 sg13g2_mux4_1 \u_neuron.u_syn/_461_  (.S0(net398),
    .A0(\u_neuron.wtab[16] ),
    .A1(\u_neuron.wtab[18] ),
    .A2(\u_neuron.wtab[20] ),
    .A3(\u_neuron.wtab[22] ),
    .S1(net391),
    .X(\u_neuron.u_syn/_091_ ));
 sg13g2_mux2_1 \u_neuron.u_syn/_462_  (.A0(\u_neuron.u_syn/_074_ ),
    .A1(\u_neuron.u_syn/_076_ ),
    .S(net396),
    .X(\u_neuron.u_syn/_092_ ));
 sg13g2_mux2_1 \u_neuron.u_syn/_463_  (.A0(\u_neuron.wtab[24] ),
    .A1(\u_neuron.wtab[26] ),
    .S(net396),
    .X(\u_neuron.u_syn/_093_ ));
 sg13g2_a21oi_1 \u_neuron.u_syn/_464_  (.A1(\u_neuron.u_syn/_077_ ),
    .A2(\u_neuron.u_syn/_093_ ),
    .Y(\u_neuron.u_syn/_094_ ),
    .B1(\u_neuron.u_syn/_078_ ));
 sg13g2_o21ai_1 \u_neuron.u_syn/_465_  (.B1(\u_neuron.u_syn/_094_ ),
    .Y(\u_neuron.u_syn/_095_ ),
    .A1(\u_neuron.u_syn/_077_ ),
    .A2(\u_neuron.u_syn/_092_ ));
 sg13g2_o21ai_1 \u_neuron.u_syn/_466_  (.B1(net387),
    .Y(\u_neuron.u_syn/_096_ ),
    .A1(net388),
    .A2(\u_neuron.u_syn/_091_ ));
 sg13g2_nand2b_1 \u_neuron.u_syn/_467_  (.Y(\u_neuron.u_syn/_097_ ),
    .B(\u_neuron.u_syn/_095_ ),
    .A_N(\u_neuron.u_syn/_096_ ));
 sg13g2_and2_1 \u_neuron.u_syn/_468_  (.A(\u_neuron.is_prog_addr ),
    .B(\u_neuron.u_syn/_097_ ),
    .X(\u_neuron.u_syn/_098_ ));
 sg13g2_xor2_1 \u_neuron.u_syn/_469_  (.B(net394),
    .A(\u_neuron.addr[5] ),
    .X(\u_neuron.u_syn/_099_ ));
 sg13g2_xnor2_1 \u_neuron.u_syn/_470_  (.Y(\u_neuron.u_syn/_100_ ),
    .A(net387),
    .B(\u_neuron.u_syn/_099_ ));
 sg13g2_xnor2_1 \u_neuron.u_syn/_471_  (.Y(\u_neuron.u_syn/_101_ ),
    .A(\u_neuron.addr[5] ),
    .B(net403));
 sg13g2_or2_1 \u_neuron.u_syn/_472_  (.X(\u_neuron.u_syn/_102_ ),
    .B(\u_neuron.u_syn/_101_ ),
    .A(net390));
 sg13g2_a21oi_1 \u_neuron.u_syn/_473_  (.A1(net390),
    .A2(\u_neuron.u_syn/_101_ ),
    .Y(\u_neuron.u_syn/_103_ ),
    .B1(\u_neuron.polarity ));
 sg13g2_a221oi_1 \u_neuron.u_syn/_474_  (.B2(\u_neuron.u_syn/_103_ ),
    .C1(\u_neuron.is_prog_addr ),
    .B1(\u_neuron.u_syn/_102_ ),
    .A1(\u_neuron.polarity ),
    .Y(\u_neuron.u_syn/_104_ ),
    .A2(\u_neuron.u_syn/_100_ ));
 sg13g2_nor2_1 \u_neuron.u_syn/_475_  (.A(net403),
    .B(\u_neuron.polarity ),
    .Y(\u_neuron.u_syn/_105_ ));
 sg13g2_a21oi_1 \u_neuron.u_syn/_476_  (.A1(\u_neuron.u_syn/_078_ ),
    .A2(\u_neuron.polarity ),
    .Y(\u_neuron.u_syn/_106_ ),
    .B1(\u_neuron.u_syn/_105_ ));
 sg13g2_xor2_1 \u_neuron.u_syn/_477_  (.B(net394),
    .A(\u_neuron.addr[4] ),
    .X(\u_neuron.u_syn/_107_ ));
 sg13g2_xnor2_1 \u_neuron.u_syn/_478_  (.Y(\u_neuron.u_syn/_108_ ),
    .A(\u_neuron.u_syn/_106_ ),
    .B(\u_neuron.u_syn/_107_ ));
 sg13g2_a22oi_1 \u_neuron.u_syn/_479_  (.Y(\u_neuron.w_eff[0] ),
    .B1(\u_neuron.u_syn/_104_ ),
    .B2(\u_neuron.u_syn/_108_ ),
    .A2(\u_neuron.u_syn/_098_ ),
    .A1(\u_neuron.u_syn/_090_ ));
 sg13g2_mux4_1 \u_neuron.u_syn/_480_  (.S0(net398),
    .A0(\u_neuron.u_syn/_065_ ),
    .A1(\u_neuron.u_syn/_067_ ),
    .A2(\u_neuron.u_syn/_069_ ),
    .A3(\u_neuron.u_syn/_071_ ),
    .S1(net391),
    .X(\u_neuron.u_syn/_109_ ));
 sg13g2_nor2b_1 \u_neuron.u_syn/_481_  (.A(\u_neuron.wtab[27] ),
    .B_N(net397),
    .Y(\u_neuron.u_syn/_110_ ));
 sg13g2_nor2_1 \u_neuron.u_syn/_482_  (.A(\u_neuron.wtab[25] ),
    .B(net397),
    .Y(\u_neuron.u_syn/_111_ ));
 sg13g2_nor3_1 \u_neuron.u_syn/_483_  (.A(net392),
    .B(\u_neuron.u_syn/_110_ ),
    .C(\u_neuron.u_syn/_111_ ),
    .Y(\u_neuron.u_syn/_112_ ));
 sg13g2_nor2b_1 \u_neuron.u_syn/_484_  (.A(\u_neuron.wtab[31] ),
    .B_N(net396),
    .Y(\u_neuron.u_syn/_113_ ));
 sg13g2_o21ai_1 \u_neuron.u_syn/_485_  (.B1(net392),
    .Y(\u_neuron.u_syn/_114_ ),
    .A1(\u_neuron.wtab[29] ),
    .A2(net396));
 sg13g2_o21ai_1 \u_neuron.u_syn/_486_  (.B1(net388),
    .Y(\u_neuron.u_syn/_115_ ),
    .A1(\u_neuron.u_syn/_113_ ),
    .A2(\u_neuron.u_syn/_114_ ));
 sg13g2_o21ai_1 \u_neuron.u_syn/_487_  (.B1(net386),
    .Y(\u_neuron.u_syn/_116_ ),
    .A1(\u_neuron.u_syn/_112_ ),
    .A2(\u_neuron.u_syn/_115_ ));
 sg13g2_a21oi_1 \u_neuron.u_syn/_488_  (.A1(\u_neuron.u_syn/_078_ ),
    .A2(\u_neuron.u_syn/_109_ ),
    .Y(\u_neuron.u_syn/_117_ ),
    .B1(\u_neuron.u_syn/_116_ ));
 sg13g2_mux4_1 \u_neuron.u_syn/_489_  (.S0(net403),
    .A0(\u_neuron.wtab[1] ),
    .A1(\u_neuron.wtab[3] ),
    .A2(\u_neuron.wtab[5] ),
    .A3(\u_neuron.wtab[7] ),
    .S1(net395),
    .X(\u_neuron.u_syn/_118_ ));
 sg13g2_inv_1 \u_neuron.u_syn/_490_  (.Y(\u_neuron.u_syn/_119_ ),
    .A(\u_neuron.u_syn/_118_ ));
 sg13g2_a21oi_1 \u_neuron.u_syn/_491_  (.A1(\u_neuron.u_syn/_064_ ),
    .A2(net400),
    .Y(\u_neuron.u_syn/_120_ ),
    .B1(\u_neuron.u_syn/_077_ ));
 sg13g2_o21ai_1 \u_neuron.u_syn/_492_  (.B1(\u_neuron.u_syn/_120_ ),
    .Y(\u_neuron.u_syn/_121_ ),
    .A1(\u_neuron.wtab[13] ),
    .A2(net401));
 sg13g2_or2_1 \u_neuron.u_syn/_493_  (.X(\u_neuron.u_syn/_122_ ),
    .B(net402),
    .A(\u_neuron.wtab[9] ));
 sg13g2_a21oi_1 \u_neuron.u_syn/_494_  (.A1(\u_neuron.u_syn/_060_ ),
    .A2(net402),
    .Y(\u_neuron.u_syn/_123_ ),
    .B1(net394));
 sg13g2_a21oi_1 \u_neuron.u_syn/_495_  (.A1(\u_neuron.u_syn/_122_ ),
    .A2(\u_neuron.u_syn/_123_ ),
    .Y(\u_neuron.u_syn/_124_ ),
    .B1(\u_neuron.u_syn/_078_ ));
 sg13g2_a221oi_1 \u_neuron.u_syn/_496_  (.B2(\u_neuron.u_syn/_124_ ),
    .C1(net387),
    .B1(\u_neuron.u_syn/_121_ ),
    .A1(\u_neuron.u_syn/_078_ ),
    .Y(\u_neuron.u_syn/_125_ ),
    .A2(\u_neuron.u_syn/_119_ ));
 sg13g2_o21ai_1 \u_neuron.u_syn/_497_  (.B1(\u_neuron.is_prog_addr ),
    .Y(\u_neuron.u_syn/_126_ ),
    .A1(\u_neuron.u_syn/_117_ ),
    .A2(\u_neuron.u_syn/_125_ ));
 sg13g2_nand2b_2 \u_neuron.u_syn/_498_  (.Y(\u_neuron.w_eff[1] ),
    .B(\u_neuron.u_syn/_126_ ),
    .A_N(\u_neuron.u_syn/_104_ ));
 sg13g2_nor3_1 \u_neuron.u_syn/_499_  (.A(net367),
    .B(\u_neuron.ltd_idx[1] ),
    .C(\u_neuron.ltd_idx[0] ),
    .Y(\u_neuron.u_syn/_127_ ));
 sg13g2_and3_2 \u_neuron.u_syn/_500_  (.X(\u_neuron.u_syn/_128_ ),
    .A(\u_neuron.u_syn/_048_ ),
    .B(\u_neuron.ltd_we ),
    .C(\u_neuron.u_syn/_127_ ));
 sg13g2_nor2_1 \u_neuron.u_syn/_501_  (.A(net408),
    .B(net409),
    .Y(\u_neuron.u_syn/_129_ ));
 sg13g2_nor3_2 \u_neuron.u_syn/_502_  (.A(net406),
    .B(net408),
    .C(net409),
    .Y(\u_neuron.u_syn/_130_ ));
 sg13g2_nor4_1 \u_neuron.u_syn/_503_  (.A(\u_neuron.pending_widx[3] ),
    .B(net406),
    .C(net408),
    .D(\u_neuron.pending_widx[0] ),
    .Y(\u_neuron.u_syn/_131_ ));
 sg13g2_nand2_1 \u_neuron.u_syn/_504_  (.Y(\u_neuron.u_syn/_132_ ),
    .A(net360),
    .B(\u_neuron.u_syn/_131_ ));
 sg13g2_nor3_2 \u_neuron.u_syn/_505_  (.A(\u_neuron.ltp_idx[2] ),
    .B(\u_neuron.ltp_idx[1] ),
    .C(\u_neuron.ltp_idx[0] ),
    .Y(\u_neuron.u_syn/_133_ ));
 sg13g2_nand2_1 \u_neuron.u_syn/_506_  (.Y(\u_neuron.u_syn/_134_ ),
    .A(\u_neuron.u_syn/_042_ ),
    .B(\u_neuron.u_syn/_133_ ));
 sg13g2_nand3_1 \u_neuron.u_syn/_507_  (.B(net321),
    .C(\u_neuron.u_syn/_133_ ),
    .A(\u_neuron.u_syn/_042_ ),
    .Y(\u_neuron.u_syn/_135_ ));
 sg13g2_mux2_1 \u_neuron.u_syn/_508_  (.A0(\u_neuron.cfg_arg[0] ),
    .A1(\u_neuron.wtab[0] ),
    .S(\u_neuron.u_syn/_132_ ),
    .X(\u_neuron.u_syn/_136_ ));
 sg13g2_mux2_1 \u_neuron.u_syn/_509_  (.A0(\u_neuron.ltp_wdata[0] ),
    .A1(\u_neuron.u_syn/_136_ ),
    .S(\u_neuron.u_syn/_135_ ),
    .X(\u_neuron.u_syn/_137_ ));
 sg13g2_a21oi_1 \u_neuron.u_syn/_510_  (.A1(\u_neuron.u_syn/_049_ ),
    .A2(\u_neuron.u_syn/_128_ ),
    .Y(\u_neuron.u_syn/_138_ ),
    .B1(net411));
 sg13g2_o21ai_1 \u_neuron.u_syn/_511_  (.B1(\u_neuron.u_syn/_138_ ),
    .Y(\u_neuron.u_syn/_139_ ),
    .A1(\u_neuron.u_syn/_128_ ),
    .A2(\u_neuron.u_syn/_137_ ));
 sg13g2_o21ai_1 \u_neuron.u_syn/_512_  (.B1(\u_neuron.u_syn/_139_ ),
    .Y(\u_neuron.u_syn/_000_ ),
    .A1(net466),
    .A2(\u_neuron.u_syn/_040_ ));
 sg13g2_mux2_1 \u_neuron.u_syn/_513_  (.A0(\u_neuron.cfg_arg[1] ),
    .A1(\u_neuron.wtab[1] ),
    .S(\u_neuron.u_syn/_132_ ),
    .X(\u_neuron.u_syn/_140_ ));
 sg13g2_mux2_1 \u_neuron.u_syn/_514_  (.A0(\u_neuron.ltp_wdata[1] ),
    .A1(\u_neuron.u_syn/_140_ ),
    .S(\u_neuron.u_syn/_135_ ),
    .X(\u_neuron.u_syn/_141_ ));
 sg13g2_a21oi_1 \u_neuron.u_syn/_515_  (.A1(\u_neuron.u_syn/_053_ ),
    .A2(\u_neuron.u_syn/_128_ ),
    .Y(\u_neuron.u_syn/_142_ ),
    .B1(net411));
 sg13g2_o21ai_1 \u_neuron.u_syn/_516_  (.B1(\u_neuron.u_syn/_142_ ),
    .Y(\u_neuron.u_syn/_143_ ),
    .A1(\u_neuron.u_syn/_128_ ),
    .A2(\u_neuron.u_syn/_141_ ));
 sg13g2_o21ai_1 \u_neuron.u_syn/_517_  (.B1(\u_neuron.u_syn/_143_ ),
    .Y(\u_neuron.u_syn/_001_ ),
    .A1(net468),
    .A2(\u_neuron.u_syn/_050_ ));
 sg13g2_xnor2_1 \u_neuron.u_syn/_518_  (.Y(\u_neuron.u_syn/_144_ ),
    .A(\u_neuron.pending_widx[3] ),
    .B(\u_neuron.u_syn/_130_ ));
 sg13g2_xnor2_1 \u_neuron.u_syn/_519_  (.Y(\u_neuron.u_syn/_145_ ),
    .A(\u_neuron.u_syn/_037_ ),
    .B(\u_neuron.u_syn/_130_ ));
 sg13g2_and2_1 \u_neuron.u_syn/_520_  (.A(net357),
    .B(\u_neuron.u_syn/_144_ ),
    .X(\u_neuron.u_syn/_146_ ));
 sg13g2_nand2_2 \u_neuron.u_syn/_521_  (.Y(\u_neuron.u_syn/_147_ ),
    .A(net359),
    .B(\u_neuron.u_syn/_144_ ));
 sg13g2_nor2b_2 \u_neuron.u_syn/_522_  (.A(\u_neuron.pending_widx[1] ),
    .B_N(net409),
    .Y(\u_neuron.u_syn/_148_ ));
 sg13g2_nor2b_2 \u_neuron.u_syn/_523_  (.A(net405),
    .B_N(\u_neuron.u_syn/_148_ ),
    .Y(\u_neuron.u_syn/_149_ ));
 sg13g2_nand3_1 \u_neuron.u_syn/_524_  (.B(\u_neuron.u_syn/_144_ ),
    .C(\u_neuron.u_syn/_149_ ),
    .A(net359),
    .Y(\u_neuron.u_syn/_150_ ));
 sg13g2_xnor2_1 \u_neuron.u_syn/_525_  (.Y(\u_neuron.u_syn/_151_ ),
    .A(\u_neuron.ltp_idx[3] ),
    .B(\u_neuron.u_syn/_133_ ));
 sg13g2_and2_1 \u_neuron.u_syn/_526_  (.A(net321),
    .B(\u_neuron.u_syn/_151_ ),
    .X(\u_neuron.u_syn/_152_ ));
 sg13g2_nor2b_2 \u_neuron.u_syn/_527_  (.A(\u_neuron.ltp_idx[1] ),
    .B_N(\u_neuron.ltp_idx[0] ),
    .Y(\u_neuron.u_syn/_153_ ));
 sg13g2_and2_1 \u_neuron.u_syn/_528_  (.A(\u_neuron.u_syn/_043_ ),
    .B(\u_neuron.u_syn/_153_ ),
    .X(\u_neuron.u_syn/_154_ ));
 sg13g2_nand2_1 \u_neuron.u_syn/_529_  (.Y(\u_neuron.u_syn/_155_ ),
    .A(\u_neuron.u_syn/_043_ ),
    .B(\u_neuron.u_syn/_153_ ));
 sg13g2_nand3_1 \u_neuron.u_syn/_530_  (.B(\u_neuron.u_syn/_151_ ),
    .C(\u_neuron.u_syn/_154_ ),
    .A(net321),
    .Y(\u_neuron.u_syn/_156_ ));
 sg13g2_and2_1 \u_neuron.u_syn/_531_  (.A(\u_neuron.cfg_arg[0] ),
    .B(\u_neuron.u_syn/_149_ ),
    .X(\u_neuron.u_syn/_157_ ));
 sg13g2_a22oi_1 \u_neuron.u_syn/_532_  (.Y(\u_neuron.u_syn/_158_ ),
    .B1(\u_neuron.u_syn/_157_ ),
    .B2(\u_neuron.u_syn/_146_ ),
    .A2(\u_neuron.u_syn/_150_ ),
    .A1(net225));
 sg13g2_xnor2_1 \u_neuron.u_syn/_533_  (.Y(\u_neuron.u_syn/_159_ ),
    .A(\u_neuron.ltd_idx[3] ),
    .B(\u_neuron.u_syn/_127_ ));
 sg13g2_and2_1 \u_neuron.u_syn/_534_  (.A(\u_neuron.ltd_we ),
    .B(\u_neuron.u_syn/_159_ ),
    .X(\u_neuron.u_syn/_160_ ));
 sg13g2_nand2_2 \u_neuron.u_syn/_535_  (.Y(\u_neuron.u_syn/_161_ ),
    .A(\u_neuron.ltd_we ),
    .B(\u_neuron.u_syn/_159_ ));
 sg13g2_nor2b_1 \u_neuron.u_syn/_536_  (.A(\u_neuron.ltd_idx[1] ),
    .B_N(\u_neuron.ltd_idx[0] ),
    .Y(\u_neuron.u_syn/_162_ ));
 sg13g2_nor2b_2 \u_neuron.u_syn/_537_  (.A(net367),
    .B_N(\u_neuron.u_syn/_162_ ),
    .Y(\u_neuron.u_syn/_163_ ));
 sg13g2_nand3_1 \u_neuron.u_syn/_538_  (.B(\u_neuron.u_syn/_159_ ),
    .C(\u_neuron.u_syn/_163_ ),
    .A(\u_neuron.ltd_we ),
    .Y(\u_neuron.u_syn/_164_ ));
 sg13g2_o21ai_1 \u_neuron.u_syn/_539_  (.B1(\u_neuron.u_syn/_164_ ),
    .Y(\u_neuron.u_syn/_165_ ),
    .A1(\u_neuron.ltp_wdata[0] ),
    .A2(\u_neuron.u_syn/_156_ ));
 sg13g2_a21o_1 \u_neuron.u_syn/_540_  (.A2(\u_neuron.u_syn/_158_ ),
    .A1(\u_neuron.u_syn/_156_ ),
    .B1(\u_neuron.u_syn/_165_ ),
    .X(\u_neuron.u_syn/_166_ ));
 sg13g2_and2_1 \u_neuron.u_syn/_541_  (.A(net332),
    .B(\u_neuron.u_syn/_163_ ),
    .X(\u_neuron.u_syn/_167_ ));
 sg13g2_a21oi_1 \u_neuron.u_syn/_542_  (.A1(net320),
    .A2(\u_neuron.u_syn/_167_ ),
    .Y(\u_neuron.u_syn/_168_ ),
    .B1(net416));
 sg13g2_a22oi_1 \u_neuron.u_syn/_543_  (.Y(\u_neuron.u_syn/_002_ ),
    .B1(\u_neuron.u_syn/_166_ ),
    .B2(\u_neuron.u_syn/_168_ ),
    .A2(\u_neuron.u_syn/_054_ ),
    .A1(net416));
 sg13g2_nand2b_1 \u_neuron.u_syn/_544_  (.Y(\u_neuron.u_syn/_169_ ),
    .B(\u_neuron.u_syn/_051_ ),
    .A_N(\u_neuron.u_syn/_150_ ));
 sg13g2_a22oi_1 \u_neuron.u_syn/_545_  (.Y(\u_neuron.u_syn/_170_ ),
    .B1(\u_neuron.u_syn/_152_ ),
    .B2(\u_neuron.u_syn/_154_ ),
    .A2(\u_neuron.u_syn/_150_ ),
    .A1(\u_neuron.u_syn/_055_ ));
 sg13g2_o21ai_1 \u_neuron.u_syn/_546_  (.B1(\u_neuron.u_syn/_164_ ),
    .Y(\u_neuron.u_syn/_171_ ),
    .A1(\u_neuron.u_syn/_052_ ),
    .A2(\u_neuron.u_syn/_156_ ));
 sg13g2_a21oi_1 \u_neuron.u_syn/_547_  (.A1(\u_neuron.u_syn/_169_ ),
    .A2(\u_neuron.u_syn/_170_ ),
    .Y(\u_neuron.u_syn/_172_ ),
    .B1(\u_neuron.u_syn/_171_ ));
 sg13g2_o21ai_1 \u_neuron.u_syn/_548_  (.B1(net468),
    .Y(\u_neuron.u_syn/_173_ ),
    .A1(\u_neuron.ltd_wdata[1] ),
    .A2(\u_neuron.u_syn/_164_ ));
 sg13g2_nand2_1 \u_neuron.u_syn/_549_  (.Y(\u_neuron.u_syn/_174_ ),
    .A(net416),
    .B(net169));
 sg13g2_o21ai_1 \u_neuron.u_syn/_550_  (.B1(\u_neuron.u_syn/_174_ ),
    .Y(\u_neuron.u_syn/_003_ ),
    .A1(\u_neuron.u_syn/_172_ ),
    .A2(\u_neuron.u_syn/_173_ ));
 sg13g2_nor2b_1 \u_neuron.u_syn/_551_  (.A(net409),
    .B_N(net408),
    .Y(\u_neuron.u_syn/_175_ ));
 sg13g2_nor2b_1 \u_neuron.u_syn/_552_  (.A(net404),
    .B_N(\u_neuron.u_syn/_175_ ),
    .Y(\u_neuron.u_syn/_176_ ));
 sg13g2_nand3_1 \u_neuron.u_syn/_553_  (.B(\u_neuron.u_syn/_144_ ),
    .C(\u_neuron.u_syn/_176_ ),
    .A(net357),
    .Y(\u_neuron.u_syn/_177_ ));
 sg13g2_nand2b_2 \u_neuron.u_syn/_554_  (.Y(\u_neuron.u_syn/_178_ ),
    .B(\u_neuron.ltp_idx[1] ),
    .A_N(\u_neuron.ltp_idx[0] ));
 sg13g2_nor2_1 \u_neuron.u_syn/_555_  (.A(\u_neuron.ltp_idx[2] ),
    .B(\u_neuron.u_syn/_178_ ),
    .Y(\u_neuron.u_syn/_179_ ));
 sg13g2_and3_2 \u_neuron.u_syn/_556_  (.X(\u_neuron.u_syn/_180_ ),
    .A(net321),
    .B(\u_neuron.u_syn/_151_ ),
    .C(\u_neuron.u_syn/_179_ ));
 sg13g2_nor4_1 \u_neuron.u_syn/_557_  (.A(net406),
    .B(\u_neuron.u_syn/_038_ ),
    .C(net409),
    .D(\u_neuron.u_syn/_041_ ),
    .Y(\u_neuron.u_syn/_181_ ));
 sg13g2_a221oi_1 \u_neuron.u_syn/_558_  (.B2(\u_neuron.u_syn/_146_ ),
    .C1(\u_neuron.u_syn/_180_ ),
    .B1(\u_neuron.u_syn/_181_ ),
    .A1(net217),
    .Y(\u_neuron.u_syn/_182_ ),
    .A2(\u_neuron.u_syn/_177_ ));
 sg13g2_nand2_2 \u_neuron.u_syn/_559_  (.Y(\u_neuron.u_syn/_183_ ),
    .A(\u_neuron.ltp_wdata[0] ),
    .B(\u_neuron.u_syn/_134_ ));
 sg13g2_nor2_1 \u_neuron.u_syn/_560_  (.A(\u_neuron.u_syn/_046_ ),
    .B(\u_neuron.ltd_idx[0] ),
    .Y(\u_neuron.u_syn/_184_ ));
 sg13g2_nor3_2 \u_neuron.u_syn/_561_  (.A(net367),
    .B(\u_neuron.u_syn/_046_ ),
    .C(\u_neuron.ltd_idx[0] ),
    .Y(\u_neuron.u_syn/_185_ ));
 sg13g2_a22oi_1 \u_neuron.u_syn/_562_  (.Y(\u_neuron.u_syn/_186_ ),
    .B1(\u_neuron.u_syn/_185_ ),
    .B2(net319),
    .A2(\u_neuron.u_syn/_183_ ),
    .A1(\u_neuron.u_syn/_180_ ));
 sg13g2_nand2b_1 \u_neuron.u_syn/_563_  (.Y(\u_neuron.u_syn/_187_ ),
    .B(\u_neuron.u_syn/_186_ ),
    .A_N(\u_neuron.u_syn/_182_ ));
 sg13g2_nor4_1 \u_neuron.u_syn/_564_  (.A(net367),
    .B(\u_neuron.u_syn/_046_ ),
    .C(\u_neuron.ltd_idx[0] ),
    .D(\u_neuron.u_syn/_049_ ),
    .Y(\u_neuron.u_syn/_188_ ));
 sg13g2_a21oi_1 \u_neuron.u_syn/_565_  (.A1(net319),
    .A2(\u_neuron.u_syn/_188_ ),
    .Y(\u_neuron.u_syn/_189_ ),
    .B1(net410));
 sg13g2_a22oi_1 \u_neuron.u_syn/_566_  (.Y(\u_neuron.u_syn/_004_ ),
    .B1(\u_neuron.u_syn/_187_ ),
    .B2(\u_neuron.u_syn/_189_ ),
    .A2(\u_neuron.u_syn/_056_ ),
    .A1(net411));
 sg13g2_nor4_1 \u_neuron.u_syn/_567_  (.A(net406),
    .B(\u_neuron.u_syn/_038_ ),
    .C(net409),
    .D(\u_neuron.u_syn/_051_ ),
    .Y(\u_neuron.u_syn/_190_ ));
 sg13g2_a221oi_1 \u_neuron.u_syn/_568_  (.B2(\u_neuron.u_syn/_146_ ),
    .C1(\u_neuron.u_syn/_180_ ),
    .B1(\u_neuron.u_syn/_190_ ),
    .A1(net202),
    .Y(\u_neuron.u_syn/_191_ ),
    .A2(\u_neuron.u_syn/_177_ ));
 sg13g2_nand2_2 \u_neuron.u_syn/_569_  (.Y(\u_neuron.u_syn/_192_ ),
    .A(net333),
    .B(\u_neuron.u_syn/_134_ ));
 sg13g2_a22oi_1 \u_neuron.u_syn/_570_  (.Y(\u_neuron.u_syn/_193_ ),
    .B1(\u_neuron.u_syn/_192_ ),
    .B2(\u_neuron.u_syn/_180_ ),
    .A2(\u_neuron.u_syn/_185_ ),
    .A1(net319));
 sg13g2_nand2b_1 \u_neuron.u_syn/_571_  (.Y(\u_neuron.u_syn/_194_ ),
    .B(\u_neuron.u_syn/_193_ ),
    .A_N(\u_neuron.u_syn/_191_ ));
 sg13g2_nor4_1 \u_neuron.u_syn/_572_  (.A(net367),
    .B(\u_neuron.u_syn/_046_ ),
    .C(\u_neuron.ltd_idx[0] ),
    .D(\u_neuron.u_syn/_053_ ),
    .Y(\u_neuron.u_syn/_195_ ));
 sg13g2_a21oi_1 \u_neuron.u_syn/_573_  (.A1(net319),
    .A2(\u_neuron.u_syn/_195_ ),
    .Y(\u_neuron.u_syn/_196_ ),
    .B1(net411));
 sg13g2_a22oi_1 \u_neuron.u_syn/_574_  (.Y(\u_neuron.u_syn/_005_ ),
    .B1(\u_neuron.u_syn/_194_ ),
    .B2(\u_neuron.u_syn/_196_ ),
    .A2(\u_neuron.u_syn/_057_ ),
    .A1(net411));
 sg13g2_and2_1 \u_neuron.u_syn/_575_  (.A(net408),
    .B(net409),
    .X(\u_neuron.u_syn/_197_ ));
 sg13g2_nor2b_2 \u_neuron.u_syn/_576_  (.A(net404),
    .B_N(\u_neuron.u_syn/_197_ ),
    .Y(\u_neuron.u_syn/_198_ ));
 sg13g2_nand3_1 \u_neuron.u_syn/_577_  (.B(\u_neuron.u_syn/_144_ ),
    .C(\u_neuron.u_syn/_198_ ),
    .A(net359),
    .Y(\u_neuron.u_syn/_199_ ));
 sg13g2_nand2b_1 \u_neuron.u_syn/_578_  (.Y(\u_neuron.u_syn/_200_ ),
    .B(\u_neuron.u_syn/_041_ ),
    .A_N(\u_neuron.u_syn/_199_ ));
 sg13g2_nand2_2 \u_neuron.u_syn/_579_  (.Y(\u_neuron.u_syn/_201_ ),
    .A(\u_neuron.ltp_idx[1] ),
    .B(\u_neuron.ltp_idx[0] ));
 sg13g2_nor2_1 \u_neuron.u_syn/_580_  (.A(\u_neuron.ltp_idx[2] ),
    .B(\u_neuron.u_syn/_201_ ),
    .Y(\u_neuron.u_syn/_202_ ));
 sg13g2_nand3_1 \u_neuron.u_syn/_581_  (.B(\u_neuron.u_syn/_151_ ),
    .C(\u_neuron.u_syn/_202_ ),
    .A(net321),
    .Y(\u_neuron.u_syn/_203_ ));
 sg13g2_a22oi_1 \u_neuron.u_syn/_582_  (.Y(\u_neuron.u_syn/_204_ ),
    .B1(\u_neuron.u_syn/_202_ ),
    .B2(\u_neuron.u_syn/_152_ ),
    .A2(\u_neuron.u_syn/_199_ ),
    .A1(\u_neuron.u_syn/_058_ ));
 sg13g2_nor3_2 \u_neuron.u_syn/_583_  (.A(net367),
    .B(\u_neuron.u_syn/_046_ ),
    .C(\u_neuron.u_syn/_047_ ),
    .Y(\u_neuron.u_syn/_205_ ));
 sg13g2_nand2_1 \u_neuron.u_syn/_584_  (.Y(\u_neuron.u_syn/_206_ ),
    .A(net320),
    .B(\u_neuron.u_syn/_205_ ));
 sg13g2_nor2_1 \u_neuron.u_syn/_585_  (.A(\u_neuron.u_syn/_044_ ),
    .B(\u_neuron.u_syn/_203_ ),
    .Y(\u_neuron.u_syn/_207_ ));
 sg13g2_a221oi_1 \u_neuron.u_syn/_586_  (.B2(net320),
    .C1(\u_neuron.u_syn/_207_ ),
    .B1(\u_neuron.u_syn/_205_ ),
    .A1(\u_neuron.u_syn/_200_ ),
    .Y(\u_neuron.u_syn/_208_ ),
    .A2(\u_neuron.u_syn/_204_ ));
 sg13g2_o21ai_1 \u_neuron.u_syn/_587_  (.B1(net468),
    .Y(\u_neuron.u_syn/_209_ ),
    .A1(net332),
    .A2(\u_neuron.u_syn/_206_ ));
 sg13g2_nand2_1 \u_neuron.u_syn/_588_  (.Y(\u_neuron.u_syn/_210_ ),
    .A(net415),
    .B(net190));
 sg13g2_o21ai_1 \u_neuron.u_syn/_589_  (.B1(\u_neuron.u_syn/_210_ ),
    .Y(\u_neuron.u_syn/_006_ ),
    .A1(\u_neuron.u_syn/_208_ ),
    .A2(\u_neuron.u_syn/_209_ ));
 sg13g2_mux2_1 \u_neuron.u_syn/_590_  (.A0(\u_neuron.cfg_arg[1] ),
    .A1(\u_neuron.wtab[7] ),
    .S(\u_neuron.u_syn/_199_ ),
    .X(\u_neuron.u_syn/_211_ ));
 sg13g2_nor2_1 \u_neuron.u_syn/_591_  (.A(\u_neuron.u_syn/_052_ ),
    .B(\u_neuron.u_syn/_203_ ),
    .Y(\u_neuron.u_syn/_212_ ));
 sg13g2_a221oi_1 \u_neuron.u_syn/_592_  (.B2(\u_neuron.u_syn/_203_ ),
    .C1(\u_neuron.u_syn/_212_ ),
    .B1(\u_neuron.u_syn/_211_ ),
    .A1(net320),
    .Y(\u_neuron.u_syn/_213_ ),
    .A2(\u_neuron.u_syn/_205_ ));
 sg13g2_o21ai_1 \u_neuron.u_syn/_593_  (.B1(net468),
    .Y(\u_neuron.u_syn/_214_ ),
    .A1(net331),
    .A2(\u_neuron.u_syn/_206_ ));
 sg13g2_nand2_1 \u_neuron.u_syn/_594_  (.Y(\u_neuron.u_syn/_215_ ),
    .A(net416),
    .B(net203));
 sg13g2_o21ai_1 \u_neuron.u_syn/_595_  (.B1(\u_neuron.u_syn/_215_ ),
    .Y(\u_neuron.u_syn/_007_ ),
    .A1(\u_neuron.u_syn/_213_ ),
    .A2(\u_neuron.u_syn/_214_ ));
 sg13g2_xor2_1 \u_neuron.u_syn/_596_  (.B(\u_neuron.u_syn/_129_ ),
    .A(net407),
    .X(\u_neuron.u_syn/_216_ ));
 sg13g2_nor4_1 \u_neuron.u_syn/_597_  (.A(\u_neuron.pending_widx[1] ),
    .B(\u_neuron.pending_widx[0] ),
    .C(\u_neuron.u_syn/_041_ ),
    .D(\u_neuron.u_syn/_131_ ),
    .Y(\u_neuron.u_syn/_217_ ));
 sg13g2_nand2b_1 \u_neuron.u_syn/_598_  (.Y(\u_neuron.u_syn/_218_ ),
    .B(\u_neuron.u_syn/_217_ ),
    .A_N(\u_neuron.u_syn/_216_ ));
 sg13g2_nand4_1 \u_neuron.u_syn/_599_  (.B(net407),
    .C(net359),
    .A(\u_neuron.u_syn/_037_ ),
    .Y(\u_neuron.u_syn/_219_ ),
    .D(\u_neuron.u_syn/_129_ ));
 sg13g2_nand2_1 \u_neuron.u_syn/_600_  (.Y(\u_neuron.u_syn/_220_ ),
    .A(net163),
    .B(\u_neuron.u_syn/_219_ ));
 sg13g2_o21ai_1 \u_neuron.u_syn/_601_  (.B1(\u_neuron.u_syn/_220_ ),
    .Y(\u_neuron.u_syn/_221_ ),
    .A1(\u_neuron.u_syn/_147_ ),
    .A2(\u_neuron.u_syn/_218_ ));
 sg13g2_nor3_2 \u_neuron.u_syn/_602_  (.A(\u_neuron.u_syn/_043_ ),
    .B(\u_neuron.ltp_idx[1] ),
    .C(\u_neuron.ltp_idx[0] ),
    .Y(\u_neuron.u_syn/_222_ ));
 sg13g2_nand2_1 \u_neuron.u_syn/_603_  (.Y(\u_neuron.u_syn/_223_ ),
    .A(\u_neuron.u_syn/_152_ ),
    .B(\u_neuron.u_syn/_222_ ));
 sg13g2_nand3_1 \u_neuron.u_syn/_604_  (.B(\u_neuron.u_syn/_046_ ),
    .C(\u_neuron.u_syn/_047_ ),
    .A(net367),
    .Y(\u_neuron.u_syn/_224_ ));
 sg13g2_nor2_1 \u_neuron.u_syn/_605_  (.A(\u_neuron.u_syn/_161_ ),
    .B(\u_neuron.u_syn/_224_ ),
    .Y(\u_neuron.u_syn/_225_ ));
 sg13g2_or2_1 \u_neuron.u_syn/_606_  (.X(\u_neuron.u_syn/_226_ ),
    .B(\u_neuron.u_syn/_224_ ),
    .A(\u_neuron.u_syn/_161_ ));
 sg13g2_and2_1 \u_neuron.u_syn/_607_  (.A(\u_neuron.ltp_wdata[0] ),
    .B(\u_neuron.u_syn/_222_ ),
    .X(\u_neuron.u_syn/_227_ ));
 sg13g2_a221oi_1 \u_neuron.u_syn/_608_  (.B2(\u_neuron.u_syn/_152_ ),
    .C1(\u_neuron.u_syn/_225_ ),
    .B1(\u_neuron.u_syn/_227_ ),
    .A1(\u_neuron.u_syn/_221_ ),
    .Y(\u_neuron.u_syn/_228_ ),
    .A2(\u_neuron.u_syn/_223_ ));
 sg13g2_o21ai_1 \u_neuron.u_syn/_609_  (.B1(net467),
    .Y(\u_neuron.u_syn/_229_ ),
    .A1(net332),
    .A2(\u_neuron.u_syn/_226_ ));
 sg13g2_nand2_1 \u_neuron.u_syn/_610_  (.Y(\u_neuron.u_syn/_230_ ),
    .A(net415),
    .B(net163));
 sg13g2_o21ai_1 \u_neuron.u_syn/_611_  (.B1(\u_neuron.u_syn/_230_ ),
    .Y(\u_neuron.u_syn/_008_ ),
    .A1(\u_neuron.u_syn/_228_ ),
    .A2(\u_neuron.u_syn/_229_ ));
 sg13g2_nor4_1 \u_neuron.u_syn/_612_  (.A(\u_neuron.pending_widx[1] ),
    .B(net238),
    .C(\u_neuron.u_syn/_051_ ),
    .D(\u_neuron.u_syn/_131_ ),
    .Y(\u_neuron.u_syn/_231_ ));
 sg13g2_nand2b_1 \u_neuron.u_syn/_613_  (.Y(\u_neuron.u_syn/_232_ ),
    .B(\u_neuron.u_syn/_231_ ),
    .A_N(\u_neuron.u_syn/_216_ ));
 sg13g2_nand2_1 \u_neuron.u_syn/_614_  (.Y(\u_neuron.u_syn/_233_ ),
    .A(net128),
    .B(\u_neuron.u_syn/_219_ ));
 sg13g2_o21ai_1 \u_neuron.u_syn/_615_  (.B1(\u_neuron.u_syn/_233_ ),
    .Y(\u_neuron.u_syn/_234_ ),
    .A1(\u_neuron.u_syn/_147_ ),
    .A2(\u_neuron.u_syn/_232_ ));
 sg13g2_and2_1 \u_neuron.u_syn/_616_  (.A(net333),
    .B(\u_neuron.u_syn/_222_ ),
    .X(\u_neuron.u_syn/_235_ ));
 sg13g2_a221oi_1 \u_neuron.u_syn/_617_  (.B2(\u_neuron.u_syn/_152_ ),
    .C1(\u_neuron.u_syn/_225_ ),
    .B1(\u_neuron.u_syn/_235_ ),
    .A1(\u_neuron.u_syn/_223_ ),
    .Y(\u_neuron.u_syn/_236_ ),
    .A2(\u_neuron.u_syn/_234_ ));
 sg13g2_o21ai_1 \u_neuron.u_syn/_618_  (.B1(net467),
    .Y(\u_neuron.u_syn/_237_ ),
    .A1(net331),
    .A2(\u_neuron.u_syn/_226_ ));
 sg13g2_nand2_1 \u_neuron.u_syn/_619_  (.Y(\u_neuron.u_syn/_238_ ),
    .A(net415),
    .B(net128));
 sg13g2_o21ai_1 \u_neuron.u_syn/_620_  (.B1(\u_neuron.u_syn/_238_ ),
    .Y(\u_neuron.u_syn/_009_ ),
    .A1(\u_neuron.u_syn/_236_ ),
    .A2(\u_neuron.u_syn/_237_ ));
 sg13g2_and2_1 \u_neuron.u_syn/_621_  (.A(net407),
    .B(\u_neuron.u_syn/_148_ ),
    .X(\u_neuron.u_syn/_239_ ));
 sg13g2_nand4_1 \u_neuron.u_syn/_622_  (.B(net407),
    .C(net360),
    .A(\u_neuron.u_syn/_037_ ),
    .Y(\u_neuron.u_syn/_240_ ),
    .D(\u_neuron.u_syn/_148_ ));
 sg13g2_nand2_1 \u_neuron.u_syn/_623_  (.Y(\u_neuron.u_syn/_241_ ),
    .A(net179),
    .B(\u_neuron.u_syn/_240_ ));
 sg13g2_nand4_1 \u_neuron.u_syn/_624_  (.B(\u_neuron.ltp_idx[2] ),
    .C(net321),
    .A(\u_neuron.u_syn/_042_ ),
    .Y(\u_neuron.u_syn/_242_ ),
    .D(\u_neuron.u_syn/_153_ ));
 sg13g2_nand4_1 \u_neuron.u_syn/_625_  (.B(net360),
    .C(\u_neuron.u_syn/_144_ ),
    .A(\u_neuron.cfg_arg[0] ),
    .Y(\u_neuron.u_syn/_243_ ),
    .D(\u_neuron.u_syn/_239_ ));
 sg13g2_nand3_1 \u_neuron.u_syn/_626_  (.B(\u_neuron.u_syn/_242_ ),
    .C(\u_neuron.u_syn/_243_ ),
    .A(\u_neuron.u_syn/_241_ ),
    .Y(\u_neuron.u_syn/_244_ ));
 sg13g2_nor2_1 \u_neuron.u_syn/_627_  (.A(\u_neuron.ltp_wdata[0] ),
    .B(\u_neuron.u_syn/_242_ ),
    .Y(\u_neuron.u_syn/_245_ ));
 sg13g2_and2_1 \u_neuron.u_syn/_628_  (.A(net368),
    .B(\u_neuron.u_syn/_162_ ),
    .X(\u_neuron.u_syn/_246_ ));
 sg13g2_a21oi_1 \u_neuron.u_syn/_629_  (.A1(\u_neuron.u_syn/_160_ ),
    .A2(\u_neuron.u_syn/_246_ ),
    .Y(\u_neuron.u_syn/_247_ ),
    .B1(\u_neuron.u_syn/_245_ ));
 sg13g2_nand2_1 \u_neuron.u_syn/_630_  (.Y(\u_neuron.u_syn/_248_ ),
    .A(\u_neuron.ltd_wdata[0] ),
    .B(\u_neuron.u_syn/_246_ ));
 sg13g2_o21ai_1 \u_neuron.u_syn/_631_  (.B1(net467),
    .Y(\u_neuron.u_syn/_249_ ),
    .A1(\u_neuron.u_syn/_161_ ),
    .A2(\u_neuron.u_syn/_248_ ));
 sg13g2_a21oi_1 \u_neuron.u_syn/_632_  (.A1(\u_neuron.u_syn/_244_ ),
    .A2(\u_neuron.u_syn/_247_ ),
    .Y(\u_neuron.u_syn/_250_ ),
    .B1(\u_neuron.u_syn/_249_ ));
 sg13g2_a21oi_1 \u_neuron.u_syn/_633_  (.A1(net416),
    .A2(\u_neuron.u_syn/_059_ ),
    .Y(\u_neuron.u_syn/_010_ ),
    .B1(\u_neuron.u_syn/_250_ ));
 sg13g2_o21ai_1 \u_neuron.u_syn/_634_  (.B1(\u_neuron.u_syn/_242_ ),
    .Y(\u_neuron.u_syn/_251_ ),
    .A1(\u_neuron.u_syn/_051_ ),
    .A2(\u_neuron.u_syn/_240_ ));
 sg13g2_a21o_1 \u_neuron.u_syn/_635_  (.A2(\u_neuron.u_syn/_240_ ),
    .A1(net184),
    .B1(\u_neuron.u_syn/_251_ ),
    .X(\u_neuron.u_syn/_252_ ));
 sg13g2_nor2_1 \u_neuron.u_syn/_636_  (.A(net333),
    .B(\u_neuron.u_syn/_242_ ),
    .Y(\u_neuron.u_syn/_253_ ));
 sg13g2_a21oi_1 \u_neuron.u_syn/_637_  (.A1(\u_neuron.u_syn/_160_ ),
    .A2(\u_neuron.u_syn/_246_ ),
    .Y(\u_neuron.u_syn/_254_ ),
    .B1(\u_neuron.u_syn/_253_ ));
 sg13g2_nand2_1 \u_neuron.u_syn/_638_  (.Y(\u_neuron.u_syn/_255_ ),
    .A(\u_neuron.ltd_wdata[1] ),
    .B(\u_neuron.u_syn/_246_ ));
 sg13g2_o21ai_1 \u_neuron.u_syn/_639_  (.B1(net467),
    .Y(\u_neuron.u_syn/_256_ ),
    .A1(\u_neuron.u_syn/_161_ ),
    .A2(\u_neuron.u_syn/_255_ ));
 sg13g2_a21oi_1 \u_neuron.u_syn/_640_  (.A1(\u_neuron.u_syn/_252_ ),
    .A2(\u_neuron.u_syn/_254_ ),
    .Y(\u_neuron.u_syn/_257_ ),
    .B1(\u_neuron.u_syn/_256_ ));
 sg13g2_a21oi_1 \u_neuron.u_syn/_641_  (.A1(net415),
    .A2(\u_neuron.u_syn/_060_ ),
    .Y(\u_neuron.u_syn/_011_ ),
    .B1(\u_neuron.u_syn/_257_ ));
 sg13g2_nand4_1 \u_neuron.u_syn/_642_  (.B(net404),
    .C(net358),
    .A(\u_neuron.u_syn/_037_ ),
    .Y(\u_neuron.u_syn/_258_ ),
    .D(\u_neuron.u_syn/_175_ ));
 sg13g2_nand2_1 \u_neuron.u_syn/_643_  (.Y(\u_neuron.u_syn/_259_ ),
    .A(net207),
    .B(\u_neuron.u_syn/_258_ ));
 sg13g2_nor4_2 \u_neuron.u_syn/_644_  (.A(\u_neuron.ltp_idx[3] ),
    .B(\u_neuron.u_syn/_043_ ),
    .C(net315),
    .Y(\u_neuron.u_syn/_260_ ),
    .D(\u_neuron.u_syn/_178_ ));
 sg13g2_nand4_1 \u_neuron.u_syn/_645_  (.B(net408),
    .C(\u_neuron.u_syn/_039_ ),
    .A(net404),
    .Y(\u_neuron.u_syn/_261_ ),
    .D(\u_neuron.cfg_arg[0] ));
 sg13g2_o21ai_1 \u_neuron.u_syn/_646_  (.B1(\u_neuron.u_syn/_259_ ),
    .Y(\u_neuron.u_syn/_262_ ),
    .A1(\u_neuron.u_syn/_147_ ),
    .A2(\u_neuron.u_syn/_261_ ));
 sg13g2_and2_1 \u_neuron.u_syn/_647_  (.A(net367),
    .B(\u_neuron.u_syn/_184_ ),
    .X(\u_neuron.u_syn/_263_ ));
 sg13g2_a22oi_1 \u_neuron.u_syn/_648_  (.Y(\u_neuron.u_syn/_264_ ),
    .B1(\u_neuron.u_syn/_263_ ),
    .B2(net319),
    .A2(\u_neuron.u_syn/_260_ ),
    .A1(\u_neuron.u_syn/_183_ ));
 sg13g2_o21ai_1 \u_neuron.u_syn/_649_  (.B1(\u_neuron.u_syn/_264_ ),
    .Y(\u_neuron.u_syn/_265_ ),
    .A1(\u_neuron.u_syn/_260_ ),
    .A2(\u_neuron.u_syn/_262_ ));
 sg13g2_and3_1 \u_neuron.u_syn/_650_  (.X(\u_neuron.u_syn/_266_ ),
    .A(net368),
    .B(net332),
    .C(\u_neuron.u_syn/_184_ ));
 sg13g2_a21oi_1 \u_neuron.u_syn/_651_  (.A1(net320),
    .A2(\u_neuron.u_syn/_266_ ),
    .Y(\u_neuron.u_syn/_267_ ),
    .B1(net413));
 sg13g2_a22oi_1 \u_neuron.u_syn/_652_  (.Y(\u_neuron.u_syn/_012_ ),
    .B1(\u_neuron.u_syn/_265_ ),
    .B2(\u_neuron.u_syn/_267_ ),
    .A2(\u_neuron.u_syn/_061_ ),
    .A1(net413));
 sg13g2_nand2_1 \u_neuron.u_syn/_653_  (.Y(\u_neuron.u_syn/_268_ ),
    .A(net172),
    .B(\u_neuron.u_syn/_258_ ));
 sg13g2_nand4_1 \u_neuron.u_syn/_654_  (.B(net408),
    .C(\u_neuron.u_syn/_039_ ),
    .A(net404),
    .Y(\u_neuron.u_syn/_269_ ),
    .D(\u_neuron.cfg_arg[1] ));
 sg13g2_o21ai_1 \u_neuron.u_syn/_655_  (.B1(\u_neuron.u_syn/_268_ ),
    .Y(\u_neuron.u_syn/_270_ ),
    .A1(\u_neuron.u_syn/_147_ ),
    .A2(\u_neuron.u_syn/_269_ ));
 sg13g2_a22oi_1 \u_neuron.u_syn/_656_  (.Y(\u_neuron.u_syn/_271_ ),
    .B1(\u_neuron.u_syn/_263_ ),
    .B2(net320),
    .A2(\u_neuron.u_syn/_260_ ),
    .A1(\u_neuron.u_syn/_192_ ));
 sg13g2_o21ai_1 \u_neuron.u_syn/_657_  (.B1(\u_neuron.u_syn/_271_ ),
    .Y(\u_neuron.u_syn/_272_ ),
    .A1(\u_neuron.u_syn/_260_ ),
    .A2(\u_neuron.u_syn/_270_ ));
 sg13g2_and3_1 \u_neuron.u_syn/_658_  (.X(\u_neuron.u_syn/_273_ ),
    .A(net368),
    .B(net331),
    .C(\u_neuron.u_syn/_184_ ));
 sg13g2_a21oi_1 \u_neuron.u_syn/_659_  (.A1(net320),
    .A2(\u_neuron.u_syn/_273_ ),
    .Y(\u_neuron.u_syn/_274_ ),
    .B1(net413));
 sg13g2_a22oi_1 \u_neuron.u_syn/_660_  (.Y(\u_neuron.u_syn/_013_ ),
    .B1(\u_neuron.u_syn/_272_ ),
    .B2(\u_neuron.u_syn/_274_ ),
    .A2(\u_neuron.u_syn/_062_ ),
    .A1(net413));
 sg13g2_nand4_1 \u_neuron.u_syn/_661_  (.B(net404),
    .C(net358),
    .A(\u_neuron.u_syn/_037_ ),
    .Y(\u_neuron.u_syn/_275_ ),
    .D(\u_neuron.u_syn/_197_ ));
 sg13g2_nor4_1 \u_neuron.u_syn/_662_  (.A(\u_neuron.ltp_idx[3] ),
    .B(\u_neuron.u_syn/_043_ ),
    .C(net315),
    .D(\u_neuron.u_syn/_201_ ),
    .Y(\u_neuron.u_syn/_276_ ));
 sg13g2_or4_1 \u_neuron.u_syn/_663_  (.A(\u_neuron.ltp_idx[3] ),
    .B(\u_neuron.u_syn/_043_ ),
    .C(net315),
    .D(\u_neuron.u_syn/_201_ ),
    .X(\u_neuron.u_syn/_277_ ));
 sg13g2_nand3_1 \u_neuron.u_syn/_664_  (.B(\u_neuron.cfg_arg[0] ),
    .C(\u_neuron.u_syn/_197_ ),
    .A(net404),
    .Y(\u_neuron.u_syn/_278_ ));
 sg13g2_a21oi_1 \u_neuron.u_syn/_665_  (.A1(net186),
    .A2(\u_neuron.u_syn/_275_ ),
    .Y(\u_neuron.u_syn/_279_ ),
    .B1(\u_neuron.u_syn/_276_ ));
 sg13g2_o21ai_1 \u_neuron.u_syn/_666_  (.B1(\u_neuron.u_syn/_279_ ),
    .Y(\u_neuron.u_syn/_280_ ),
    .A1(\u_neuron.u_syn/_147_ ),
    .A2(\u_neuron.u_syn/_278_ ));
 sg13g2_and3_2 \u_neuron.u_syn/_667_  (.X(\u_neuron.u_syn/_281_ ),
    .A(net368),
    .B(\u_neuron.ltd_idx[1] ),
    .C(\u_neuron.ltd_idx[0] ));
 sg13g2_nand2_1 \u_neuron.u_syn/_668_  (.Y(\u_neuron.u_syn/_282_ ),
    .A(net319),
    .B(\u_neuron.u_syn/_281_ ));
 sg13g2_nand2_1 \u_neuron.u_syn/_669_  (.Y(\u_neuron.u_syn/_283_ ),
    .A(\u_neuron.u_syn/_044_ ),
    .B(\u_neuron.u_syn/_276_ ));
 sg13g2_nand3_1 \u_neuron.u_syn/_670_  (.B(\u_neuron.u_syn/_282_ ),
    .C(\u_neuron.u_syn/_283_ ),
    .A(\u_neuron.u_syn/_280_ ),
    .Y(\u_neuron.u_syn/_284_ ));
 sg13g2_and2_1 \u_neuron.u_syn/_671_  (.A(net332),
    .B(\u_neuron.u_syn/_281_ ),
    .X(\u_neuron.u_syn/_285_ ));
 sg13g2_a21oi_1 \u_neuron.u_syn/_672_  (.A1(net319),
    .A2(\u_neuron.u_syn/_285_ ),
    .Y(\u_neuron.u_syn/_286_ ),
    .B1(net412));
 sg13g2_a22oi_1 \u_neuron.u_syn/_673_  (.Y(\u_neuron.u_syn/_014_ ),
    .B1(\u_neuron.u_syn/_284_ ),
    .B2(\u_neuron.u_syn/_286_ ),
    .A2(\u_neuron.u_syn/_063_ ),
    .A1(net413));
 sg13g2_o21ai_1 \u_neuron.u_syn/_674_  (.B1(\u_neuron.u_syn/_277_ ),
    .Y(\u_neuron.u_syn/_287_ ),
    .A1(\u_neuron.cfg_arg[1] ),
    .A2(\u_neuron.u_syn/_275_ ));
 sg13g2_a21oi_1 \u_neuron.u_syn/_675_  (.A1(\u_neuron.u_syn/_064_ ),
    .A2(\u_neuron.u_syn/_275_ ),
    .Y(\u_neuron.u_syn/_288_ ),
    .B1(\u_neuron.u_syn/_287_ ));
 sg13g2_a221oi_1 \u_neuron.u_syn/_676_  (.B2(net319),
    .C1(\u_neuron.u_syn/_288_ ),
    .B1(\u_neuron.u_syn/_281_ ),
    .A1(net333),
    .Y(\u_neuron.u_syn/_289_ ),
    .A2(\u_neuron.u_syn/_276_ ));
 sg13g2_o21ai_1 \u_neuron.u_syn/_677_  (.B1(net465),
    .Y(\u_neuron.u_syn/_290_ ),
    .A1(net331),
    .A2(\u_neuron.u_syn/_282_ ));
 sg13g2_nand2_1 \u_neuron.u_syn/_678_  (.Y(\u_neuron.u_syn/_291_ ),
    .A(net413),
    .B(net111));
 sg13g2_o21ai_1 \u_neuron.u_syn/_679_  (.B1(\u_neuron.u_syn/_291_ ),
    .Y(\u_neuron.u_syn/_015_ ),
    .A1(\u_neuron.u_syn/_289_ ),
    .A2(\u_neuron.u_syn/_290_ ));
 sg13g2_nor2_1 \u_neuron.u_syn/_680_  (.A(net465),
    .B(net174),
    .Y(\u_neuron.u_syn/_292_ ));
 sg13g2_nand3_1 \u_neuron.u_syn/_681_  (.B(\u_neuron.u_syn/_216_ ),
    .C(\u_neuron.u_syn/_217_ ),
    .A(net359),
    .Y(\u_neuron.u_syn/_293_ ));
 sg13g2_and3_2 \u_neuron.u_syn/_682_  (.X(\u_neuron.u_syn/_294_ ),
    .A(\u_neuron.ltp_idx[3] ),
    .B(net321),
    .C(\u_neuron.u_syn/_133_ ));
 sg13g2_nand3_1 \u_neuron.u_syn/_683_  (.B(net358),
    .C(\u_neuron.u_syn/_130_ ),
    .A(\u_neuron.pending_widx[3] ),
    .Y(\u_neuron.u_syn/_295_ ));
 sg13g2_a21oi_1 \u_neuron.u_syn/_684_  (.A1(net174),
    .A2(\u_neuron.u_syn/_295_ ),
    .Y(\u_neuron.u_syn/_296_ ),
    .B1(\u_neuron.u_syn/_294_ ));
 sg13g2_nand2_1 \u_neuron.u_syn/_685_  (.Y(\u_neuron.u_syn/_297_ ),
    .A(\u_neuron.u_syn/_293_ ),
    .B(\u_neuron.u_syn/_296_ ));
 sg13g2_and3_2 \u_neuron.u_syn/_686_  (.X(\u_neuron.u_syn/_298_ ),
    .A(\u_neuron.ltd_idx[3] ),
    .B(\u_neuron.ltd_we ),
    .C(\u_neuron.u_syn/_127_ ));
 sg13g2_a21oi_1 \u_neuron.u_syn/_687_  (.A1(\u_neuron.u_syn/_044_ ),
    .A2(\u_neuron.u_syn/_294_ ),
    .Y(\u_neuron.u_syn/_299_ ),
    .B1(\u_neuron.u_syn/_298_ ));
 sg13g2_a22oi_1 \u_neuron.u_syn/_688_  (.Y(\u_neuron.u_syn/_300_ ),
    .B1(\u_neuron.u_syn/_299_ ),
    .B2(\u_neuron.u_syn/_297_ ),
    .A2(\u_neuron.u_syn/_298_ ),
    .A1(net332));
 sg13g2_a21oi_1 \u_neuron.u_syn/_689_  (.A1(net465),
    .A2(\u_neuron.u_syn/_300_ ),
    .Y(\u_neuron.u_syn/_016_ ),
    .B1(\u_neuron.u_syn/_292_ ));
 sg13g2_nand3_1 \u_neuron.u_syn/_690_  (.B(\u_neuron.u_syn/_216_ ),
    .C(\u_neuron.u_syn/_231_ ),
    .A(net359),
    .Y(\u_neuron.u_syn/_301_ ));
 sg13g2_a21oi_1 \u_neuron.u_syn/_691_  (.A1(net205),
    .A2(\u_neuron.u_syn/_295_ ),
    .Y(\u_neuron.u_syn/_302_ ),
    .B1(\u_neuron.u_syn/_294_ ));
 sg13g2_a221oi_1 \u_neuron.u_syn/_692_  (.B2(\u_neuron.u_syn/_302_ ),
    .C1(\u_neuron.u_syn/_298_ ),
    .B1(\u_neuron.u_syn/_301_ ),
    .A1(\u_neuron.u_syn/_052_ ),
    .Y(\u_neuron.u_syn/_303_ ),
    .A2(\u_neuron.u_syn/_294_ ));
 sg13g2_nand2_1 \u_neuron.u_syn/_693_  (.Y(\u_neuron.u_syn/_304_ ),
    .A(net331),
    .B(\u_neuron.u_syn/_298_ ));
 sg13g2_nor2_1 \u_neuron.u_syn/_694_  (.A(net411),
    .B(\u_neuron.u_syn/_303_ ),
    .Y(\u_neuron.u_syn/_305_ ));
 sg13g2_a22oi_1 \u_neuron.u_syn/_695_  (.Y(\u_neuron.u_syn/_017_ ),
    .B1(\u_neuron.u_syn/_304_ ),
    .B2(\u_neuron.u_syn/_305_ ),
    .A2(\u_neuron.u_syn/_065_ ),
    .A1(net414));
 sg13g2_and2_1 \u_neuron.u_syn/_696_  (.A(net357),
    .B(\u_neuron.u_syn/_145_ ),
    .X(\u_neuron.u_syn/_306_ ));
 sg13g2_nand2_2 \u_neuron.u_syn/_697_  (.Y(\u_neuron.u_syn/_307_ ),
    .A(net358),
    .B(\u_neuron.u_syn/_145_ ));
 sg13g2_nand3_1 \u_neuron.u_syn/_698_  (.B(\u_neuron.u_syn/_145_ ),
    .C(\u_neuron.u_syn/_149_ ),
    .A(net358),
    .Y(\u_neuron.u_syn/_308_ ));
 sg13g2_nor2_1 \u_neuron.u_syn/_699_  (.A(\u_neuron.u_syn/_045_ ),
    .B(\u_neuron.u_syn/_151_ ),
    .Y(\u_neuron.u_syn/_309_ ));
 sg13g2_nor3_2 \u_neuron.u_syn/_700_  (.A(net315),
    .B(\u_neuron.u_syn/_151_ ),
    .C(\u_neuron.u_syn/_155_ ),
    .Y(\u_neuron.u_syn/_310_ ));
 sg13g2_a221oi_1 \u_neuron.u_syn/_701_  (.B2(net204),
    .C1(\u_neuron.u_syn/_310_ ),
    .B1(\u_neuron.u_syn/_308_ ),
    .A1(\u_neuron.u_syn/_157_ ),
    .Y(\u_neuron.u_syn/_311_ ),
    .A2(\u_neuron.u_syn/_306_ ));
 sg13g2_nor2b_1 \u_neuron.u_syn/_702_  (.A(\u_neuron.u_syn/_159_ ),
    .B_N(\u_neuron.ltd_we ),
    .Y(\u_neuron.u_syn/_312_ ));
 sg13g2_nand2b_2 \u_neuron.u_syn/_703_  (.Y(\u_neuron.u_syn/_313_ ),
    .B(\u_neuron.ltd_we ),
    .A_N(\u_neuron.u_syn/_159_ ));
 sg13g2_and2_1 \u_neuron.u_syn/_704_  (.A(\u_neuron.u_syn/_163_ ),
    .B(net316),
    .X(\u_neuron.u_syn/_314_ ));
 sg13g2_a22oi_1 \u_neuron.u_syn/_705_  (.Y(\u_neuron.u_syn/_315_ ),
    .B1(net318),
    .B2(\u_neuron.u_syn/_163_ ),
    .A2(\u_neuron.u_syn/_310_ ),
    .A1(\u_neuron.u_syn/_044_ ));
 sg13g2_nand2b_1 \u_neuron.u_syn/_706_  (.Y(\u_neuron.u_syn/_316_ ),
    .B(\u_neuron.u_syn/_315_ ),
    .A_N(\u_neuron.u_syn/_311_ ));
 sg13g2_a21oi_1 \u_neuron.u_syn/_707_  (.A1(\u_neuron.u_syn/_167_ ),
    .A2(net318),
    .Y(\u_neuron.u_syn/_317_ ),
    .B1(net414));
 sg13g2_a22oi_1 \u_neuron.u_syn/_708_  (.Y(\u_neuron.u_syn/_018_ ),
    .B1(\u_neuron.u_syn/_316_ ),
    .B2(\u_neuron.u_syn/_317_ ),
    .A2(\u_neuron.u_syn/_066_ ),
    .A1(net414));
 sg13g2_nand2b_1 \u_neuron.u_syn/_709_  (.Y(\u_neuron.u_syn/_318_ ),
    .B(\u_neuron.u_syn/_051_ ),
    .A_N(\u_neuron.u_syn/_308_ ));
 sg13g2_a21oi_1 \u_neuron.u_syn/_710_  (.A1(\u_neuron.u_syn/_067_ ),
    .A2(\u_neuron.u_syn/_308_ ),
    .Y(\u_neuron.u_syn/_319_ ),
    .B1(\u_neuron.u_syn/_310_ ));
 sg13g2_a221oi_1 \u_neuron.u_syn/_711_  (.B2(\u_neuron.u_syn/_319_ ),
    .C1(\u_neuron.u_syn/_314_ ),
    .B1(\u_neuron.u_syn/_318_ ),
    .A1(net333),
    .Y(\u_neuron.u_syn/_320_ ),
    .A2(\u_neuron.u_syn/_310_ ));
 sg13g2_a21o_1 \u_neuron.u_syn/_712_  (.A2(\u_neuron.u_syn/_314_ ),
    .A1(\u_neuron.u_syn/_053_ ),
    .B1(net411),
    .X(\u_neuron.u_syn/_321_ ));
 sg13g2_nand2_1 \u_neuron.u_syn/_713_  (.Y(\u_neuron.u_syn/_322_ ),
    .A(net410),
    .B(net129));
 sg13g2_o21ai_1 \u_neuron.u_syn/_714_  (.B1(\u_neuron.u_syn/_322_ ),
    .Y(\u_neuron.u_syn/_019_ ),
    .A1(\u_neuron.u_syn/_320_ ),
    .A2(\u_neuron.u_syn/_321_ ));
 sg13g2_nand3_1 \u_neuron.u_syn/_715_  (.B(\u_neuron.u_syn/_145_ ),
    .C(\u_neuron.u_syn/_176_ ),
    .A(net357),
    .Y(\u_neuron.u_syn/_323_ ));
 sg13g2_nor4_2 \u_neuron.u_syn/_716_  (.A(\u_neuron.ltp_idx[2] ),
    .B(net315),
    .C(\u_neuron.u_syn/_151_ ),
    .Y(\u_neuron.u_syn/_324_ ),
    .D(\u_neuron.u_syn/_178_ ));
 sg13g2_a221oi_1 \u_neuron.u_syn/_717_  (.B2(net185),
    .C1(\u_neuron.u_syn/_324_ ),
    .B1(\u_neuron.u_syn/_323_ ),
    .A1(\u_neuron.u_syn/_181_ ),
    .Y(\u_neuron.u_syn/_325_ ),
    .A2(\u_neuron.u_syn/_306_ ));
 sg13g2_a22oi_1 \u_neuron.u_syn/_718_  (.Y(\u_neuron.u_syn/_326_ ),
    .B1(\u_neuron.u_syn/_324_ ),
    .B2(\u_neuron.u_syn/_183_ ),
    .A2(net316),
    .A1(\u_neuron.u_syn/_185_ ));
 sg13g2_nand2b_1 \u_neuron.u_syn/_719_  (.Y(\u_neuron.u_syn/_327_ ),
    .B(\u_neuron.u_syn/_326_ ),
    .A_N(\u_neuron.u_syn/_325_ ));
 sg13g2_a21oi_1 \u_neuron.u_syn/_720_  (.A1(\u_neuron.u_syn/_188_ ),
    .A2(net316),
    .Y(\u_neuron.u_syn/_328_ ),
    .B1(net410));
 sg13g2_a22oi_1 \u_neuron.u_syn/_721_  (.Y(\u_neuron.u_syn/_020_ ),
    .B1(\u_neuron.u_syn/_327_ ),
    .B2(\u_neuron.u_syn/_328_ ),
    .A2(\u_neuron.u_syn/_068_ ),
    .A1(net410));
 sg13g2_a221oi_1 \u_neuron.u_syn/_722_  (.B2(net208),
    .C1(\u_neuron.u_syn/_324_ ),
    .B1(\u_neuron.u_syn/_323_ ),
    .A1(\u_neuron.u_syn/_190_ ),
    .Y(\u_neuron.u_syn/_329_ ),
    .A2(\u_neuron.u_syn/_306_ ));
 sg13g2_a22oi_1 \u_neuron.u_syn/_723_  (.Y(\u_neuron.u_syn/_330_ ),
    .B1(\u_neuron.u_syn/_324_ ),
    .B2(\u_neuron.u_syn/_192_ ),
    .A2(net316),
    .A1(\u_neuron.u_syn/_185_ ));
 sg13g2_nand2b_1 \u_neuron.u_syn/_724_  (.Y(\u_neuron.u_syn/_331_ ),
    .B(\u_neuron.u_syn/_330_ ),
    .A_N(\u_neuron.u_syn/_329_ ));
 sg13g2_a21oi_1 \u_neuron.u_syn/_725_  (.A1(\u_neuron.u_syn/_195_ ),
    .A2(net316),
    .Y(\u_neuron.u_syn/_332_ ),
    .B1(net410));
 sg13g2_a22oi_1 \u_neuron.u_syn/_726_  (.Y(\u_neuron.u_syn/_021_ ),
    .B1(\u_neuron.u_syn/_331_ ),
    .B2(\u_neuron.u_syn/_332_ ),
    .A2(\u_neuron.u_syn/_069_ ),
    .A1(net410));
 sg13g2_nand3_1 \u_neuron.u_syn/_727_  (.B(\u_neuron.u_syn/_145_ ),
    .C(\u_neuron.u_syn/_198_ ),
    .A(net357),
    .Y(\u_neuron.u_syn/_333_ ));
 sg13g2_nand2b_1 \u_neuron.u_syn/_728_  (.Y(\u_neuron.u_syn/_334_ ),
    .B(\u_neuron.u_syn/_041_ ),
    .A_N(\u_neuron.u_syn/_333_ ));
 sg13g2_nor4_2 \u_neuron.u_syn/_729_  (.A(\u_neuron.ltp_idx[2] ),
    .B(net315),
    .C(\u_neuron.u_syn/_151_ ),
    .Y(\u_neuron.u_syn/_335_ ),
    .D(\u_neuron.u_syn/_201_ ));
 sg13g2_a21oi_1 \u_neuron.u_syn/_730_  (.A1(\u_neuron.u_syn/_070_ ),
    .A2(\u_neuron.u_syn/_333_ ),
    .Y(\u_neuron.u_syn/_336_ ),
    .B1(\u_neuron.u_syn/_335_ ));
 sg13g2_and2_1 \u_neuron.u_syn/_731_  (.A(\u_neuron.u_syn/_205_ ),
    .B(net316),
    .X(\u_neuron.u_syn/_337_ ));
 sg13g2_nand2_1 \u_neuron.u_syn/_732_  (.Y(\u_neuron.u_syn/_338_ ),
    .A(\u_neuron.u_syn/_205_ ),
    .B(net316));
 sg13g2_a221oi_1 \u_neuron.u_syn/_733_  (.B2(\u_neuron.u_syn/_334_ ),
    .C1(\u_neuron.u_syn/_337_ ),
    .B1(\u_neuron.u_syn/_336_ ),
    .A1(\u_neuron.ltp_wdata[0] ),
    .Y(\u_neuron.u_syn/_339_ ),
    .A2(\u_neuron.u_syn/_335_ ));
 sg13g2_o21ai_1 \u_neuron.u_syn/_734_  (.B1(net466),
    .Y(\u_neuron.u_syn/_340_ ),
    .A1(net332),
    .A2(\u_neuron.u_syn/_338_ ));
 sg13g2_nand2_1 \u_neuron.u_syn/_735_  (.Y(\u_neuron.u_syn/_341_ ),
    .A(net410),
    .B(net148));
 sg13g2_o21ai_1 \u_neuron.u_syn/_736_  (.B1(\u_neuron.u_syn/_341_ ),
    .Y(\u_neuron.u_syn/_022_ ),
    .A1(\u_neuron.u_syn/_339_ ),
    .A2(\u_neuron.u_syn/_340_ ));
 sg13g2_nand2_1 \u_neuron.u_syn/_737_  (.Y(\u_neuron.u_syn/_342_ ),
    .A(\u_neuron.u_syn/_071_ ),
    .B(\u_neuron.u_syn/_333_ ));
 sg13g2_nand4_1 \u_neuron.u_syn/_738_  (.B(\u_neuron.u_syn/_051_ ),
    .C(\u_neuron.u_syn/_145_ ),
    .A(net357),
    .Y(\u_neuron.u_syn/_343_ ),
    .D(\u_neuron.u_syn/_198_ ));
 sg13g2_nor2b_1 \u_neuron.u_syn/_739_  (.A(\u_neuron.u_syn/_335_ ),
    .B_N(\u_neuron.u_syn/_343_ ),
    .Y(\u_neuron.u_syn/_344_ ));
 sg13g2_a221oi_1 \u_neuron.u_syn/_740_  (.B2(\u_neuron.u_syn/_344_ ),
    .C1(\u_neuron.u_syn/_337_ ),
    .B1(\u_neuron.u_syn/_342_ ),
    .A1(net333),
    .Y(\u_neuron.u_syn/_345_ ),
    .A2(\u_neuron.u_syn/_335_ ));
 sg13g2_o21ai_1 \u_neuron.u_syn/_741_  (.B1(net466),
    .Y(\u_neuron.u_syn/_346_ ),
    .A1(net331),
    .A2(\u_neuron.u_syn/_338_ ));
 sg13g2_nand2_1 \u_neuron.u_syn/_742_  (.Y(\u_neuron.u_syn/_347_ ),
    .A(net410),
    .B(net147));
 sg13g2_o21ai_1 \u_neuron.u_syn/_743_  (.B1(\u_neuron.u_syn/_347_ ),
    .Y(\u_neuron.u_syn/_023_ ),
    .A1(\u_neuron.u_syn/_345_ ),
    .A2(\u_neuron.u_syn/_346_ ));
 sg13g2_nand4_1 \u_neuron.u_syn/_744_  (.B(net407),
    .C(net359),
    .A(\u_neuron.pending_widx[3] ),
    .Y(\u_neuron.u_syn/_348_ ),
    .D(\u_neuron.u_syn/_129_ ));
 sg13g2_nand2_1 \u_neuron.u_syn/_745_  (.Y(\u_neuron.u_syn/_349_ ),
    .A(net183),
    .B(\u_neuron.u_syn/_348_ ));
 sg13g2_o21ai_1 \u_neuron.u_syn/_746_  (.B1(\u_neuron.u_syn/_349_ ),
    .Y(\u_neuron.u_syn/_350_ ),
    .A1(\u_neuron.u_syn/_218_ ),
    .A2(\u_neuron.u_syn/_307_ ));
 sg13g2_nand2_1 \u_neuron.u_syn/_747_  (.Y(\u_neuron.u_syn/_351_ ),
    .A(\u_neuron.u_syn/_222_ ),
    .B(\u_neuron.u_syn/_309_ ));
 sg13g2_nor2_1 \u_neuron.u_syn/_748_  (.A(\u_neuron.u_syn/_224_ ),
    .B(\u_neuron.u_syn/_313_ ),
    .Y(\u_neuron.u_syn/_352_ ));
 sg13g2_nand2b_1 \u_neuron.u_syn/_749_  (.Y(\u_neuron.u_syn/_353_ ),
    .B(net318),
    .A_N(\u_neuron.u_syn/_224_ ));
 sg13g2_a221oi_1 \u_neuron.u_syn/_750_  (.B2(\u_neuron.u_syn/_351_ ),
    .C1(\u_neuron.u_syn/_352_ ),
    .B1(\u_neuron.u_syn/_350_ ),
    .A1(\u_neuron.u_syn/_227_ ),
    .Y(\u_neuron.u_syn/_354_ ),
    .A2(\u_neuron.u_syn/_309_ ));
 sg13g2_o21ai_1 \u_neuron.u_syn/_751_  (.B1(net467),
    .Y(\u_neuron.u_syn/_355_ ),
    .A1(\u_neuron.ltd_wdata[0] ),
    .A2(\u_neuron.u_syn/_353_ ));
 sg13g2_nand2_1 \u_neuron.u_syn/_752_  (.Y(\u_neuron.u_syn/_356_ ),
    .A(net415),
    .B(net183));
 sg13g2_o21ai_1 \u_neuron.u_syn/_753_  (.B1(\u_neuron.u_syn/_356_ ),
    .Y(\u_neuron.u_syn/_024_ ),
    .A1(\u_neuron.u_syn/_354_ ),
    .A2(\u_neuron.u_syn/_355_ ));
 sg13g2_nand2_1 \u_neuron.u_syn/_754_  (.Y(\u_neuron.u_syn/_357_ ),
    .A(net193),
    .B(\u_neuron.u_syn/_348_ ));
 sg13g2_o21ai_1 \u_neuron.u_syn/_755_  (.B1(\u_neuron.u_syn/_357_ ),
    .Y(\u_neuron.u_syn/_358_ ),
    .A1(\u_neuron.u_syn/_232_ ),
    .A2(\u_neuron.u_syn/_307_ ));
 sg13g2_a221oi_1 \u_neuron.u_syn/_756_  (.B2(\u_neuron.u_syn/_358_ ),
    .C1(\u_neuron.u_syn/_352_ ),
    .B1(\u_neuron.u_syn/_351_ ),
    .A1(\u_neuron.u_syn/_235_ ),
    .Y(\u_neuron.u_syn/_359_ ),
    .A2(\u_neuron.u_syn/_309_ ));
 sg13g2_o21ai_1 \u_neuron.u_syn/_757_  (.B1(net467),
    .Y(\u_neuron.u_syn/_360_ ),
    .A1(\u_neuron.ltd_wdata[1] ),
    .A2(\u_neuron.u_syn/_353_ ));
 sg13g2_nand2_1 \u_neuron.u_syn/_758_  (.Y(\u_neuron.u_syn/_361_ ),
    .A(net415),
    .B(net193));
 sg13g2_o21ai_1 \u_neuron.u_syn/_759_  (.B1(\u_neuron.u_syn/_361_ ),
    .Y(\u_neuron.u_syn/_025_ ),
    .A1(\u_neuron.u_syn/_359_ ),
    .A2(\u_neuron.u_syn/_360_ ));
 sg13g2_nand4_1 \u_neuron.u_syn/_760_  (.B(net405),
    .C(net359),
    .A(\u_neuron.pending_widx[3] ),
    .Y(\u_neuron.u_syn/_362_ ),
    .D(\u_neuron.u_syn/_148_ ));
 sg13g2_nand4_1 \u_neuron.u_syn/_761_  (.B(\u_neuron.ltp_idx[2] ),
    .C(\u_neuron.ltp_we ),
    .A(\u_neuron.ltp_idx[3] ),
    .Y(\u_neuron.u_syn/_363_ ),
    .D(\u_neuron.u_syn/_153_ ));
 sg13g2_o21ai_1 \u_neuron.u_syn/_762_  (.B1(\u_neuron.u_syn/_363_ ),
    .Y(\u_neuron.u_syn/_364_ ),
    .A1(\u_neuron.u_syn/_041_ ),
    .A2(\u_neuron.u_syn/_362_ ));
 sg13g2_a21o_1 \u_neuron.u_syn/_763_  (.A2(\u_neuron.u_syn/_362_ ),
    .A1(net197),
    .B1(\u_neuron.u_syn/_364_ ),
    .X(\u_neuron.u_syn/_365_ ));
 sg13g2_nor2_1 \u_neuron.u_syn/_764_  (.A(\u_neuron.ltp_wdata[0] ),
    .B(\u_neuron.u_syn/_363_ ),
    .Y(\u_neuron.u_syn/_366_ ));
 sg13g2_a21oi_1 \u_neuron.u_syn/_765_  (.A1(\u_neuron.u_syn/_246_ ),
    .A2(net318),
    .Y(\u_neuron.u_syn/_367_ ),
    .B1(\u_neuron.u_syn/_366_ ));
 sg13g2_o21ai_1 \u_neuron.u_syn/_766_  (.B1(net467),
    .Y(\u_neuron.u_syn/_368_ ),
    .A1(\u_neuron.u_syn/_248_ ),
    .A2(\u_neuron.u_syn/_313_ ));
 sg13g2_a21oi_1 \u_neuron.u_syn/_767_  (.A1(\u_neuron.u_syn/_365_ ),
    .A2(\u_neuron.u_syn/_367_ ),
    .Y(\u_neuron.u_syn/_369_ ),
    .B1(\u_neuron.u_syn/_368_ ));
 sg13g2_a21oi_1 \u_neuron.u_syn/_768_  (.A1(net415),
    .A2(\u_neuron.u_syn/_072_ ),
    .Y(\u_neuron.u_syn/_026_ ),
    .B1(\u_neuron.u_syn/_369_ ));
 sg13g2_o21ai_1 \u_neuron.u_syn/_769_  (.B1(\u_neuron.u_syn/_363_ ),
    .Y(\u_neuron.u_syn/_370_ ),
    .A1(\u_neuron.u_syn/_051_ ),
    .A2(\u_neuron.u_syn/_362_ ));
 sg13g2_a21o_1 \u_neuron.u_syn/_770_  (.A2(\u_neuron.u_syn/_362_ ),
    .A1(net198),
    .B1(\u_neuron.u_syn/_370_ ),
    .X(\u_neuron.u_syn/_371_ ));
 sg13g2_nor2_1 \u_neuron.u_syn/_771_  (.A(net333),
    .B(\u_neuron.u_syn/_363_ ),
    .Y(\u_neuron.u_syn/_372_ ));
 sg13g2_a21oi_1 \u_neuron.u_syn/_772_  (.A1(\u_neuron.u_syn/_246_ ),
    .A2(net318),
    .Y(\u_neuron.u_syn/_373_ ),
    .B1(\u_neuron.u_syn/_372_ ));
 sg13g2_o21ai_1 \u_neuron.u_syn/_773_  (.B1(net467),
    .Y(\u_neuron.u_syn/_374_ ),
    .A1(\u_neuron.u_syn/_255_ ),
    .A2(\u_neuron.u_syn/_313_ ));
 sg13g2_a21oi_1 \u_neuron.u_syn/_774_  (.A1(\u_neuron.u_syn/_371_ ),
    .A2(\u_neuron.u_syn/_373_ ),
    .Y(\u_neuron.u_syn/_375_ ),
    .B1(\u_neuron.u_syn/_374_ ));
 sg13g2_a21oi_1 \u_neuron.u_syn/_775_  (.A1(net415),
    .A2(\u_neuron.u_syn/_073_ ),
    .Y(\u_neuron.u_syn/_027_ ),
    .B1(\u_neuron.u_syn/_375_ ));
 sg13g2_nand4_1 \u_neuron.u_syn/_776_  (.B(net404),
    .C(net357),
    .A(\u_neuron.pending_widx[3] ),
    .Y(\u_neuron.u_syn/_376_ ),
    .D(\u_neuron.u_syn/_175_ ));
 sg13g2_nor4_2 \u_neuron.u_syn/_777_  (.A(\u_neuron.u_syn/_042_ ),
    .B(\u_neuron.u_syn/_043_ ),
    .C(net315),
    .Y(\u_neuron.u_syn/_377_ ),
    .D(\u_neuron.u_syn/_178_ ));
 sg13g2_a21oi_1 \u_neuron.u_syn/_778_  (.A1(net189),
    .A2(\u_neuron.u_syn/_376_ ),
    .Y(\u_neuron.u_syn/_378_ ),
    .B1(\u_neuron.u_syn/_377_ ));
 sg13g2_o21ai_1 \u_neuron.u_syn/_779_  (.B1(\u_neuron.u_syn/_378_ ),
    .Y(\u_neuron.u_syn/_379_ ),
    .A1(\u_neuron.u_syn/_261_ ),
    .A2(\u_neuron.u_syn/_307_ ));
 sg13g2_a22oi_1 \u_neuron.u_syn/_780_  (.Y(\u_neuron.u_syn/_380_ ),
    .B1(\u_neuron.u_syn/_377_ ),
    .B2(\u_neuron.u_syn/_183_ ),
    .A2(net317),
    .A1(\u_neuron.u_syn/_263_ ));
 sg13g2_a221oi_1 \u_neuron.u_syn/_781_  (.B2(\u_neuron.u_syn/_380_ ),
    .C1(net412),
    .B1(\u_neuron.u_syn/_379_ ),
    .A1(\u_neuron.u_syn/_266_ ),
    .Y(\u_neuron.u_syn/_381_ ),
    .A2(net317));
 sg13g2_a21oi_1 \u_neuron.u_syn/_782_  (.A1(net412),
    .A2(\u_neuron.u_syn/_074_ ),
    .Y(\u_neuron.u_syn/_028_ ),
    .B1(\u_neuron.u_syn/_381_ ));
 sg13g2_nand2_1 \u_neuron.u_syn/_783_  (.Y(\u_neuron.u_syn/_382_ ),
    .A(net211),
    .B(\u_neuron.u_syn/_376_ ));
 sg13g2_o21ai_1 \u_neuron.u_syn/_784_  (.B1(\u_neuron.u_syn/_382_ ),
    .Y(\u_neuron.u_syn/_383_ ),
    .A1(\u_neuron.u_syn/_269_ ),
    .A2(\u_neuron.u_syn/_307_ ));
 sg13g2_a22oi_1 \u_neuron.u_syn/_785_  (.Y(\u_neuron.u_syn/_384_ ),
    .B1(\u_neuron.u_syn/_377_ ),
    .B2(\u_neuron.u_syn/_192_ ),
    .A2(net317),
    .A1(\u_neuron.u_syn/_263_ ));
 sg13g2_o21ai_1 \u_neuron.u_syn/_786_  (.B1(\u_neuron.u_syn/_384_ ),
    .Y(\u_neuron.u_syn/_385_ ),
    .A1(\u_neuron.u_syn/_377_ ),
    .A2(\u_neuron.u_syn/_383_ ));
 sg13g2_a21oi_1 \u_neuron.u_syn/_787_  (.A1(\u_neuron.u_syn/_273_ ),
    .A2(net317),
    .Y(\u_neuron.u_syn/_386_ ),
    .B1(net412));
 sg13g2_a22oi_1 \u_neuron.u_syn/_788_  (.Y(\u_neuron.u_syn/_029_ ),
    .B1(\u_neuron.u_syn/_385_ ),
    .B2(\u_neuron.u_syn/_386_ ),
    .A2(\u_neuron.u_syn/_075_ ),
    .A1(net412));
 sg13g2_nand4_1 \u_neuron.u_syn/_789_  (.B(net405),
    .C(net357),
    .A(\u_neuron.pending_widx[3] ),
    .Y(\u_neuron.u_syn/_387_ ),
    .D(\u_neuron.u_syn/_197_ ));
 sg13g2_nand2_1 \u_neuron.u_syn/_790_  (.Y(\u_neuron.u_syn/_388_ ),
    .A(net194),
    .B(\u_neuron.u_syn/_387_ ));
 sg13g2_nor4_2 \u_neuron.u_syn/_791_  (.A(\u_neuron.u_syn/_042_ ),
    .B(\u_neuron.u_syn/_043_ ),
    .C(net315),
    .Y(\u_neuron.u_syn/_389_ ),
    .D(\u_neuron.u_syn/_201_ ));
 sg13g2_o21ai_1 \u_neuron.u_syn/_792_  (.B1(\u_neuron.u_syn/_388_ ),
    .Y(\u_neuron.u_syn/_390_ ),
    .A1(\u_neuron.u_syn/_278_ ),
    .A2(\u_neuron.u_syn/_307_ ));
 sg13g2_nand2_1 \u_neuron.u_syn/_793_  (.Y(\u_neuron.u_syn/_391_ ),
    .A(\u_neuron.u_syn/_281_ ),
    .B(net316));
 sg13g2_a22oi_1 \u_neuron.u_syn/_794_  (.Y(\u_neuron.u_syn/_392_ ),
    .B1(\u_neuron.u_syn/_389_ ),
    .B2(\u_neuron.u_syn/_044_ ),
    .A2(net317),
    .A1(\u_neuron.u_syn/_281_ ));
 sg13g2_o21ai_1 \u_neuron.u_syn/_795_  (.B1(\u_neuron.u_syn/_392_ ),
    .Y(\u_neuron.u_syn/_393_ ),
    .A1(\u_neuron.u_syn/_389_ ),
    .A2(\u_neuron.u_syn/_390_ ));
 sg13g2_a21oi_1 \u_neuron.u_syn/_796_  (.A1(\u_neuron.u_syn/_285_ ),
    .A2(net317),
    .Y(\u_neuron.u_syn/_394_ ),
    .B1(net412));
 sg13g2_a22oi_1 \u_neuron.u_syn/_797_  (.Y(\u_neuron.u_syn/_030_ ),
    .B1(\u_neuron.u_syn/_393_ ),
    .B2(\u_neuron.u_syn/_394_ ),
    .A2(\u_neuron.u_syn/_076_ ),
    .A1(net412));
 sg13g2_nor2b_1 \u_neuron.u_syn/_798_  (.A(net146),
    .B_N(\u_neuron.u_syn/_387_ ),
    .Y(\u_neuron.u_syn/_395_ ));
 sg13g2_nor2_1 \u_neuron.u_syn/_799_  (.A(\u_neuron.cfg_arg[1] ),
    .B(\u_neuron.u_syn/_387_ ),
    .Y(\u_neuron.u_syn/_396_ ));
 sg13g2_nor3_1 \u_neuron.u_syn/_800_  (.A(\u_neuron.u_syn/_389_ ),
    .B(\u_neuron.u_syn/_395_ ),
    .C(\u_neuron.u_syn/_396_ ),
    .Y(\u_neuron.u_syn/_397_ ));
 sg13g2_a221oi_1 \u_neuron.u_syn/_801_  (.B2(net333),
    .C1(\u_neuron.u_syn/_397_ ),
    .B1(\u_neuron.u_syn/_389_ ),
    .A1(\u_neuron.u_syn/_281_ ),
    .Y(\u_neuron.u_syn/_398_ ),
    .A2(net317));
 sg13g2_o21ai_1 \u_neuron.u_syn/_802_  (.B1(net466),
    .Y(\u_neuron.u_syn/_399_ ),
    .A1(net331),
    .A2(\u_neuron.u_syn/_391_ ));
 sg13g2_nand2_1 \u_neuron.u_syn/_803_  (.Y(\u_neuron.u_syn/_400_ ),
    .A(net412),
    .B(net146));
 sg13g2_o21ai_1 \u_neuron.u_syn/_804_  (.B1(\u_neuron.u_syn/_400_ ),
    .Y(\u_neuron.u_syn/_031_ ),
    .A1(\u_neuron.u_syn/_398_ ),
    .A2(\u_neuron.u_syn/_399_ ));
 sg13g2_nand2_2 \u_neuron.u_syn/_805_  (.Y(\u_neuron.u_syn/_401_ ),
    .A(_000_),
    .B(net469));
 sg13g2_nor2_1 \u_neuron.u_syn/_806_  (.A(\u_neuron.cfg_arg[0] ),
    .B(\u_neuron.u_syn/_401_ ),
    .Y(\u_neuron.u_syn/_402_ ));
 sg13g2_a21oi_1 \u_neuron.u_syn/_807_  (.A1(\u_neuron.u_syn/_039_ ),
    .A2(\u_neuron.u_syn/_401_ ),
    .Y(\u_neuron.u_syn/_032_ ),
    .B1(\u_neuron.u_syn/_402_ ));
 sg13g2_nor2_1 \u_neuron.u_syn/_808_  (.A(\u_neuron.cfg_arg[1] ),
    .B(\u_neuron.u_syn/_401_ ),
    .Y(\u_neuron.u_syn/_403_ ));
 sg13g2_a21oi_1 \u_neuron.u_syn/_809_  (.A1(\u_neuron.u_syn/_038_ ),
    .A2(\u_neuron.u_syn/_401_ ),
    .Y(\u_neuron.u_syn/_033_ ),
    .B1(net229));
 sg13g2_mux2_1 \u_neuron.u_syn/_810_  (.A0(\u_neuron.cfg_arg[2] ),
    .A1(net407),
    .S(\u_neuron.u_syn/_401_ ),
    .X(\u_neuron.u_syn/_034_ ));
 sg13g2_nor2_1 \u_neuron.u_syn/_811_  (.A(\u_neuron.cfg_arg[3] ),
    .B(\u_neuron.u_syn/_401_ ),
    .Y(\u_neuron.u_syn/_404_ ));
 sg13g2_a21oi_1 \u_neuron.u_syn/_812_  (.A1(\u_neuron.u_syn/_037_ ),
    .A2(\u_neuron.u_syn/_401_ ),
    .Y(\u_neuron.u_syn/_035_ ),
    .B1(\u_neuron.u_syn/_404_ ));
 sg13g2_dfrbpq_2 \u_neuron.u_syn/_813_  (.RESET_B(net456),
    .D(\u_neuron.u_syn/_000_ ),
    .Q(\u_neuron.wtab[0] ),
    .CLK(clknet_5_6__leaf_clk));
 sg13g2_dfrbpq_2 \u_neuron.u_syn/_814_  (.RESET_B(net456),
    .D(\u_neuron.u_syn/_001_ ),
    .Q(\u_neuron.wtab[1] ),
    .CLK(clknet_5_30__leaf_clk));
 sg13g2_dfrbpq_2 \u_neuron.u_syn/_815_  (.RESET_B(net456),
    .D(\u_neuron.u_syn/_002_ ),
    .Q(\u_neuron.wtab[2] ),
    .CLK(clknet_5_30__leaf_clk));
 sg13g2_dfrbpq_2 \u_neuron.u_syn/_816_  (.RESET_B(net460),
    .D(\u_neuron.u_syn/_003_ ),
    .Q(\u_neuron.wtab[3] ),
    .CLK(clknet_5_28__leaf_clk));
 sg13g2_dfrbpq_2 \u_neuron.u_syn/_817_  (.RESET_B(net447),
    .D(\u_neuron.u_syn/_004_ ),
    .Q(\u_neuron.wtab[4] ),
    .CLK(clknet_5_13__leaf_clk));
 sg13g2_dfrbpq_2 \u_neuron.u_syn/_818_  (.RESET_B(net445),
    .D(\u_neuron.u_syn/_005_ ),
    .Q(\u_neuron.wtab[5] ),
    .CLK(clknet_5_5__leaf_clk));
 sg13g2_dfrbpq_2 \u_neuron.u_syn/_819_  (.RESET_B(net463),
    .D(\u_neuron.u_syn/_006_ ),
    .Q(\u_neuron.wtab[6] ),
    .CLK(clknet_5_30__leaf_clk));
 sg13g2_dfrbpq_2 \u_neuron.u_syn/_820_  (.RESET_B(net463),
    .D(\u_neuron.u_syn/_007_ ),
    .Q(\u_neuron.wtab[7] ),
    .CLK(clknet_5_30__leaf_clk));
 sg13g2_dfrbpq_2 \u_neuron.u_syn/_821_  (.RESET_B(net457),
    .D(\u_neuron.u_syn/_008_ ),
    .Q(\u_neuron.wtab[8] ),
    .CLK(clknet_5_27__leaf_clk));
 sg13g2_dfrbpq_2 \u_neuron.u_syn/_822_  (.RESET_B(net457),
    .D(\u_neuron.u_syn/_009_ ),
    .Q(\u_neuron.wtab[9] ),
    .CLK(clknet_5_26__leaf_clk));
 sg13g2_dfrbpq_2 \u_neuron.u_syn/_823_  (.RESET_B(net463),
    .D(\u_neuron.u_syn/_010_ ),
    .Q(\u_neuron.wtab[10] ),
    .CLK(clknet_5_30__leaf_clk));
 sg13g2_dfrbpq_2 \u_neuron.u_syn/_824_  (.RESET_B(net456),
    .D(\u_neuron.u_syn/_011_ ),
    .Q(\u_neuron.wtab[11] ),
    .CLK(clknet_5_26__leaf_clk));
 sg13g2_dfrbpq_2 \u_neuron.u_syn/_825_  (.RESET_B(net446),
    .D(\u_neuron.u_syn/_012_ ),
    .Q(\u_neuron.wtab[12] ),
    .CLK(clknet_5_15__leaf_clk));
 sg13g2_dfrbpq_2 \u_neuron.u_syn/_826_  (.RESET_B(net446),
    .D(\u_neuron.u_syn/_013_ ),
    .Q(\u_neuron.wtab[13] ),
    .CLK(clknet_5_15__leaf_clk));
 sg13g2_dfrbpq_2 \u_neuron.u_syn/_827_  (.RESET_B(net446),
    .D(net187),
    .Q(\u_neuron.wtab[14] ),
    .CLK(clknet_5_26__leaf_clk));
 sg13g2_dfrbpq_2 \u_neuron.u_syn/_828_  (.RESET_B(net457),
    .D(\u_neuron.u_syn/_015_ ),
    .Q(\u_neuron.wtab[15] ),
    .CLK(clknet_5_26__leaf_clk));
 sg13g2_dfrbpq_2 \u_neuron.u_syn/_829_  (.RESET_B(net445),
    .D(\u_neuron.u_syn/_016_ ),
    .Q(\u_neuron.wtab[16] ),
    .CLK(clknet_5_13__leaf_clk));
 sg13g2_dfrbpq_2 \u_neuron.u_syn/_830_  (.RESET_B(net445),
    .D(\u_neuron.u_syn/_017_ ),
    .Q(\u_neuron.wtab[17] ),
    .CLK(clknet_5_14__leaf_clk));
 sg13g2_dfrbpq_2 \u_neuron.u_syn/_831_  (.RESET_B(net445),
    .D(\u_neuron.u_syn/_018_ ),
    .Q(\u_neuron.wtab[18] ),
    .CLK(clknet_5_6__leaf_clk));
 sg13g2_dfrbpq_1 \u_neuron.u_syn/_832_  (.RESET_B(net446),
    .D(\u_neuron.u_syn/_019_ ),
    .Q(\u_neuron.wtab[19] ),
    .CLK(clknet_5_14__leaf_clk));
 sg13g2_dfrbpq_2 \u_neuron.u_syn/_833_  (.RESET_B(net445),
    .D(\u_neuron.u_syn/_020_ ),
    .Q(\u_neuron.wtab[20] ),
    .CLK(clknet_5_4__leaf_clk));
 sg13g2_dfrbpq_2 \u_neuron.u_syn/_834_  (.RESET_B(net445),
    .D(\u_neuron.u_syn/_021_ ),
    .Q(\u_neuron.wtab[21] ),
    .CLK(clknet_5_13__leaf_clk));
 sg13g2_dfrbpq_2 \u_neuron.u_syn/_835_  (.RESET_B(net445),
    .D(\u_neuron.u_syn/_022_ ),
    .Q(\u_neuron.wtab[22] ),
    .CLK(clknet_5_14__leaf_clk));
 sg13g2_dfrbpq_2 \u_neuron.u_syn/_836_  (.RESET_B(net445),
    .D(\u_neuron.u_syn/_023_ ),
    .Q(\u_neuron.wtab[23] ),
    .CLK(clknet_5_14__leaf_clk));
 sg13g2_dfrbpq_2 \u_neuron.u_syn/_837_  (.RESET_B(net457),
    .D(\u_neuron.u_syn/_024_ ),
    .Q(\u_neuron.wtab[24] ),
    .CLK(clknet_5_27__leaf_clk));
 sg13g2_dfrbpq_2 \u_neuron.u_syn/_838_  (.RESET_B(net457),
    .D(\u_neuron.u_syn/_025_ ),
    .Q(\u_neuron.wtab[25] ),
    .CLK(clknet_5_26__leaf_clk));
 sg13g2_dfrbpq_2 \u_neuron.u_syn/_839_  (.RESET_B(net456),
    .D(\u_neuron.u_syn/_026_ ),
    .Q(\u_neuron.wtab[26] ),
    .CLK(clknet_5_27__leaf_clk));
 sg13g2_dfrbpq_2 \u_neuron.u_syn/_840_  (.RESET_B(net457),
    .D(\u_neuron.u_syn/_027_ ),
    .Q(\u_neuron.wtab[27] ),
    .CLK(clknet_5_24__leaf_clk));
 sg13g2_dfrbpq_2 \u_neuron.u_syn/_841_  (.RESET_B(net446),
    .D(\u_neuron.u_syn/_028_ ),
    .Q(\u_neuron.wtab[28] ),
    .CLK(clknet_5_15__leaf_clk));
 sg13g2_dfrbpq_2 \u_neuron.u_syn/_842_  (.RESET_B(net447),
    .D(\u_neuron.u_syn/_029_ ),
    .Q(\u_neuron.wtab[29] ),
    .CLK(clknet_5_14__leaf_clk));
 sg13g2_dfrbpq_2 \u_neuron.u_syn/_843_  (.RESET_B(net446),
    .D(\u_neuron.u_syn/_030_ ),
    .Q(\u_neuron.wtab[30] ),
    .CLK(clknet_5_15__leaf_clk));
 sg13g2_dfrbpq_2 \u_neuron.u_syn/_844_  (.RESET_B(net446),
    .D(\u_neuron.u_syn/_031_ ),
    .Q(\u_neuron.wtab[31] ),
    .CLK(clknet_5_15__leaf_clk));
 sg13g2_dfrbpq_2 \u_neuron.u_syn/_845_  (.RESET_B(net456),
    .D(net227),
    .Q(\u_neuron.pending_widx[0] ),
    .CLK(clknet_5_6__leaf_clk));
 sg13g2_dfrbpq_2 \u_neuron.u_syn/_846_  (.RESET_B(net456),
    .D(net230),
    .Q(\u_neuron.pending_widx[1] ),
    .CLK(clknet_5_6__leaf_clk));
 sg13g2_dfrbpq_1 \u_neuron.u_syn/_847_  (.RESET_B(net460),
    .D(net220),
    .Q(\u_neuron.pending_widx[2] ),
    .CLK(clknet_5_28__leaf_clk));
 sg13g2_dfrbpq_2 \u_neuron.u_syn/_848_  (.RESET_B(net456),
    .D(net216),
    .Q(\u_neuron.pending_widx[3] ),
    .CLK(clknet_5_28__leaf_clk));
 sg13g2_inv_1 \u_neuron.u_td/_096_  (.Y(\u_neuron.u_td/_058_ ),
    .A(net182));
 sg13g2_inv_1 \u_neuron.u_td/_097_  (.Y(\u_neuron.u_td/_059_ ),
    .A(net166));
 sg13g2_inv_1 \u_neuron.u_td/_098_  (.Y(\u_neuron.u_td/_060_ ),
    .A(net170));
 sg13g2_inv_1 \u_neuron.u_td/_099_  (.Y(\u_neuron.u_td/_061_ ),
    .A(net156));
 sg13g2_inv_1 \u_neuron.u_td/_100_  (.Y(\u_neuron.u_td/_062_ ),
    .A(net162));
 sg13g2_inv_1 \u_neuron.u_td/_101_  (.Y(\u_neuron.u_td/_063_ ),
    .A(net178));
 sg13g2_inv_1 \u_neuron.u_td/_102_  (.Y(\u_neuron.u_td/_064_ ),
    .A(\u_neuron.stream_act ));
 sg13g2_nor2b_1 \u_neuron.u_td/_103_  (.A(\u_neuron.td_prev[1] ),
    .B_N(\u_neuron.td_curr[1] ),
    .Y(\u_neuron.u_td/_065_ ));
 sg13g2_nand2b_2 \u_neuron.u_td/_104_  (.Y(\u_neuron.u_td/_066_ ),
    .B(\u_neuron.td_prev[0] ),
    .A_N(\u_neuron.td_curr[0] ));
 sg13g2_xnor2_1 \u_neuron.u_td/_105_  (.Y(\u_neuron.u_td/_067_ ),
    .A(\u_neuron.td_prev[1] ),
    .B(\u_neuron.td_curr[1] ));
 sg13g2_a21oi_1 \u_neuron.u_td/_106_  (.A1(\u_neuron.u_td/_066_ ),
    .A2(\u_neuron.u_td/_067_ ),
    .Y(\u_neuron.u_td/_068_ ),
    .B1(\u_neuron.u_td/_065_ ));
 sg13g2_a21o_1 \u_neuron.u_td/_107_  (.A2(\u_neuron.u_td/_067_ ),
    .A1(\u_neuron.u_td/_066_ ),
    .B1(\u_neuron.u_td/_065_ ),
    .X(\u_neuron.u_td/_069_ ));
 sg13g2_nor2b_1 \u_neuron.u_td/_108_  (.A(\u_neuron.td_prev[2] ),
    .B_N(\u_neuron.td_curr[2] ),
    .Y(\u_neuron.u_td/_070_ ));
 sg13g2_xnor2_1 \u_neuron.u_td/_109_  (.Y(\u_neuron.u_td/_071_ ),
    .A(\u_neuron.td_prev[2] ),
    .B(\u_neuron.td_curr[2] ));
 sg13g2_nor2b_1 \u_neuron.u_td/_110_  (.A(\u_neuron.td_prev[3] ),
    .B_N(\u_neuron.td_curr[3] ),
    .Y(\u_neuron.u_td/_072_ ));
 sg13g2_nand2b_1 \u_neuron.u_td/_111_  (.Y(\u_neuron.u_td/_073_ ),
    .B(\u_neuron.td_prev[3] ),
    .A_N(\u_neuron.td_curr[3] ));
 sg13g2_xnor2_1 \u_neuron.u_td/_112_  (.Y(\u_neuron.u_td/_074_ ),
    .A(\u_neuron.td_prev[3] ),
    .B(\u_neuron.td_curr[3] ));
 sg13g2_nand2_1 \u_neuron.u_td/_113_  (.Y(\u_neuron.u_td/_075_ ),
    .A(\u_neuron.u_td/_071_ ),
    .B(\u_neuron.u_td/_074_ ));
 sg13g2_a21oi_1 \u_neuron.u_td/_114_  (.A1(\u_neuron.u_td/_070_ ),
    .A2(\u_neuron.u_td/_073_ ),
    .Y(\u_neuron.u_td/_076_ ),
    .B1(\u_neuron.u_td/_072_ ));
 sg13g2_o21ai_1 \u_neuron.u_td/_115_  (.B1(\u_neuron.u_td/_076_ ),
    .Y(\u_neuron.u_td/_077_ ),
    .A1(\u_neuron.u_td/_068_ ),
    .A2(\u_neuron.u_td/_075_ ));
 sg13g2_nand2b_1 \u_neuron.u_td/_116_  (.Y(\u_neuron.u_td/_078_ ),
    .B(\u_neuron.td_prev[5] ),
    .A_N(\u_neuron.td_curr[5] ));
 sg13g2_nor2b_1 \u_neuron.u_td/_117_  (.A(\u_neuron.td_prev[5] ),
    .B_N(\u_neuron.td_curr[5] ),
    .Y(\u_neuron.u_td/_079_ ));
 sg13g2_xor2_1 \u_neuron.u_td/_118_  (.B(\u_neuron.td_curr[5] ),
    .A(\u_neuron.td_prev[5] ),
    .X(\u_neuron.u_td/_080_ ));
 sg13g2_nor2b_1 \u_neuron.u_td/_119_  (.A(\u_neuron.td_prev[4] ),
    .B_N(\u_neuron.td_curr[4] ),
    .Y(\u_neuron.u_td/_081_ ));
 sg13g2_nand2b_1 \u_neuron.u_td/_120_  (.Y(\u_neuron.u_td/_082_ ),
    .B(\u_neuron.td_curr[4] ),
    .A_N(\u_neuron.td_prev[4] ));
 sg13g2_xnor2_1 \u_neuron.u_td/_121_  (.Y(\u_neuron.u_td/_083_ ),
    .A(\u_neuron.td_prev[4] ),
    .B(\u_neuron.td_curr[4] ));
 sg13g2_nor2b_1 \u_neuron.u_td/_122_  (.A(\u_neuron.u_td/_080_ ),
    .B_N(\u_neuron.u_td/_083_ ),
    .Y(\u_neuron.u_td/_084_ ));
 sg13g2_a21oi_1 \u_neuron.u_td/_123_  (.A1(\u_neuron.u_td/_078_ ),
    .A2(\u_neuron.u_td/_081_ ),
    .Y(\u_neuron.u_td/_085_ ),
    .B1(\u_neuron.u_td/_079_ ));
 sg13g2_inv_1 \u_neuron.u_td/_124_  (.Y(\u_neuron.u_td/_086_ ),
    .A(\u_neuron.u_td/_085_ ));
 sg13g2_nor2b_1 \u_neuron.u_td/_125_  (.A(\u_neuron.td_prev[7] ),
    .B_N(\u_neuron.td_curr[7] ),
    .Y(\u_neuron.u_td/_087_ ));
 sg13g2_nand2b_1 \u_neuron.u_td/_126_  (.Y(\u_neuron.u_td/_088_ ),
    .B(\u_neuron.td_prev[7] ),
    .A_N(\u_neuron.td_curr[7] ));
 sg13g2_nor2b_1 \u_neuron.u_td/_127_  (.A(\u_neuron.td_prev[6] ),
    .B_N(\u_neuron.td_curr[6] ),
    .Y(\u_neuron.u_td/_089_ ));
 sg13g2_a21oi_1 \u_neuron.u_td/_128_  (.A1(\u_neuron.u_td/_088_ ),
    .A2(\u_neuron.u_td/_089_ ),
    .Y(\u_neuron.u_td/_090_ ),
    .B1(\u_neuron.u_td/_087_ ));
 sg13g2_nand2_1 \u_neuron.u_td/_129_  (.Y(\u_neuron.u_td/_091_ ),
    .A(\u_neuron.u_td/_085_ ),
    .B(\u_neuron.u_td/_090_ ));
 sg13g2_a21oi_2 \u_neuron.u_td/_130_  (.B1(\u_neuron.u_td/_091_ ),
    .Y(\u_neuron.u_td/_092_ ),
    .A2(\u_neuron.u_td/_084_ ),
    .A1(\u_neuron.u_td/_077_ ));
 sg13g2_nand2b_1 \u_neuron.u_td/_131_  (.Y(\u_neuron.u_td/_093_ ),
    .B(\u_neuron.td_prev[6] ),
    .A_N(\u_neuron.td_curr[6] ));
 sg13g2_o21ai_1 \u_neuron.u_td/_132_  (.B1(\u_neuron.u_td/_088_ ),
    .Y(\u_neuron.u_td/_094_ ),
    .A1(\u_neuron.u_td/_087_ ),
    .A2(\u_neuron.u_td/_093_ ));
 sg13g2_nor2_1 \u_neuron.u_td/_133_  (.A(\u_neuron.u_td/_092_ ),
    .B(\u_neuron.u_td/_094_ ),
    .Y(\u_neuron.u_td/_095_ ));
 sg13g2_a21oi_1 \u_neuron.u_td/_134_  (.A1(\u_neuron.u_td/_069_ ),
    .A2(\u_neuron.u_td/_071_ ),
    .Y(\u_neuron.u_td/_000_ ),
    .B1(\u_neuron.u_td/_070_ ));
 sg13g2_xor2_1 \u_neuron.u_td/_135_  (.B(\u_neuron.u_td/_000_ ),
    .A(\u_neuron.u_td/_074_ ),
    .X(\u_neuron.u_td/_001_ ));
 sg13g2_nor3_2 \u_neuron.u_td/_136_  (.A(\u_neuron.u_td/_092_ ),
    .B(\u_neuron.u_td/_094_ ),
    .C(\u_neuron.u_td/_001_ ),
    .Y(\u_neuron.td_emit_data[3] ));
 sg13g2_xnor2_1 \u_neuron.u_td/_137_  (.Y(\u_neuron.u_td/_002_ ),
    .A(\u_neuron.td_prev[0] ),
    .B(\u_neuron.td_curr[0] ));
 sg13g2_nor3_1 \u_neuron.u_td/_138_  (.A(\u_neuron.u_td/_092_ ),
    .B(\u_neuron.u_td/_094_ ),
    .C(\u_neuron.u_td/_002_ ),
    .Y(\u_neuron.td_emit_data[0] ));
 sg13g2_xnor2_1 \u_neuron.u_td/_139_  (.Y(\u_neuron.u_td/_003_ ),
    .A(\u_neuron.u_td/_066_ ),
    .B(\u_neuron.u_td/_067_ ));
 sg13g2_nor3_2 \u_neuron.u_td/_140_  (.A(\u_neuron.u_td/_092_ ),
    .B(\u_neuron.u_td/_094_ ),
    .C(\u_neuron.u_td/_003_ ),
    .Y(\u_neuron.td_emit_data[1] ));
 sg13g2_xnor2_1 \u_neuron.u_td/_141_  (.Y(\u_neuron.u_td/_004_ ),
    .A(\u_neuron.u_td/_069_ ),
    .B(\u_neuron.u_td/_071_ ));
 sg13g2_nor3_2 \u_neuron.u_td/_142_  (.A(\u_neuron.u_td/_092_ ),
    .B(\u_neuron.u_td/_094_ ),
    .C(\u_neuron.u_td/_004_ ),
    .Y(\u_neuron.td_emit_data[2] ));
 sg13g2_nand2_1 \u_neuron.u_td/_143_  (.Y(\u_neuron.u_td/_005_ ),
    .A(net385),
    .B(net355));
 sg13g2_or2_1 \u_neuron.u_td/_144_  (.X(\u_neuron.u_td/_006_ ),
    .B(net328),
    .A(net417));
 sg13g2_nand2_1 \u_neuron.u_td/_145_  (.Y(\u_neuron.u_td/_007_ ),
    .A(\u_neuron.u_td/_077_ ),
    .B(\u_neuron.u_td/_083_ ));
 sg13g2_xnor2_1 \u_neuron.u_td/_146_  (.Y(\u_neuron.u_td/_008_ ),
    .A(\u_neuron.u_td/_077_ ),
    .B(\u_neuron.u_td/_083_ ));
 sg13g2_nor3_1 \u_neuron.u_td/_147_  (.A(\u_neuron.u_td/_092_ ),
    .B(\u_neuron.u_td/_094_ ),
    .C(\u_neuron.u_td/_008_ ),
    .Y(\u_neuron.u_td/_009_ ));
 sg13g2_nor3_1 \u_neuron.u_td/_148_  (.A(\u_neuron.td_emit_data[3] ),
    .B(\u_neuron.td_emit_data[2] ),
    .C(\u_neuron.u_td/_009_ ),
    .Y(\u_neuron.u_td/_010_ ));
 sg13g2_nand2b_1 \u_neuron.u_td/_149_  (.Y(\u_neuron.u_td/_011_ ),
    .B(\u_neuron.u_td/_093_ ),
    .A_N(\u_neuron.u_td/_089_ ));
 sg13g2_a21oi_1 \u_neuron.u_td/_150_  (.A1(\u_neuron.u_td/_077_ ),
    .A2(\u_neuron.u_td/_084_ ),
    .Y(\u_neuron.u_td/_012_ ),
    .B1(\u_neuron.u_td/_086_ ));
 sg13g2_nand2_1 \u_neuron.u_td/_151_  (.Y(\u_neuron.u_td/_013_ ),
    .A(\u_neuron.u_td/_011_ ),
    .B(\u_neuron.u_td/_012_ ));
 sg13g2_nor2_1 \u_neuron.u_td/_152_  (.A(\u_neuron.u_td/_011_ ),
    .B(\u_neuron.u_td/_012_ ),
    .Y(\u_neuron.u_td/_014_ ));
 sg13g2_nand3b_1 \u_neuron.u_td/_153_  (.B(\u_neuron.u_td/_095_ ),
    .C(\u_neuron.u_td/_013_ ),
    .Y(\u_neuron.u_td/_015_ ),
    .A_N(\u_neuron.u_td/_014_ ));
 sg13g2_o21ai_1 \u_neuron.u_td/_154_  (.B1(\u_neuron.u_td/_087_ ),
    .Y(\u_neuron.u_td/_016_ ),
    .A1(\u_neuron.u_td/_089_ ),
    .A2(\u_neuron.u_td/_014_ ));
 sg13g2_nand3_1 \u_neuron.u_td/_155_  (.B(\u_neuron.u_td/_082_ ),
    .C(\u_neuron.u_td/_007_ ),
    .A(\u_neuron.u_td/_080_ ),
    .Y(\u_neuron.u_td/_017_ ));
 sg13g2_a21o_1 \u_neuron.u_td/_156_  (.A2(\u_neuron.u_td/_007_ ),
    .A1(\u_neuron.u_td/_082_ ),
    .B1(\u_neuron.u_td/_080_ ),
    .X(\u_neuron.u_td/_018_ ));
 sg13g2_nand3_1 \u_neuron.u_td/_157_  (.B(\u_neuron.u_td/_017_ ),
    .C(\u_neuron.u_td/_018_ ),
    .A(\u_neuron.u_td/_095_ ),
    .Y(\u_neuron.u_td/_019_ ));
 sg13g2_and4_1 \u_neuron.u_td/_158_  (.A(\u_neuron.u_td/_010_ ),
    .B(\u_neuron.u_td/_015_ ),
    .C(\u_neuron.u_td/_016_ ),
    .D(\u_neuron.u_td/_019_ ),
    .X(\u_neuron.u_td/_020_ ));
 sg13g2_nor2_1 \u_neuron.u_td/_159_  (.A(\u_neuron.u_td/_006_ ),
    .B(\u_neuron.u_td/_020_ ),
    .Y(\u_neuron.td_post_spike ));
 sg13g2_or2_1 \u_neuron.u_td/_160_  (.X(\u_neuron.td_emit_data[6] ),
    .B(\u_neuron.u_td/_020_ ),
    .A(\u_neuron.u_td/_006_ ));
 sg13g2_a21oi_1 \u_neuron.u_td/_161_  (.A1(\u_neuron.u_td/_064_ ),
    .A2(\u_neuron.u_td/_020_ ),
    .Y(\u_neuron.td_emit_valid ),
    .B1(\u_neuron.u_td/_006_ ));
 sg13g2_nand2_1 \u_neuron.u_td/_162_  (.Y(\u_neuron.u_td/_021_ ),
    .A(\u_neuron.td_curr[1] ),
    .B(\u_neuron.w_eff[1] ));
 sg13g2_nand2_1 \u_neuron.u_td/_163_  (.Y(\u_neuron.u_td/_022_ ),
    .A(\u_neuron.td_curr[0] ),
    .B(\u_neuron.w_eff[0] ));
 sg13g2_nor2_1 \u_neuron.u_td/_164_  (.A(\u_neuron.td_curr[1] ),
    .B(\u_neuron.w_eff[1] ),
    .Y(\u_neuron.u_td/_023_ ));
 sg13g2_xor2_1 \u_neuron.u_td/_165_  (.B(\u_neuron.w_eff[1] ),
    .A(\u_neuron.td_curr[1] ),
    .X(\u_neuron.u_td/_024_ ));
 sg13g2_o21ai_1 \u_neuron.u_td/_166_  (.B1(\u_neuron.u_td/_021_ ),
    .Y(\u_neuron.u_td/_025_ ),
    .A1(\u_neuron.u_td/_022_ ),
    .A2(\u_neuron.u_td/_023_ ));
 sg13g2_nand3_1 \u_neuron.u_td/_167_  (.B(\u_neuron.td_curr[2] ),
    .C(\u_neuron.u_td/_025_ ),
    .A(\u_neuron.td_curr[3] ),
    .Y(\u_neuron.u_td/_026_ ));
 sg13g2_nand4_1 \u_neuron.u_td/_168_  (.B(\u_neuron.td_curr[2] ),
    .C(\u_neuron.td_curr[4] ),
    .A(\u_neuron.td_curr[3] ),
    .Y(\u_neuron.u_td/_027_ ),
    .D(\u_neuron.u_td/_025_ ));
 sg13g2_nor2_1 \u_neuron.u_td/_169_  (.A(\u_neuron.u_td/_062_ ),
    .B(\u_neuron.u_td/_027_ ),
    .Y(\u_neuron.u_td/_028_ ));
 sg13g2_and2_1 \u_neuron.u_td/_170_  (.A(\u_neuron.td_curr[6] ),
    .B(\u_neuron.u_td/_028_ ),
    .X(\u_neuron.u_td/_029_ ));
 sg13g2_and2_1 \u_neuron.u_td/_171_  (.A(\u_neuron.td_curr[7] ),
    .B(\u_neuron.u_td/_029_ ),
    .X(\u_neuron.u_td/_030_ ));
 sg13g2_xor2_1 \u_neuron.u_td/_172_  (.B(\u_neuron.w_eff[0] ),
    .A(\u_neuron.td_curr[0] ),
    .X(\u_neuron.u_td/_031_ ));
 sg13g2_nor2b_2 \u_neuron.u_td/_173_  (.A(net382),
    .B_N(net354),
    .Y(\u_neuron.u_td/_032_ ));
 sg13g2_o21ai_1 \u_neuron.u_td/_174_  (.B1(\u_neuron.u_td/_032_ ),
    .Y(\u_neuron.u_td/_033_ ),
    .A1(\u_neuron.u_td/_030_ ),
    .A2(\u_neuron.u_td/_031_ ));
 sg13g2_o21ai_1 \u_neuron.u_td/_175_  (.B1(\u_neuron.u_td/_033_ ),
    .Y(\u_neuron.td_curr_next[0] ),
    .A1(\u_neuron.u_td/_061_ ),
    .A2(net354));
 sg13g2_xnor2_1 \u_neuron.u_td/_176_  (.Y(\u_neuron.u_td/_034_ ),
    .A(\u_neuron.u_td/_022_ ),
    .B(\u_neuron.u_td/_024_ ));
 sg13g2_o21ai_1 \u_neuron.u_td/_177_  (.B1(\u_neuron.u_td/_032_ ),
    .Y(\u_neuron.u_td/_035_ ),
    .A1(\u_neuron.u_td/_030_ ),
    .A2(\u_neuron.u_td/_034_ ));
 sg13g2_o21ai_1 \u_neuron.u_td/_178_  (.B1(\u_neuron.u_td/_035_ ),
    .Y(\u_neuron.td_curr_next[1] ),
    .A1(\u_neuron.u_td/_060_ ),
    .A2(net354));
 sg13g2_xnor2_1 \u_neuron.u_td/_179_  (.Y(\u_neuron.u_td/_036_ ),
    .A(\u_neuron.u_td/_059_ ),
    .B(\u_neuron.u_td/_025_ ));
 sg13g2_o21ai_1 \u_neuron.u_td/_180_  (.B1(\u_neuron.u_td/_032_ ),
    .Y(\u_neuron.u_td/_037_ ),
    .A1(\u_neuron.u_td/_030_ ),
    .A2(\u_neuron.u_td/_036_ ));
 sg13g2_o21ai_1 \u_neuron.u_td/_181_  (.B1(\u_neuron.u_td/_037_ ),
    .Y(\u_neuron.td_curr_next[2] ),
    .A1(\u_neuron.u_td/_059_ ),
    .A2(net354));
 sg13g2_a21o_1 \u_neuron.u_td/_182_  (.A2(\u_neuron.u_td/_025_ ),
    .A1(\u_neuron.td_curr[2] ),
    .B1(\u_neuron.td_curr[3] ),
    .X(\u_neuron.u_td/_038_ ));
 sg13g2_and2_1 \u_neuron.u_td/_183_  (.A(\u_neuron.u_td/_026_ ),
    .B(\u_neuron.u_td/_038_ ),
    .X(\u_neuron.u_td/_039_ ));
 sg13g2_o21ai_1 \u_neuron.u_td/_184_  (.B1(\u_neuron.u_td/_032_ ),
    .Y(\u_neuron.u_td/_040_ ),
    .A1(\u_neuron.u_td/_030_ ),
    .A2(\u_neuron.u_td/_039_ ));
 sg13g2_o21ai_1 \u_neuron.u_td/_185_  (.B1(\u_neuron.u_td/_040_ ),
    .Y(\u_neuron.td_curr_next[3] ),
    .A1(\u_neuron.u_td/_058_ ),
    .A2(net354));
 sg13g2_xnor2_1 \u_neuron.u_td/_186_  (.Y(\u_neuron.u_td/_041_ ),
    .A(\u_neuron.td_curr[4] ),
    .B(\u_neuron.u_td/_026_ ));
 sg13g2_o21ai_1 \u_neuron.u_td/_187_  (.B1(\u_neuron.u_td/_032_ ),
    .Y(\u_neuron.u_td/_042_ ),
    .A1(\u_neuron.u_td/_030_ ),
    .A2(\u_neuron.u_td/_041_ ));
 sg13g2_o21ai_1 \u_neuron.u_td/_188_  (.B1(\u_neuron.u_td/_042_ ),
    .Y(\u_neuron.td_curr_next[4] ),
    .A1(\u_neuron.u_td/_063_ ),
    .A2(net354));
 sg13g2_xnor2_1 \u_neuron.u_td/_189_  (.Y(\u_neuron.u_td/_043_ ),
    .A(\u_neuron.td_curr[5] ),
    .B(\u_neuron.u_td/_027_ ));
 sg13g2_o21ai_1 \u_neuron.u_td/_190_  (.B1(\u_neuron.u_td/_032_ ),
    .Y(\u_neuron.u_td/_044_ ),
    .A1(\u_neuron.u_td/_030_ ),
    .A2(\u_neuron.u_td/_043_ ));
 sg13g2_o21ai_1 \u_neuron.u_td/_191_  (.B1(\u_neuron.u_td/_044_ ),
    .Y(\u_neuron.td_curr_next[5] ),
    .A1(\u_neuron.u_td/_062_ ),
    .A2(net354));
 sg13g2_nand2b_1 \u_neuron.u_td/_192_  (.Y(\u_neuron.u_td/_045_ ),
    .B(net155),
    .A_N(net354));
 sg13g2_nor2b_1 \u_neuron.u_td/_193_  (.A(net153),
    .B_N(\u_neuron.u_td/_029_ ),
    .Y(\u_neuron.u_td/_046_ ));
 sg13g2_o21ai_1 \u_neuron.u_td/_194_  (.B1(\u_neuron.u_td/_032_ ),
    .Y(\u_neuron.u_td/_047_ ),
    .A1(net155),
    .A2(\u_neuron.u_td/_028_ ));
 sg13g2_o21ai_1 \u_neuron.u_td/_195_  (.B1(\u_neuron.u_td/_045_ ),
    .Y(\u_neuron.td_curr_next[6] ),
    .A1(\u_neuron.u_td/_046_ ),
    .A2(\u_neuron.u_td/_047_ ));
 sg13g2_a21oi_1 \u_neuron.u_td/_196_  (.A1(net355),
    .A2(\u_neuron.u_td/_029_ ),
    .Y(\u_neuron.u_td/_048_ ),
    .B1(net153));
 sg13g2_a21oi_1 \u_neuron.u_td/_197_  (.A1(net382),
    .A2(net355),
    .Y(\u_neuron.td_curr_next[7] ),
    .B1(\u_neuron.u_td/_048_ ));
 sg13g2_nand2_1 \u_neuron.u_td/_198_  (.Y(\u_neuron.u_td/_049_ ),
    .A(net126),
    .B(net327));
 sg13g2_o21ai_1 \u_neuron.u_td/_199_  (.B1(\u_neuron.u_td/_049_ ),
    .Y(\u_neuron.td_prev_next[0] ),
    .A1(\u_neuron.u_td/_061_ ),
    .A2(net327));
 sg13g2_nand2_1 \u_neuron.u_td/_200_  (.Y(\u_neuron.u_td/_050_ ),
    .A(net114),
    .B(net326));
 sg13g2_o21ai_1 \u_neuron.u_td/_201_  (.B1(\u_neuron.u_td/_050_ ),
    .Y(\u_neuron.td_prev_next[1] ),
    .A1(\u_neuron.u_td/_060_ ),
    .A2(net326));
 sg13g2_nand2_1 \u_neuron.u_td/_202_  (.Y(\u_neuron.u_td/_051_ ),
    .A(net118),
    .B(net326));
 sg13g2_o21ai_1 \u_neuron.u_td/_203_  (.B1(\u_neuron.u_td/_051_ ),
    .Y(\u_neuron.td_prev_next[2] ),
    .A1(\u_neuron.u_td/_059_ ),
    .A2(net326));
 sg13g2_nand2_1 \u_neuron.u_td/_204_  (.Y(\u_neuron.u_td/_052_ ),
    .A(net140),
    .B(net327));
 sg13g2_o21ai_1 \u_neuron.u_td/_205_  (.B1(\u_neuron.u_td/_052_ ),
    .Y(\u_neuron.td_prev_next[3] ),
    .A1(\u_neuron.u_td/_058_ ),
    .A2(net327));
 sg13g2_nand2_1 \u_neuron.u_td/_206_  (.Y(\u_neuron.u_td/_053_ ),
    .A(net151),
    .B(net326));
 sg13g2_o21ai_1 \u_neuron.u_td/_207_  (.B1(\u_neuron.u_td/_053_ ),
    .Y(\u_neuron.td_prev_next[4] ),
    .A1(\u_neuron.u_td/_063_ ),
    .A2(net326));
 sg13g2_nand2_1 \u_neuron.u_td/_208_  (.Y(\u_neuron.u_td/_054_ ),
    .A(net144),
    .B(net326));
 sg13g2_o21ai_1 \u_neuron.u_td/_209_  (.B1(\u_neuron.u_td/_054_ ),
    .Y(\u_neuron.td_prev_next[5] ),
    .A1(\u_neuron.u_td/_062_ ),
    .A2(net326));
 sg13g2_mux2_1 \u_neuron.u_td/_210_  (.A0(\u_neuron.td_curr[6] ),
    .A1(net112),
    .S(net329),
    .X(\u_neuron.td_prev_next[6] ));
 sg13g2_mux2_1 \u_neuron.u_td/_211_  (.A0(\u_neuron.td_curr[7] ),
    .A1(net131),
    .S(net327),
    .X(\u_neuron.td_prev_next[7] ));
 sg13g2_mux2_1 \u_neuron.u_td/_212_  (.A0(\u_neuron.td_emit_data[0] ),
    .A1(net68),
    .S(net328),
    .X(\u_neuron.td_last_diff_next[0] ));
 sg13g2_mux2_1 \u_neuron.u_td/_213_  (.A0(\u_neuron.td_emit_data[1] ),
    .A1(net75),
    .S(net328),
    .X(\u_neuron.td_last_diff_next[1] ));
 sg13g2_mux2_1 \u_neuron.u_td/_214_  (.A0(\u_neuron.td_emit_data[2] ),
    .A1(net84),
    .S(net329),
    .X(\u_neuron.td_last_diff_next[2] ));
 sg13g2_mux2_1 \u_neuron.u_td/_215_  (.A0(\u_neuron.td_emit_data[3] ),
    .A1(net79),
    .S(net329),
    .X(\u_neuron.td_last_diff_next[3] ));
 sg13g2_mux2_1 \u_neuron.u_td/_216_  (.A0(\u_neuron.u_td/_009_ ),
    .A1(net61),
    .S(net328),
    .X(\u_neuron.td_last_diff_next[4] ));
 sg13g2_nand2_1 \u_neuron.u_td/_217_  (.Y(\u_neuron.u_td/_055_ ),
    .A(net80),
    .B(net327));
 sg13g2_o21ai_1 \u_neuron.u_td/_218_  (.B1(\u_neuron.u_td/_055_ ),
    .Y(\u_neuron.td_last_diff_next[5] ),
    .A1(net327),
    .A2(\u_neuron.u_td/_019_ ));
 sg13g2_nand2_1 \u_neuron.u_td/_219_  (.Y(\u_neuron.u_td/_056_ ),
    .A(net87),
    .B(net328));
 sg13g2_o21ai_1 \u_neuron.u_td/_220_  (.B1(\u_neuron.u_td/_056_ ),
    .Y(\u_neuron.td_last_diff_next[6] ),
    .A1(net328),
    .A2(\u_neuron.u_td/_015_ ));
 sg13g2_nand2_1 \u_neuron.u_td/_221_  (.Y(\u_neuron.u_td/_057_ ),
    .A(net64),
    .B(net328));
 sg13g2_o21ai_1 \u_neuron.u_td/_222_  (.B1(\u_neuron.u_td/_057_ ),
    .Y(\u_neuron.td_last_diff_next[7] ),
    .A1(net328),
    .A2(\u_neuron.u_td/_016_ ));
 sg13g2_buf_8 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_tielo \u_neuron.u_mode_sel/_00__36  (.L_LO(net36));
 sg13g2_tiehi \u_neuron.u_mode_sel/_09__37  (.L_HI(net37));
 sg13g2_buf_1 \u_neuron.u_td/_226_  (.A(\u_neuron.td_emit_data[6] ),
    .X(\u_neuron.td_emit_data[4] ));
 sg13g2_buf_8 fanout314 (.A(\u_neuron.u_outq/_20_ ),
    .X(net314));
 sg13g2_buf_8 fanout315 (.A(\u_neuron.u_syn/_045_ ),
    .X(net315));
 sg13g2_buf_8 fanout316 (.A(net318),
    .X(net316));
 sg13g2_buf_2 fanout317 (.A(net318),
    .X(net317));
 sg13g2_buf_8 fanout318 (.A(\u_neuron.u_syn/_312_ ),
    .X(net318));
 sg13g2_buf_8 fanout319 (.A(net320),
    .X(net319));
 sg13g2_buf_8 fanout320 (.A(\u_neuron.u_syn/_160_ ),
    .X(net320));
 sg13g2_buf_8 fanout321 (.A(\u_neuron.ltp_we ),
    .X(net321));
 sg13g2_buf_8 fanout322 (.A(\u_neuron.u_fst/_019_ ),
    .X(net322));
 sg13g2_buf_8 fanout323 (.A(\u_neuron.u_fst/_019_ ),
    .X(net323));
 sg13g2_buf_8 fanout324 (.A(\u_neuron.u_conv/_03_ ),
    .X(net324));
 sg13g2_buf_1 fanout325 (.A(\u_neuron.u_conv/_03_ ),
    .X(net325));
 sg13g2_buf_8 fanout326 (.A(net327),
    .X(net326));
 sg13g2_buf_8 fanout327 (.A(net329),
    .X(net327));
 sg13g2_buf_8 fanout328 (.A(net329),
    .X(net328));
 sg13g2_buf_8 fanout329 (.A(\u_neuron.u_td/_005_ ),
    .X(net329));
 sg13g2_buf_8 fanout330 (.A(\u_neuron.u_learning/_027_ ),
    .X(net330));
 sg13g2_buf_8 fanout331 (.A(\u_neuron.ltd_wdata[1] ),
    .X(net331));
 sg13g2_buf_8 fanout332 (.A(\u_neuron.ltd_wdata[0] ),
    .X(net332));
 sg13g2_buf_8 fanout333 (.A(\u_neuron.ltp_wdata[1] ),
    .X(net333));
 sg13g2_buf_8 fanout334 (.A(net336),
    .X(net334));
 sg13g2_buf_1 fanout335 (.A(net336),
    .X(net335));
 sg13g2_buf_8 fanout336 (.A(net352),
    .X(net336));
 sg13g2_buf_8 fanout337 (.A(net339),
    .X(net337));
 sg13g2_buf_1 fanout338 (.A(net339),
    .X(net338));
 sg13g2_buf_8 fanout339 (.A(net352),
    .X(net339));
 sg13g2_buf_8 fanout340 (.A(net343),
    .X(net340));
 sg13g2_buf_1 fanout341 (.A(net343),
    .X(net341));
 sg13g2_buf_8 fanout342 (.A(net343),
    .X(net342));
 sg13g2_buf_8 fanout343 (.A(net352),
    .X(net343));
 sg13g2_buf_8 fanout344 (.A(net345),
    .X(net344));
 sg13g2_buf_8 fanout345 (.A(net346),
    .X(net345));
 sg13g2_buf_8 fanout346 (.A(net352),
    .X(net346));
 sg13g2_buf_8 fanout347 (.A(net350),
    .X(net347));
 sg13g2_buf_8 fanout348 (.A(net350),
    .X(net348));
 sg13g2_buf_2 fanout349 (.A(net350),
    .X(net349));
 sg13g2_buf_8 fanout350 (.A(net351),
    .X(net350));
 sg13g2_buf_2 fanout351 (.A(net352),
    .X(net351));
 sg13g2_buf_8 fanout352 (.A(_129_),
    .X(net352));
 sg13g2_buf_8 fanout353 (.A(\u_neuron.mode_lif_evt ),
    .X(net353));
 sg13g2_buf_8 fanout354 (.A(net355),
    .X(net354));
 sg13g2_buf_2 fanout355 (.A(\u_neuron.mode_td_evt ),
    .X(net355));
 sg13g2_buf_8 fanout356 (.A(\u_neuron.normal_event ),
    .X(net356));
 sg13g2_buf_2 fanout357 (.A(net360),
    .X(net357));
 sg13g2_buf_1 fanout358 (.A(net360),
    .X(net358));
 sg13g2_buf_8 fanout359 (.A(net360),
    .X(net359));
 sg13g2_buf_8 fanout360 (.A(_001_),
    .X(net360));
 sg13g2_buf_8 fanout361 (.A(net362),
    .X(net361));
 sg13g2_buf_2 fanout362 (.A(net363),
    .X(net362));
 sg13g2_buf_8 fanout363 (.A(\u_neuron.u_learning/_118_ ),
    .X(net363));
 sg13g2_buf_8 fanout364 (.A(net366),
    .X(net364));
 sg13g2_buf_1 fanout365 (.A(net366),
    .X(net365));
 sg13g2_buf_8 fanout366 (.A(\u_neuron.u_learning/_025_ ),
    .X(net366));
 sg13g2_buf_8 fanout367 (.A(\u_neuron.ltd_idx[2] ),
    .X(net367));
 sg13g2_buf_1 fanout368 (.A(\u_neuron.ltd_idx[2] ),
    .X(net368));
 sg13g2_buf_2 fanout369 (.A(net370),
    .X(net369));
 sg13g2_buf_8 fanout370 (.A(net371),
    .X(net370));
 sg13g2_buf_2 fanout371 (.A(net379),
    .X(net371));
 sg13g2_buf_2 fanout372 (.A(net373),
    .X(net372));
 sg13g2_buf_1 fanout373 (.A(net379),
    .X(net373));
 sg13g2_buf_2 fanout374 (.A(net375),
    .X(net374));
 sg13g2_buf_1 fanout375 (.A(net379),
    .X(net375));
 sg13g2_buf_1 fanout376 (.A(net377),
    .X(net376));
 sg13g2_buf_8 fanout377 (.A(net378),
    .X(net377));
 sg13g2_buf_1 fanout378 (.A(net379),
    .X(net378));
 sg13g2_buf_2 fanout379 (.A(\u_neuron.is_reset_cmd ),
    .X(net379));
 sg13g2_buf_8 fanout380 (.A(\u_neuron.u_learning/_119_ ),
    .X(net380));
 sg13g2_buf_1 fanout381 (.A(\u_neuron.u_learning/_119_ ),
    .X(net381));
 sg13g2_buf_8 fanout382 (.A(net384),
    .X(net382));
 sg13g2_buf_1 fanout383 (.A(net384),
    .X(net383));
 sg13g2_buf_8 fanout384 (.A(\u_neuron.is_tick ),
    .X(net384));
 sg13g2_buf_8 fanout385 (.A(\u_neuron.is_tick ),
    .X(net385));
 sg13g2_buf_8 fanout386 (.A(net387),
    .X(net386));
 sg13g2_buf_8 fanout387 (.A(\u_neuron.addr[3] ),
    .X(net387));
 sg13g2_buf_8 fanout388 (.A(net390),
    .X(net388));
 sg13g2_buf_1 fanout389 (.A(net390),
    .X(net389));
 sg13g2_buf_8 fanout390 (.A(\u_neuron.addr[2] ),
    .X(net390));
 sg13g2_buf_8 fanout391 (.A(net393),
    .X(net391));
 sg13g2_buf_1 fanout392 (.A(net393),
    .X(net392));
 sg13g2_buf_8 fanout393 (.A(net395),
    .X(net393));
 sg13g2_buf_8 fanout394 (.A(net395),
    .X(net394));
 sg13g2_buf_8 fanout395 (.A(\u_neuron.addr[1] ),
    .X(net395));
 sg13g2_buf_8 fanout396 (.A(net398),
    .X(net396));
 sg13g2_buf_1 fanout397 (.A(net398),
    .X(net397));
 sg13g2_buf_8 fanout398 (.A(net399),
    .X(net398));
 sg13g2_buf_8 fanout399 (.A(\u_neuron.addr[0] ),
    .X(net399));
 sg13g2_buf_8 fanout400 (.A(net401),
    .X(net400));
 sg13g2_buf_1 fanout401 (.A(\u_neuron.addr[0] ),
    .X(net401));
 sg13g2_buf_8 fanout402 (.A(net403),
    .X(net402));
 sg13g2_buf_8 fanout403 (.A(\u_neuron.addr[0] ),
    .X(net403));
 sg13g2_buf_8 fanout404 (.A(net405),
    .X(net404));
 sg13g2_buf_2 fanout405 (.A(net406),
    .X(net405));
 sg13g2_buf_1 fanout406 (.A(net407),
    .X(net406));
 sg13g2_buf_8 fanout407 (.A(\u_neuron.pending_widx[2] ),
    .X(net407));
 sg13g2_buf_8 fanout408 (.A(\u_neuron.pending_widx[1] ),
    .X(net408));
 sg13g2_buf_8 fanout409 (.A(net226),
    .X(net409));
 sg13g2_buf_8 fanout410 (.A(net411),
    .X(net410));
 sg13g2_buf_8 fanout411 (.A(net414),
    .X(net411));
 sg13g2_buf_8 fanout412 (.A(net413),
    .X(net412));
 sg13g2_buf_8 fanout413 (.A(net414),
    .X(net413));
 sg13g2_buf_8 fanout414 (.A(\u_neuron.u_syn/_036_ ),
    .X(net414));
 sg13g2_buf_8 fanout415 (.A(net416),
    .X(net415));
 sg13g2_buf_8 fanout416 (.A(\u_neuron.u_syn/_036_ ),
    .X(net416));
 sg13g2_buf_8 fanout417 (.A(\u_neuron.have_out ),
    .X(net417));
 sg13g2_buf_1 fanout418 (.A(net233),
    .X(net418));
 sg13g2_buf_8 fanout419 (.A(net224),
    .X(net419));
 sg13g2_buf_2 fanout420 (.A(\u_neuron.learn_ptr[3] ),
    .X(net420));
 sg13g2_buf_8 fanout421 (.A(net422),
    .X(net421));
 sg13g2_buf_1 fanout422 (.A(net423),
    .X(net422));
 sg13g2_buf_8 fanout423 (.A(\u_neuron.learn_ptr[2] ),
    .X(net423));
 sg13g2_buf_8 fanout424 (.A(net425),
    .X(net424));
 sg13g2_buf_2 fanout425 (.A(net426),
    .X(net425));
 sg13g2_buf_8 fanout426 (.A(\u_neuron.learn_ptr[1] ),
    .X(net426));
 sg13g2_buf_8 fanout427 (.A(net428),
    .X(net427));
 sg13g2_buf_8 fanout428 (.A(net218),
    .X(net428));
 sg13g2_buf_8 fanout429 (.A(net430),
    .X(net429));
 sg13g2_buf_8 fanout430 (.A(\u_neuron.learn_ptr[0] ),
    .X(net430));
 sg13g2_buf_8 fanout431 (.A(net432),
    .X(net431));
 sg13g2_buf_8 fanout432 (.A(net231),
    .X(net432));
 sg13g2_buf_8 fanout433 (.A(net434),
    .X(net433));
 sg13g2_buf_8 fanout434 (.A(\u_neuron.mode[0] ),
    .X(net434));
 sg13g2_buf_8 fanout435 (.A(\u_neuron.fst_t[0] ),
    .X(net435));
 sg13g2_buf_8 fanout436 (.A(net448),
    .X(net436));
 sg13g2_buf_8 fanout437 (.A(net448),
    .X(net437));
 sg13g2_buf_8 fanout438 (.A(net440),
    .X(net438));
 sg13g2_buf_2 fanout439 (.A(net440),
    .X(net439));
 sg13g2_buf_8 fanout440 (.A(net448),
    .X(net440));
 sg13g2_buf_8 fanout441 (.A(net444),
    .X(net441));
 sg13g2_buf_8 fanout442 (.A(net443),
    .X(net442));
 sg13g2_buf_8 fanout443 (.A(net444),
    .X(net443));
 sg13g2_buf_8 fanout444 (.A(net447),
    .X(net444));
 sg13g2_buf_8 fanout445 (.A(net446),
    .X(net445));
 sg13g2_buf_8 fanout446 (.A(net447),
    .X(net446));
 sg13g2_buf_8 fanout447 (.A(net448),
    .X(net447));
 sg13g2_buf_8 fanout448 (.A(rst_n),
    .X(net448));
 sg13g2_buf_8 fanout449 (.A(net450),
    .X(net449));
 sg13g2_buf_8 fanout450 (.A(net455),
    .X(net450));
 sg13g2_buf_8 fanout451 (.A(net455),
    .X(net451));
 sg13g2_buf_8 fanout452 (.A(net455),
    .X(net452));
 sg13g2_buf_8 fanout453 (.A(net454),
    .X(net453));
 sg13g2_buf_8 fanout454 (.A(net455),
    .X(net454));
 sg13g2_buf_8 fanout455 (.A(rst_n),
    .X(net455));
 sg13g2_buf_8 fanout456 (.A(net464),
    .X(net456));
 sg13g2_buf_8 fanout457 (.A(net464),
    .X(net457));
 sg13g2_buf_8 fanout458 (.A(net460),
    .X(net458));
 sg13g2_buf_8 fanout459 (.A(net460),
    .X(net459));
 sg13g2_buf_8 fanout460 (.A(net464),
    .X(net460));
 sg13g2_buf_8 fanout461 (.A(net462),
    .X(net461));
 sg13g2_buf_8 fanout462 (.A(net463),
    .X(net462));
 sg13g2_buf_2 fanout463 (.A(net464),
    .X(net463));
 sg13g2_buf_8 fanout464 (.A(rst_n),
    .X(net464));
 sg13g2_buf_8 fanout465 (.A(ena),
    .X(net465));
 sg13g2_buf_1 fanout466 (.A(ena),
    .X(net466));
 sg13g2_buf_8 fanout467 (.A(net468),
    .X(net467));
 sg13g2_buf_8 fanout468 (.A(net469),
    .X(net468));
 sg13g2_buf_8 fanout469 (.A(ena),
    .X(net469));
 sg13g2_buf_1 input1 (.A(ui_in[0]),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[1]),
    .X(net2));
 sg13g2_buf_1 input3 (.A(ui_in[2]),
    .X(net3));
 sg13g2_buf_1 input4 (.A(ui_in[3]),
    .X(net4));
 sg13g2_buf_1 input5 (.A(ui_in[4]),
    .X(net5));
 sg13g2_buf_1 input6 (.A(ui_in[5]),
    .X(net6));
 sg13g2_buf_1 input7 (.A(ui_in[6]),
    .X(net7));
 sg13g2_buf_1 input8 (.A(ui_in[7]),
    .X(net8));
 sg13g2_buf_1 input9 (.A(uio_in[0]),
    .X(net9));
 sg13g2_buf_1 input10 (.A(uio_in[1]),
    .X(net10));
 sg13g2_buf_1 input11 (.A(uio_in[2]),
    .X(net11));
 sg13g2_buf_1 input12 (.A(uio_in[3]),
    .X(net12));
 sg13g2_buf_1 input13 (.A(uio_in[4]),
    .X(net13));
 sg13g2_buf_1 input14 (.A(uio_in[5]),
    .X(net14));
 sg13g2_buf_1 input15 (.A(uio_in[6]),
    .X(net15));
 sg13g2_buf_1 input16 (.A(uio_in[7]),
    .X(net16));
 sg13g2_tielo \u_neuron.u_mode_sel/_05__17  (.L_LO(net17));
 sg13g2_buf_8 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sg13g2_buf_8 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sg13g2_buf_8 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sg13g2_buf_8 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sg13g2_buf_8 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sg13g2_buf_8 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sg13g2_buf_8 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sg13g2_buf_8 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sg13g2_buf_8 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sg13g2_buf_8 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sg13g2_buf_8 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sg13g2_buf_8 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sg13g2_buf_8 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sg13g2_buf_8 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sg13g2_buf_8 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sg13g2_buf_8 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sg13g2_buf_8 clkbuf_5_0__f_clk (.A(clknet_4_0_0_clk),
    .X(clknet_5_0__leaf_clk));
 sg13g2_buf_8 clkbuf_5_1__f_clk (.A(clknet_4_0_0_clk),
    .X(clknet_5_1__leaf_clk));
 sg13g2_buf_8 clkbuf_5_2__f_clk (.A(clknet_4_1_0_clk),
    .X(clknet_5_2__leaf_clk));
 sg13g2_buf_8 clkbuf_5_3__f_clk (.A(clknet_4_1_0_clk),
    .X(clknet_5_3__leaf_clk));
 sg13g2_buf_8 clkbuf_5_4__f_clk (.A(clknet_4_2_0_clk),
    .X(clknet_5_4__leaf_clk));
 sg13g2_buf_8 clkbuf_5_5__f_clk (.A(clknet_4_2_0_clk),
    .X(clknet_5_5__leaf_clk));
 sg13g2_buf_8 clkbuf_5_6__f_clk (.A(clknet_4_3_0_clk),
    .X(clknet_5_6__leaf_clk));
 sg13g2_buf_8 clkbuf_5_7__f_clk (.A(clknet_4_3_0_clk),
    .X(clknet_5_7__leaf_clk));
 sg13g2_buf_8 clkbuf_5_8__f_clk (.A(clknet_4_4_0_clk),
    .X(clknet_5_8__leaf_clk));
 sg13g2_buf_8 clkbuf_5_9__f_clk (.A(clknet_4_4_0_clk),
    .X(clknet_5_9__leaf_clk));
 sg13g2_buf_8 clkbuf_5_10__f_clk (.A(clknet_4_5_0_clk),
    .X(clknet_5_10__leaf_clk));
 sg13g2_buf_8 clkbuf_5_11__f_clk (.A(clknet_4_5_0_clk),
    .X(clknet_5_11__leaf_clk));
 sg13g2_buf_8 clkbuf_5_12__f_clk (.A(clknet_4_6_0_clk),
    .X(clknet_5_12__leaf_clk));
 sg13g2_buf_8 clkbuf_5_13__f_clk (.A(clknet_4_6_0_clk),
    .X(clknet_5_13__leaf_clk));
 sg13g2_buf_8 clkbuf_5_14__f_clk (.A(clknet_4_7_0_clk),
    .X(clknet_5_14__leaf_clk));
 sg13g2_buf_8 clkbuf_5_15__f_clk (.A(clknet_4_7_0_clk),
    .X(clknet_5_15__leaf_clk));
 sg13g2_buf_8 clkbuf_5_16__f_clk (.A(clknet_4_8_0_clk),
    .X(clknet_5_16__leaf_clk));
 sg13g2_buf_8 clkbuf_5_17__f_clk (.A(clknet_4_8_0_clk),
    .X(clknet_5_17__leaf_clk));
 sg13g2_buf_8 clkbuf_5_18__f_clk (.A(clknet_4_9_0_clk),
    .X(clknet_5_18__leaf_clk));
 sg13g2_buf_8 clkbuf_5_19__f_clk (.A(clknet_4_9_0_clk),
    .X(clknet_5_19__leaf_clk));
 sg13g2_buf_8 clkbuf_5_20__f_clk (.A(clknet_4_10_0_clk),
    .X(clknet_5_20__leaf_clk));
 sg13g2_buf_8 clkbuf_5_21__f_clk (.A(clknet_4_10_0_clk),
    .X(clknet_5_21__leaf_clk));
 sg13g2_buf_8 clkbuf_5_22__f_clk (.A(clknet_4_11_0_clk),
    .X(clknet_5_22__leaf_clk));
 sg13g2_buf_8 clkbuf_5_23__f_clk (.A(clknet_4_11_0_clk),
    .X(clknet_5_23__leaf_clk));
 sg13g2_buf_8 clkbuf_5_24__f_clk (.A(clknet_4_12_0_clk),
    .X(clknet_5_24__leaf_clk));
 sg13g2_buf_8 clkbuf_5_25__f_clk (.A(clknet_4_12_0_clk),
    .X(clknet_5_25__leaf_clk));
 sg13g2_buf_8 clkbuf_5_26__f_clk (.A(clknet_4_13_0_clk),
    .X(clknet_5_26__leaf_clk));
 sg13g2_buf_8 clkbuf_5_27__f_clk (.A(clknet_4_13_0_clk),
    .X(clknet_5_27__leaf_clk));
 sg13g2_buf_8 clkbuf_5_28__f_clk (.A(clknet_4_14_0_clk),
    .X(clknet_5_28__leaf_clk));
 sg13g2_buf_8 clkbuf_5_29__f_clk (.A(clknet_4_14_0_clk),
    .X(clknet_5_29__leaf_clk));
 sg13g2_buf_8 clkbuf_5_30__f_clk (.A(clknet_4_15_0_clk),
    .X(clknet_5_30__leaf_clk));
 sg13g2_buf_8 clkbuf_5_31__f_clk (.A(clknet_4_15_0_clk),
    .X(clknet_5_31__leaf_clk));
 sg13g2_inv_1 clkload0 (.A(clknet_5_1__leaf_clk));
 sg13g2_buf_1 clkload1 (.A(clknet_5_3__leaf_clk));
 sg13g2_buf_1 clkload2 (.A(clknet_5_4__leaf_clk));
 sg13g2_buf_1 clkload3 (.A(clknet_5_7__leaf_clk));
 sg13g2_buf_1 clkload4 (.A(clknet_5_8__leaf_clk));
 sg13g2_buf_1 clkload5 (.A(clknet_5_14__leaf_clk));
 sg13g2_buf_1 clkload6 (.A(clknet_5_16__leaf_clk));
 sg13g2_buf_1 clkload7 (.A(clknet_5_19__leaf_clk));
 sg13g2_buf_1 clkload8 (.A(clknet_5_27__leaf_clk));
 sg13g2_buf_1 clkload9 (.A(clknet_5_29__leaf_clk));
 sg13g2_buf_1 clkload10 (.A(clknet_5_31__leaf_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(\u_neuron.u_frontend/uio_in_meta[6] ),
    .X(net43));
 sg13g2_dlygate4sd3_1 hold2 (.A(\u_neuron.u_frontend/uio_in_meta[7] ),
    .X(net44));
 sg13g2_dlygate4sd3_1 hold3 (.A(\u_neuron.u_frontend/uio_in_meta[5] ),
    .X(net45));
 sg13g2_dlygate4sd3_1 hold4 (.A(\u_neuron.u_frontend/ui_in_meta[2] ),
    .X(net46));
 sg13g2_dlygate4sd3_1 hold5 (.A(\u_neuron.u_frontend/uio_in_meta[2] ),
    .X(net47));
 sg13g2_dlygate4sd3_1 hold6 (.A(\u_neuron.u_frontend/ui_in_meta[6] ),
    .X(net48));
 sg13g2_dlygate4sd3_1 hold7 (.A(\u_neuron.u_frontend/ui_in_meta[3] ),
    .X(net49));
 sg13g2_dlygate4sd3_1 hold8 (.A(\u_neuron.u_frontend/uio_in_meta[3] ),
    .X(net50));
 sg13g2_dlygate4sd3_1 hold9 (.A(\u_neuron.u_frontend/ui_in_meta[4] ),
    .X(net51));
 sg13g2_dlygate4sd3_1 hold10 (.A(\u_neuron.u_frontend/ui_in_meta[5] ),
    .X(net52));
 sg13g2_dlygate4sd3_1 hold11 (.A(\u_neuron.u_frontend/ui_in_meta[0] ),
    .X(net53));
 sg13g2_dlygate4sd3_1 hold12 (.A(\u_neuron.u_frontend/ui_in_meta[1] ),
    .X(net54));
 sg13g2_dlygate4sd3_1 hold13 (.A(\u_neuron.u_frontend/ui_in_meta[7] ),
    .X(net55));
 sg13g2_dlygate4sd3_1 hold14 (.A(\u_neuron.u_frontend/uio_in_meta[0] ),
    .X(net56));
 sg13g2_dlygate4sd3_1 hold15 (.A(\u_neuron.u_frontend/uio_in_meta[1] ),
    .X(net57));
 sg13g2_dlygate4sd3_1 hold16 (.A(\u_neuron.u_frontend/uio_in_meta[4] ),
    .X(net58));
 sg13g2_dlygate4sd3_1 hold17 (.A(\u_neuron.fst_last_t[0] ),
    .X(net59));
 sg13g2_dlygate4sd3_1 hold18 (.A(_030_),
    .X(net60));
 sg13g2_dlygate4sd3_1 hold19 (.A(\u_neuron.td_last_diff[4] ),
    .X(net61));
 sg13g2_dlygate4sd3_1 hold20 (.A(\u_neuron.fst_last_t[4] ),
    .X(net62));
 sg13g2_dlygate4sd3_1 hold21 (.A(_034_),
    .X(net63));
 sg13g2_dlygate4sd3_1 hold22 (.A(\u_neuron.td_last_diff[7] ),
    .X(net64));
 sg13g2_dlygate4sd3_1 hold23 (.A(_013_),
    .X(net65));
 sg13g2_dlygate4sd3_1 hold24 (.A(\u_neuron.fst_last_t[5] ),
    .X(net66));
 sg13g2_dlygate4sd3_1 hold25 (.A(_035_),
    .X(net67));
 sg13g2_dlygate4sd3_1 hold26 (.A(\u_neuron.td_last_diff[0] ),
    .X(net68));
 sg13g2_dlygate4sd3_1 hold27 (.A(\u_neuron.in_req_seen ),
    .X(net69));
 sg13g2_dlygate4sd3_1 hold28 (.A(\u_neuron.u_frontend/_03_ ),
    .X(net70));
 sg13g2_dlygate4sd3_1 hold29 (.A(\u_neuron.u_frontend/_00_ ),
    .X(net71));
 sg13g2_dlygate4sd3_1 hold30 (.A(\u_neuron.conv_last_sum[2] ),
    .X(net72));
 sg13g2_dlygate4sd3_1 hold31 (.A(\u_neuron.fst_last_t[6] ),
    .X(net73));
 sg13g2_dlygate4sd3_1 hold32 (.A(_036_),
    .X(net74));
 sg13g2_dlygate4sd3_1 hold33 (.A(\u_neuron.td_last_diff[1] ),
    .X(net75));
 sg13g2_dlygate4sd3_1 hold34 (.A(\u_neuron.conv_last_sum[0] ),
    .X(net76));
 sg13g2_dlygate4sd3_1 hold35 (.A(\u_neuron.conv_shift[3] ),
    .X(net77));
 sg13g2_dlygate4sd3_1 hold36 (.A(_058_),
    .X(net78));
 sg13g2_dlygate4sd3_1 hold37 (.A(\u_neuron.td_last_diff[3] ),
    .X(net79));
 sg13g2_dlygate4sd3_1 hold38 (.A(\u_neuron.td_last_diff[5] ),
    .X(net80));
 sg13g2_dlygate4sd3_1 hold39 (.A(\u_neuron.fst_last_t[7] ),
    .X(net81));
 sg13g2_dlygate4sd3_1 hold40 (.A(_037_),
    .X(net82));
 sg13g2_dlygate4sd3_1 hold41 (.A(\u_neuron.conv_last_sum[1] ),
    .X(net83));
 sg13g2_dlygate4sd3_1 hold42 (.A(\u_neuron.td_last_diff[2] ),
    .X(net84));
 sg13g2_dlygate4sd3_1 hold43 (.A(\u_neuron.pre_trace[0] ),
    .X(net85));
 sg13g2_dlygate4sd3_1 hold44 (.A(\u_neuron.u_learning/_034_ ),
    .X(net86));
 sg13g2_dlygate4sd3_1 hold45 (.A(\u_neuron.td_last_diff[6] ),
    .X(net87));
 sg13g2_dlygate4sd3_1 hold46 (.A(\u_neuron.fst_last_t[3] ),
    .X(net88));
 sg13g2_dlygate4sd3_1 hold47 (.A(_033_),
    .X(net89));
 sg13g2_dlygate4sd3_1 hold48 (.A(\u_neuron.pre_trace[2] ),
    .X(net90));
 sg13g2_dlygate4sd3_1 hold49 (.A(\u_neuron.pre_trace[1] ),
    .X(net91));
 sg13g2_dlygate4sd3_1 hold50 (.A(\u_neuron.pre_trace[9] ),
    .X(net92));
 sg13g2_dlygate4sd3_1 hold51 (.A(\u_neuron.pre_trace[12] ),
    .X(net93));
 sg13g2_dlygate4sd3_1 hold52 (.A(\u_neuron.pre_trace[3] ),
    .X(net94));
 sg13g2_dlygate4sd3_1 hold53 (.A(\u_neuron.pre_trace[13] ),
    .X(net95));
 sg13g2_dlygate4sd3_1 hold54 (.A(\u_neuron.pre_trace[7] ),
    .X(net96));
 sg13g2_dlygate4sd3_1 hold55 (.A(\u_neuron.u_learning/_007_ ),
    .X(net97));
 sg13g2_dlygate4sd3_1 hold56 (.A(\u_neuron.conv_shift[2] ),
    .X(net98));
 sg13g2_dlygate4sd3_1 hold57 (.A(_057_),
    .X(net99));
 sg13g2_dlygate4sd3_1 hold58 (.A(\u_neuron.pre_trace[10] ),
    .X(net100));
 sg13g2_dlygate4sd3_1 hold59 (.A(\u_neuron.pre_trace[4] ),
    .X(net101));
 sg13g2_dlygate4sd3_1 hold60 (.A(\u_neuron.pre_trace[6] ),
    .X(net102));
 sg13g2_dlygate4sd3_1 hold61 (.A(\u_neuron.pre_trace[14] ),
    .X(net103));
 sg13g2_dlygate4sd3_1 hold62 (.A(\u_neuron.fst_last_t[2] ),
    .X(net104));
 sg13g2_dlygate4sd3_1 hold63 (.A(_032_),
    .X(net105));
 sg13g2_dlygate4sd3_1 hold64 (.A(\u_neuron.pre_trace[5] ),
    .X(net106));
 sg13g2_dlygate4sd3_1 hold65 (.A(\u_neuron.pre_trace[8] ),
    .X(net107));
 sg13g2_dlygate4sd3_1 hold66 (.A(\u_neuron.u_learning/_081_ ),
    .X(net108));
 sg13g2_dlygate4sd3_1 hold67 (.A(\u_neuron.fst_last_t[1] ),
    .X(net109));
 sg13g2_dlygate4sd3_1 hold68 (.A(_031_),
    .X(net110));
 sg13g2_dlygate4sd3_1 hold69 (.A(\u_neuron.wtab[15] ),
    .X(net111));
 sg13g2_dlygate4sd3_1 hold70 (.A(\u_neuron.td_prev[6] ),
    .X(net112));
 sg13g2_dlygate4sd3_1 hold71 (.A(_028_),
    .X(net113));
 sg13g2_dlygate4sd3_1 hold72 (.A(\u_neuron.td_prev[1] ),
    .X(net114));
 sg13g2_dlygate4sd3_1 hold73 (.A(_023_),
    .X(net115));
 sg13g2_dlygate4sd3_1 hold74 (.A(\u_neuron.fst_t[5] ),
    .X(net116));
 sg13g2_dlygate4sd3_1 hold75 (.A(_019_),
    .X(net117));
 sg13g2_dlygate4sd3_1 hold76 (.A(\u_neuron.td_prev[2] ),
    .X(net118));
 sg13g2_dlygate4sd3_1 hold77 (.A(_024_),
    .X(net119));
 sg13g2_dlygate4sd3_1 hold78 (.A(\u_neuron.lif_V[7] ),
    .X(net120));
 sg13g2_dlygate4sd3_1 hold79 (.A(_053_),
    .X(net121));
 sg13g2_dlygate4sd3_1 hold80 (.A(\u_neuron.pre_trace[11] ),
    .X(net122));
 sg13g2_dlygate4sd3_1 hold81 (.A(\u_neuron.fst_t[3] ),
    .X(net123));
 sg13g2_dlygate4sd3_1 hold82 (.A(\u_neuron.conv_shift[0] ),
    .X(net124));
 sg13g2_dlygate4sd3_1 hold83 (.A(_055_),
    .X(net125));
 sg13g2_dlygate4sd3_1 hold84 (.A(\u_neuron.td_prev[0] ),
    .X(net126));
 sg13g2_dlygate4sd3_1 hold85 (.A(_022_),
    .X(net127));
 sg13g2_dlygate4sd3_1 hold86 (.A(\u_neuron.wtab[9] ),
    .X(net128));
 sg13g2_dlygate4sd3_1 hold87 (.A(\u_neuron.wtab[19] ),
    .X(net129));
 sg13g2_dlygate4sd3_1 hold88 (.A(\u_neuron.fst_t[0] ),
    .X(net130));
 sg13g2_dlygate4sd3_1 hold89 (.A(\u_neuron.td_prev[7] ),
    .X(net131));
 sg13g2_dlygate4sd3_1 hold90 (.A(_029_),
    .X(net132));
 sg13g2_dlygate4sd3_1 hold91 (.A(\u_neuron.fst_t[7] ),
    .X(net133));
 sg13g2_dlygate4sd3_1 hold92 (.A(_021_),
    .X(net134));
 sg13g2_dlygate4sd3_1 hold93 (.A(\u_neuron.fst_t[2] ),
    .X(net135));
 sg13g2_dlygate4sd3_1 hold94 (.A(\u_neuron.fst_t[6] ),
    .X(net136));
 sg13g2_dlygate4sd3_1 hold95 (.A(_002_),
    .X(net137));
 sg13g2_dlygate4sd3_1 hold96 (.A(_242_),
    .X(net138));
 sg13g2_dlygate4sd3_1 hold97 (.A(_059_),
    .X(net139));
 sg13g2_dlygate4sd3_1 hold98 (.A(\u_neuron.td_prev[3] ),
    .X(net140));
 sg13g2_dlygate4sd3_1 hold99 (.A(_025_),
    .X(net141));
 sg13g2_dlygate4sd3_1 hold100 (.A(\u_neuron.lif_V[0] ),
    .X(net142));
 sg13g2_dlygate4sd3_1 hold101 (.A(_046_),
    .X(net143));
 sg13g2_dlygate4sd3_1 hold102 (.A(\u_neuron.td_prev[5] ),
    .X(net144));
 sg13g2_dlygate4sd3_1 hold103 (.A(_027_),
    .X(net145));
 sg13g2_dlygate4sd3_1 hold104 (.A(\u_neuron.wtab[31] ),
    .X(net146));
 sg13g2_dlygate4sd3_1 hold105 (.A(\u_neuron.wtab[23] ),
    .X(net147));
 sg13g2_dlygate4sd3_1 hold106 (.A(\u_neuron.wtab[22] ),
    .X(net148));
 sg13g2_dlygate4sd3_1 hold107 (.A(\u_neuron.lif_V[6] ),
    .X(net149));
 sg13g2_dlygate4sd3_1 hold108 (.A(_052_),
    .X(net150));
 sg13g2_dlygate4sd3_1 hold109 (.A(\u_neuron.td_prev[4] ),
    .X(net151));
 sg13g2_dlygate4sd3_1 hold110 (.A(_026_),
    .X(net152));
 sg13g2_dlygate4sd3_1 hold111 (.A(\u_neuron.td_curr[7] ),
    .X(net153));
 sg13g2_dlygate4sd3_1 hold112 (.A(_045_),
    .X(net154));
 sg13g2_dlygate4sd3_1 hold113 (.A(\u_neuron.td_curr[6] ),
    .X(net155));
 sg13g2_dlygate4sd3_1 hold114 (.A(\u_neuron.td_curr[0] ),
    .X(net156));
 sg13g2_dlygate4sd3_1 hold115 (.A(_038_),
    .X(net157));
 sg13g2_dlygate4sd3_1 hold116 (.A(\u_neuron.fst_armed ),
    .X(net158));
 sg13g2_dlygate4sd3_1 hold117 (.A(\u_neuron.fst_t[4] ),
    .X(net159));
 sg13g2_dlygate4sd3_1 hold118 (.A(uo_out[7]),
    .X(net160));
 sg13g2_dlygate4sd3_1 hold119 (.A(\u_neuron.lif_V[3] ),
    .X(net161));
 sg13g2_dlygate4sd3_1 hold120 (.A(\u_neuron.td_curr[5] ),
    .X(net162));
 sg13g2_dlygate4sd3_1 hold121 (.A(\u_neuron.wtab[8] ),
    .X(net163));
 sg13g2_dlygate4sd3_1 hold122 (.A(uo_out[6]),
    .X(net164));
 sg13g2_dlygate4sd3_1 hold123 (.A(\u_neuron.spike_seen_this_tick ),
    .X(net165));
 sg13g2_dlygate4sd3_1 hold124 (.A(\u_neuron.td_curr[2] ),
    .X(net166));
 sg13g2_dlygate4sd3_1 hold125 (.A(uo_out[5]),
    .X(net167));
 sg13g2_dlygate4sd3_1 hold126 (.A(uo_out[2]),
    .X(net168));
 sg13g2_dlygate4sd3_1 hold127 (.A(\u_neuron.wtab[3] ),
    .X(net169));
 sg13g2_dlygate4sd3_1 hold128 (.A(\u_neuron.td_curr[1] ),
    .X(net170));
 sg13g2_dlygate4sd3_1 hold129 (.A(uo_out[4]),
    .X(net171));
 sg13g2_dlygate4sd3_1 hold130 (.A(\u_neuron.wtab[13] ),
    .X(net172));
 sg13g2_dlygate4sd3_1 hold131 (.A(\u_neuron.lif_V[1] ),
    .X(net173));
 sg13g2_dlygate4sd3_1 hold132 (.A(\u_neuron.wtab[16] ),
    .X(net174));
 sg13g2_dlygate4sd3_1 hold133 (.A(uo_out[1]),
    .X(net175));
 sg13g2_dlygate4sd3_1 hold134 (.A(uo_out[3]),
    .X(net176));
 sg13g2_dlygate4sd3_1 hold135 (.A(\u_neuron.u_outq/_03_ ),
    .X(net177));
 sg13g2_dlygate4sd3_1 hold136 (.A(\u_neuron.td_curr[4] ),
    .X(net178));
 sg13g2_dlygate4sd3_1 hold137 (.A(\u_neuron.wtab[10] ),
    .X(net179));
 sg13g2_dlygate4sd3_1 hold138 (.A(uo_out[0]),
    .X(net180));
 sg13g2_dlygate4sd3_1 hold139 (.A(\u_neuron.conv_shift[1] ),
    .X(net181));
 sg13g2_dlygate4sd3_1 hold140 (.A(\u_neuron.td_curr[3] ),
    .X(net182));
 sg13g2_dlygate4sd3_1 hold141 (.A(\u_neuron.wtab[24] ),
    .X(net183));
 sg13g2_dlygate4sd3_1 hold142 (.A(\u_neuron.wtab[11] ),
    .X(net184));
 sg13g2_dlygate4sd3_1 hold143 (.A(\u_neuron.wtab[20] ),
    .X(net185));
 sg13g2_dlygate4sd3_1 hold144 (.A(\u_neuron.wtab[14] ),
    .X(net186));
 sg13g2_dlygate4sd3_1 hold145 (.A(\u_neuron.u_syn/_014_ ),
    .X(net187));
 sg13g2_dlygate4sd3_1 hold146 (.A(\u_neuron.wtab[1] ),
    .X(net188));
 sg13g2_dlygate4sd3_1 hold147 (.A(\u_neuron.wtab[28] ),
    .X(net189));
 sg13g2_dlygate4sd3_1 hold148 (.A(\u_neuron.wtab[6] ),
    .X(net190));
 sg13g2_dlygate4sd3_1 hold149 (.A(\u_neuron.lif_V[2] ),
    .X(net191));
 sg13g2_dlygate4sd3_1 hold150 (.A(\u_neuron.fst_t[1] ),
    .X(net192));
 sg13g2_dlygate4sd3_1 hold151 (.A(\u_neuron.wtab[25] ),
    .X(net193));
 sg13g2_dlygate4sd3_1 hold152 (.A(\u_neuron.wtab[30] ),
    .X(net194));
 sg13g2_dlygate4sd3_1 hold153 (.A(\u_neuron.lif_V[5] ),
    .X(net195));
 sg13g2_dlygate4sd3_1 hold154 (.A(\u_neuron.wtab[0] ),
    .X(net196));
 sg13g2_dlygate4sd3_1 hold155 (.A(\u_neuron.wtab[26] ),
    .X(net197));
 sg13g2_dlygate4sd3_1 hold156 (.A(\u_neuron.wtab[27] ),
    .X(net198));
 sg13g2_dlygate4sd3_1 hold157 (.A(\u_neuron.lif_V[4] ),
    .X(net199));
 sg13g2_dlygate4sd3_1 hold158 (.A(\u_neuron.learn_pending ),
    .X(net200));
 sg13g2_dlygate4sd3_1 hold159 (.A(\u_neuron.u_learning/_017_ ),
    .X(net201));
 sg13g2_dlygate4sd3_1 hold160 (.A(\u_neuron.wtab[5] ),
    .X(net202));
 sg13g2_dlygate4sd3_1 hold161 (.A(\u_neuron.wtab[7] ),
    .X(net203));
 sg13g2_dlygate4sd3_1 hold162 (.A(\u_neuron.wtab[18] ),
    .X(net204));
 sg13g2_dlygate4sd3_1 hold163 (.A(\u_neuron.wtab[17] ),
    .X(net205));
 sg13g2_dlygate4sd3_1 hold164 (.A(\u_neuron.post_trace ),
    .X(net206));
 sg13g2_dlygate4sd3_1 hold165 (.A(\u_neuron.wtab[12] ),
    .X(net207));
 sg13g2_dlygate4sd3_1 hold166 (.A(\u_neuron.wtab[21] ),
    .X(net208));
 sg13g2_dlygate4sd3_1 hold167 (.A(\u_neuron.learn_en ),
    .X(net209));
 sg13g2_dlygate4sd3_1 hold168 (.A(_054_),
    .X(net210));
 sg13g2_dlygate4sd3_1 hold169 (.A(\u_neuron.wtab[29] ),
    .X(net211));
 sg13g2_dlygate4sd3_1 hold170 (.A(\u_neuron.pre_trace[15] ),
    .X(net212));
 sg13g2_dlygate4sd3_1 hold171 (.A(\u_neuron.u_learning/_105_ ),
    .X(net213));
 sg13g2_dlygate4sd3_1 hold172 (.A(\u_neuron.u_learning/_015_ ),
    .X(net214));
 sg13g2_dlygate4sd3_1 hold173 (.A(\u_neuron.pending_widx[3] ),
    .X(net215));
 sg13g2_dlygate4sd3_1 hold174 (.A(\u_neuron.u_syn/_035_ ),
    .X(net216));
 sg13g2_dlygate4sd3_1 hold175 (.A(\u_neuron.wtab[4] ),
    .X(net217));
 sg13g2_dlygate4sd3_1 hold176 (.A(\u_neuron.learn_ptr[0] ),
    .X(net218));
 sg13g2_dlygate4sd3_1 hold177 (.A(\u_neuron.uio_in_sync[6] ),
    .X(net219));
 sg13g2_dlygate4sd3_1 hold178 (.A(\u_neuron.u_syn/_034_ ),
    .X(net220));
 sg13g2_dlygate4sd3_1 hold179 (.A(\u_neuron.uio_in_sync[4] ),
    .X(net221));
 sg13g2_dlygate4sd3_1 hold180 (.A(_243_),
    .X(net222));
 sg13g2_dlygate4sd3_1 hold181 (.A(_060_),
    .X(net223));
 sg13g2_dlygate4sd3_1 hold182 (.A(\u_neuron.learn_ptr[3] ),
    .X(net224));
 sg13g2_dlygate4sd3_1 hold183 (.A(\u_neuron.wtab[2] ),
    .X(net225));
 sg13g2_dlygate4sd3_1 hold184 (.A(\u_neuron.pending_widx[0] ),
    .X(net226));
 sg13g2_dlygate4sd3_1 hold185 (.A(\u_neuron.u_syn/_032_ ),
    .X(net227));
 sg13g2_dlygate4sd3_1 hold186 (.A(\u_neuron.uio_in_sync[5] ),
    .X(net228));
 sg13g2_dlygate4sd3_1 hold187 (.A(\u_neuron.u_syn/_403_ ),
    .X(net229));
 sg13g2_dlygate4sd3_1 hold188 (.A(\u_neuron.u_syn/_033_ ),
    .X(net230));
 sg13g2_dlygate4sd3_1 hold189 (.A(\u_neuron.mode[1] ),
    .X(net231));
 sg13g2_dlygate4sd3_1 hold190 (.A(_061_),
    .X(net232));
 sg13g2_dlygate4sd3_1 hold191 (.A(\u_neuron.have_out ),
    .X(net233));
 sg13g2_dlygate4sd3_1 hold192 (.A(\u_neuron.u_outq/_08_ ),
    .X(net234));
 sg13g2_dlygate4sd3_1 hold193 (.A(\u_neuron.learn_pending ),
    .X(net235));
 sg13g2_dlygate4sd3_1 hold194 (.A(\u_neuron.conv_shift[0] ),
    .X(net236));
 sg13g2_dlygate4sd3_1 hold195 (.A(\u_neuron.spike_seen_this_tick ),
    .X(net237));
 sg13g2_dlygate4sd3_1 hold196 (.A(\u_neuron.pending_widx[0] ),
    .X(net238));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_fill_2 FILLER_0_406 ();
 sg13g2_fill_1 FILLER_0_408 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_fill_2 FILLER_1_406 ();
 sg13g2_fill_1 FILLER_1_408 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_fill_2 FILLER_2_329 ();
 sg13g2_fill_1 FILLER_2_331 ();
 sg13g2_decap_8 FILLER_2_359 ();
 sg13g2_decap_8 FILLER_2_366 ();
 sg13g2_decap_8 FILLER_2_373 ();
 sg13g2_decap_8 FILLER_2_380 ();
 sg13g2_decap_8 FILLER_2_387 ();
 sg13g2_decap_8 FILLER_2_394 ();
 sg13g2_decap_8 FILLER_2_401 ();
 sg13g2_fill_1 FILLER_2_408 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_252 ();
 sg13g2_decap_8 FILLER_3_259 ();
 sg13g2_decap_8 FILLER_3_266 ();
 sg13g2_decap_8 FILLER_3_273 ();
 sg13g2_decap_8 FILLER_3_280 ();
 sg13g2_decap_8 FILLER_3_287 ();
 sg13g2_decap_8 FILLER_3_294 ();
 sg13g2_decap_8 FILLER_3_301 ();
 sg13g2_decap_4 FILLER_3_308 ();
 sg13g2_decap_8 FILLER_3_366 ();
 sg13g2_decap_8 FILLER_3_373 ();
 sg13g2_decap_8 FILLER_3_380 ();
 sg13g2_decap_8 FILLER_3_387 ();
 sg13g2_decap_8 FILLER_3_394 ();
 sg13g2_decap_8 FILLER_3_401 ();
 sg13g2_fill_1 FILLER_3_408 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_224 ();
 sg13g2_decap_8 FILLER_4_231 ();
 sg13g2_decap_8 FILLER_4_238 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_decap_8 FILLER_4_252 ();
 sg13g2_decap_8 FILLER_4_259 ();
 sg13g2_decap_8 FILLER_4_266 ();
 sg13g2_decap_8 FILLER_4_273 ();
 sg13g2_decap_8 FILLER_4_280 ();
 sg13g2_decap_8 FILLER_4_287 ();
 sg13g2_fill_2 FILLER_4_294 ();
 sg13g2_fill_2 FILLER_4_347 ();
 sg13g2_decap_8 FILLER_4_362 ();
 sg13g2_decap_8 FILLER_4_369 ();
 sg13g2_decap_8 FILLER_4_376 ();
 sg13g2_decap_8 FILLER_4_383 ();
 sg13g2_decap_8 FILLER_4_390 ();
 sg13g2_decap_8 FILLER_4_397 ();
 sg13g2_decap_4 FILLER_4_404 ();
 sg13g2_fill_1 FILLER_4_408 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_decap_8 FILLER_5_175 ();
 sg13g2_decap_8 FILLER_5_182 ();
 sg13g2_decap_8 FILLER_5_189 ();
 sg13g2_decap_8 FILLER_5_196 ();
 sg13g2_decap_8 FILLER_5_203 ();
 sg13g2_decap_8 FILLER_5_210 ();
 sg13g2_decap_8 FILLER_5_217 ();
 sg13g2_decap_8 FILLER_5_224 ();
 sg13g2_decap_8 FILLER_5_231 ();
 sg13g2_decap_8 FILLER_5_238 ();
 sg13g2_decap_8 FILLER_5_245 ();
 sg13g2_decap_8 FILLER_5_252 ();
 sg13g2_decap_8 FILLER_5_259 ();
 sg13g2_decap_8 FILLER_5_266 ();
 sg13g2_decap_8 FILLER_5_273 ();
 sg13g2_decap_8 FILLER_5_280 ();
 sg13g2_decap_8 FILLER_5_287 ();
 sg13g2_decap_8 FILLER_5_294 ();
 sg13g2_fill_2 FILLER_5_301 ();
 sg13g2_decap_8 FILLER_5_365 ();
 sg13g2_decap_8 FILLER_5_372 ();
 sg13g2_decap_8 FILLER_5_379 ();
 sg13g2_decap_8 FILLER_5_386 ();
 sg13g2_decap_8 FILLER_5_393 ();
 sg13g2_decap_8 FILLER_5_400 ();
 sg13g2_fill_2 FILLER_5_407 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_147 ();
 sg13g2_decap_8 FILLER_6_154 ();
 sg13g2_decap_8 FILLER_6_161 ();
 sg13g2_decap_8 FILLER_6_168 ();
 sg13g2_decap_8 FILLER_6_175 ();
 sg13g2_decap_8 FILLER_6_182 ();
 sg13g2_decap_8 FILLER_6_189 ();
 sg13g2_decap_8 FILLER_6_196 ();
 sg13g2_decap_8 FILLER_6_203 ();
 sg13g2_decap_8 FILLER_6_210 ();
 sg13g2_decap_8 FILLER_6_217 ();
 sg13g2_decap_8 FILLER_6_224 ();
 sg13g2_decap_8 FILLER_6_231 ();
 sg13g2_decap_8 FILLER_6_238 ();
 sg13g2_decap_8 FILLER_6_245 ();
 sg13g2_decap_8 FILLER_6_252 ();
 sg13g2_decap_8 FILLER_6_259 ();
 sg13g2_decap_8 FILLER_6_266 ();
 sg13g2_decap_8 FILLER_6_273 ();
 sg13g2_decap_8 FILLER_6_280 ();
 sg13g2_decap_8 FILLER_6_287 ();
 sg13g2_decap_8 FILLER_6_294 ();
 sg13g2_decap_4 FILLER_6_301 ();
 sg13g2_decap_4 FILLER_6_310 ();
 sg13g2_fill_1 FILLER_6_318 ();
 sg13g2_decap_4 FILLER_6_323 ();
 sg13g2_fill_1 FILLER_6_327 ();
 sg13g2_decap_8 FILLER_6_349 ();
 sg13g2_decap_8 FILLER_6_356 ();
 sg13g2_decap_8 FILLER_6_363 ();
 sg13g2_decap_8 FILLER_6_370 ();
 sg13g2_decap_8 FILLER_6_377 ();
 sg13g2_decap_8 FILLER_6_384 ();
 sg13g2_decap_8 FILLER_6_391 ();
 sg13g2_decap_8 FILLER_6_398 ();
 sg13g2_decap_4 FILLER_6_405 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_8 FILLER_7_140 ();
 sg13g2_decap_8 FILLER_7_147 ();
 sg13g2_decap_8 FILLER_7_154 ();
 sg13g2_decap_8 FILLER_7_161 ();
 sg13g2_decap_8 FILLER_7_168 ();
 sg13g2_decap_8 FILLER_7_175 ();
 sg13g2_decap_8 FILLER_7_182 ();
 sg13g2_decap_8 FILLER_7_189 ();
 sg13g2_decap_8 FILLER_7_196 ();
 sg13g2_decap_8 FILLER_7_203 ();
 sg13g2_decap_8 FILLER_7_210 ();
 sg13g2_decap_8 FILLER_7_217 ();
 sg13g2_decap_8 FILLER_7_224 ();
 sg13g2_decap_8 FILLER_7_231 ();
 sg13g2_decap_8 FILLER_7_238 ();
 sg13g2_decap_8 FILLER_7_245 ();
 sg13g2_decap_8 FILLER_7_252 ();
 sg13g2_decap_8 FILLER_7_259 ();
 sg13g2_decap_8 FILLER_7_266 ();
 sg13g2_decap_8 FILLER_7_273 ();
 sg13g2_decap_8 FILLER_7_280 ();
 sg13g2_decap_8 FILLER_7_287 ();
 sg13g2_decap_8 FILLER_7_294 ();
 sg13g2_decap_8 FILLER_7_301 ();
 sg13g2_fill_1 FILLER_7_308 ();
 sg13g2_fill_1 FILLER_7_328 ();
 sg13g2_fill_2 FILLER_7_334 ();
 sg13g2_decap_8 FILLER_7_372 ();
 sg13g2_decap_8 FILLER_7_379 ();
 sg13g2_decap_8 FILLER_7_386 ();
 sg13g2_decap_8 FILLER_7_393 ();
 sg13g2_decap_8 FILLER_7_400 ();
 sg13g2_fill_2 FILLER_7_407 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_decap_8 FILLER_8_119 ();
 sg13g2_decap_8 FILLER_8_126 ();
 sg13g2_decap_8 FILLER_8_133 ();
 sg13g2_decap_8 FILLER_8_140 ();
 sg13g2_decap_8 FILLER_8_147 ();
 sg13g2_decap_8 FILLER_8_154 ();
 sg13g2_decap_8 FILLER_8_161 ();
 sg13g2_decap_8 FILLER_8_168 ();
 sg13g2_decap_8 FILLER_8_175 ();
 sg13g2_decap_8 FILLER_8_182 ();
 sg13g2_decap_8 FILLER_8_189 ();
 sg13g2_decap_8 FILLER_8_196 ();
 sg13g2_decap_8 FILLER_8_203 ();
 sg13g2_decap_8 FILLER_8_210 ();
 sg13g2_decap_8 FILLER_8_217 ();
 sg13g2_decap_8 FILLER_8_224 ();
 sg13g2_decap_8 FILLER_8_231 ();
 sg13g2_decap_8 FILLER_8_238 ();
 sg13g2_decap_8 FILLER_8_245 ();
 sg13g2_decap_8 FILLER_8_252 ();
 sg13g2_decap_8 FILLER_8_259 ();
 sg13g2_decap_8 FILLER_8_266 ();
 sg13g2_decap_8 FILLER_8_273 ();
 sg13g2_decap_8 FILLER_8_280 ();
 sg13g2_decap_4 FILLER_8_287 ();
 sg13g2_decap_4 FILLER_8_352 ();
 sg13g2_fill_2 FILLER_8_356 ();
 sg13g2_decap_8 FILLER_8_367 ();
 sg13g2_decap_8 FILLER_8_374 ();
 sg13g2_decap_8 FILLER_8_381 ();
 sg13g2_decap_8 FILLER_8_388 ();
 sg13g2_decap_8 FILLER_8_395 ();
 sg13g2_decap_8 FILLER_8_402 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_91 ();
 sg13g2_decap_8 FILLER_9_98 ();
 sg13g2_decap_8 FILLER_9_105 ();
 sg13g2_decap_8 FILLER_9_112 ();
 sg13g2_decap_8 FILLER_9_119 ();
 sg13g2_decap_8 FILLER_9_126 ();
 sg13g2_decap_8 FILLER_9_133 ();
 sg13g2_decap_8 FILLER_9_140 ();
 sg13g2_decap_8 FILLER_9_147 ();
 sg13g2_decap_8 FILLER_9_154 ();
 sg13g2_decap_8 FILLER_9_161 ();
 sg13g2_decap_8 FILLER_9_168 ();
 sg13g2_decap_8 FILLER_9_175 ();
 sg13g2_decap_8 FILLER_9_182 ();
 sg13g2_decap_8 FILLER_9_189 ();
 sg13g2_decap_8 FILLER_9_196 ();
 sg13g2_decap_8 FILLER_9_203 ();
 sg13g2_decap_8 FILLER_9_210 ();
 sg13g2_decap_8 FILLER_9_217 ();
 sg13g2_decap_8 FILLER_9_224 ();
 sg13g2_decap_8 FILLER_9_231 ();
 sg13g2_decap_8 FILLER_9_238 ();
 sg13g2_decap_8 FILLER_9_245 ();
 sg13g2_decap_8 FILLER_9_252 ();
 sg13g2_decap_8 FILLER_9_259 ();
 sg13g2_decap_8 FILLER_9_266 ();
 sg13g2_decap_8 FILLER_9_273 ();
 sg13g2_decap_8 FILLER_9_280 ();
 sg13g2_decap_8 FILLER_9_287 ();
 sg13g2_fill_1 FILLER_9_294 ();
 sg13g2_decap_8 FILLER_9_347 ();
 sg13g2_decap_8 FILLER_9_354 ();
 sg13g2_fill_1 FILLER_9_361 ();
 sg13g2_decap_8 FILLER_9_375 ();
 sg13g2_decap_8 FILLER_9_382 ();
 sg13g2_decap_8 FILLER_9_389 ();
 sg13g2_decap_8 FILLER_9_396 ();
 sg13g2_decap_4 FILLER_9_403 ();
 sg13g2_fill_2 FILLER_9_407 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_decap_8 FILLER_10_77 ();
 sg13g2_decap_8 FILLER_10_84 ();
 sg13g2_decap_8 FILLER_10_91 ();
 sg13g2_decap_8 FILLER_10_98 ();
 sg13g2_decap_8 FILLER_10_105 ();
 sg13g2_decap_8 FILLER_10_112 ();
 sg13g2_decap_8 FILLER_10_119 ();
 sg13g2_decap_8 FILLER_10_126 ();
 sg13g2_decap_8 FILLER_10_133 ();
 sg13g2_decap_8 FILLER_10_140 ();
 sg13g2_decap_8 FILLER_10_147 ();
 sg13g2_decap_8 FILLER_10_154 ();
 sg13g2_decap_8 FILLER_10_161 ();
 sg13g2_decap_8 FILLER_10_168 ();
 sg13g2_decap_8 FILLER_10_175 ();
 sg13g2_decap_8 FILLER_10_182 ();
 sg13g2_decap_8 FILLER_10_189 ();
 sg13g2_decap_8 FILLER_10_196 ();
 sg13g2_decap_8 FILLER_10_203 ();
 sg13g2_decap_8 FILLER_10_210 ();
 sg13g2_decap_8 FILLER_10_217 ();
 sg13g2_decap_8 FILLER_10_224 ();
 sg13g2_decap_8 FILLER_10_231 ();
 sg13g2_decap_8 FILLER_10_238 ();
 sg13g2_decap_8 FILLER_10_245 ();
 sg13g2_decap_8 FILLER_10_252 ();
 sg13g2_decap_8 FILLER_10_259 ();
 sg13g2_decap_8 FILLER_10_266 ();
 sg13g2_decap_8 FILLER_10_273 ();
 sg13g2_decap_8 FILLER_10_280 ();
 sg13g2_fill_2 FILLER_10_287 ();
 sg13g2_fill_1 FILLER_10_289 ();
 sg13g2_decap_8 FILLER_10_294 ();
 sg13g2_fill_2 FILLER_10_301 ();
 sg13g2_decap_4 FILLER_10_308 ();
 sg13g2_fill_1 FILLER_10_312 ();
 sg13g2_decap_4 FILLER_10_323 ();
 sg13g2_fill_2 FILLER_10_327 ();
 sg13g2_fill_2 FILLER_10_332 ();
 sg13g2_decap_8 FILLER_10_384 ();
 sg13g2_decap_8 FILLER_10_391 ();
 sg13g2_decap_8 FILLER_10_398 ();
 sg13g2_decap_4 FILLER_10_405 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_63 ();
 sg13g2_decap_8 FILLER_11_70 ();
 sg13g2_decap_8 FILLER_11_77 ();
 sg13g2_decap_8 FILLER_11_84 ();
 sg13g2_decap_8 FILLER_11_91 ();
 sg13g2_decap_8 FILLER_11_98 ();
 sg13g2_decap_8 FILLER_11_105 ();
 sg13g2_decap_8 FILLER_11_112 ();
 sg13g2_decap_8 FILLER_11_119 ();
 sg13g2_decap_8 FILLER_11_126 ();
 sg13g2_decap_8 FILLER_11_133 ();
 sg13g2_decap_8 FILLER_11_140 ();
 sg13g2_decap_8 FILLER_11_147 ();
 sg13g2_decap_8 FILLER_11_154 ();
 sg13g2_decap_8 FILLER_11_161 ();
 sg13g2_decap_8 FILLER_11_168 ();
 sg13g2_decap_8 FILLER_11_175 ();
 sg13g2_decap_8 FILLER_11_182 ();
 sg13g2_decap_8 FILLER_11_189 ();
 sg13g2_decap_8 FILLER_11_196 ();
 sg13g2_decap_8 FILLER_11_203 ();
 sg13g2_decap_8 FILLER_11_210 ();
 sg13g2_decap_8 FILLER_11_217 ();
 sg13g2_decap_8 FILLER_11_224 ();
 sg13g2_decap_8 FILLER_11_231 ();
 sg13g2_decap_8 FILLER_11_238 ();
 sg13g2_decap_8 FILLER_11_245 ();
 sg13g2_decap_8 FILLER_11_252 ();
 sg13g2_decap_8 FILLER_11_259 ();
 sg13g2_fill_1 FILLER_11_266 ();
 sg13g2_fill_1 FILLER_11_294 ();
 sg13g2_fill_2 FILLER_11_300 ();
 sg13g2_fill_1 FILLER_11_302 ();
 sg13g2_decap_8 FILLER_11_313 ();
 sg13g2_decap_8 FILLER_11_320 ();
 sg13g2_fill_1 FILLER_11_327 ();
 sg13g2_fill_2 FILLER_11_347 ();
 sg13g2_decap_8 FILLER_11_376 ();
 sg13g2_decap_8 FILLER_11_383 ();
 sg13g2_decap_8 FILLER_11_390 ();
 sg13g2_decap_8 FILLER_11_397 ();
 sg13g2_decap_4 FILLER_11_404 ();
 sg13g2_fill_1 FILLER_11_408 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_decap_8 FILLER_12_56 ();
 sg13g2_decap_8 FILLER_12_63 ();
 sg13g2_decap_8 FILLER_12_70 ();
 sg13g2_decap_8 FILLER_12_77 ();
 sg13g2_decap_8 FILLER_12_84 ();
 sg13g2_decap_8 FILLER_12_91 ();
 sg13g2_decap_8 FILLER_12_98 ();
 sg13g2_decap_8 FILLER_12_105 ();
 sg13g2_decap_8 FILLER_12_112 ();
 sg13g2_decap_8 FILLER_12_119 ();
 sg13g2_decap_8 FILLER_12_126 ();
 sg13g2_decap_8 FILLER_12_133 ();
 sg13g2_decap_8 FILLER_12_140 ();
 sg13g2_decap_8 FILLER_12_147 ();
 sg13g2_decap_8 FILLER_12_154 ();
 sg13g2_decap_8 FILLER_12_161 ();
 sg13g2_decap_8 FILLER_12_168 ();
 sg13g2_decap_8 FILLER_12_175 ();
 sg13g2_decap_8 FILLER_12_182 ();
 sg13g2_decap_8 FILLER_12_189 ();
 sg13g2_decap_8 FILLER_12_196 ();
 sg13g2_decap_8 FILLER_12_203 ();
 sg13g2_decap_8 FILLER_12_210 ();
 sg13g2_decap_8 FILLER_12_217 ();
 sg13g2_decap_8 FILLER_12_224 ();
 sg13g2_decap_8 FILLER_12_231 ();
 sg13g2_decap_8 FILLER_12_238 ();
 sg13g2_decap_8 FILLER_12_245 ();
 sg13g2_decap_8 FILLER_12_252 ();
 sg13g2_decap_8 FILLER_12_259 ();
 sg13g2_decap_4 FILLER_12_266 ();
 sg13g2_fill_2 FILLER_12_312 ();
 sg13g2_fill_1 FILLER_12_318 ();
 sg13g2_fill_1 FILLER_12_347 ();
 sg13g2_decap_8 FILLER_12_375 ();
 sg13g2_decap_8 FILLER_12_382 ();
 sg13g2_decap_8 FILLER_12_389 ();
 sg13g2_decap_8 FILLER_12_396 ();
 sg13g2_decap_4 FILLER_12_403 ();
 sg13g2_fill_2 FILLER_12_407 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_decap_8 FILLER_13_49 ();
 sg13g2_decap_8 FILLER_13_56 ();
 sg13g2_decap_8 FILLER_13_63 ();
 sg13g2_decap_8 FILLER_13_70 ();
 sg13g2_decap_8 FILLER_13_77 ();
 sg13g2_decap_8 FILLER_13_84 ();
 sg13g2_decap_8 FILLER_13_91 ();
 sg13g2_decap_8 FILLER_13_98 ();
 sg13g2_decap_8 FILLER_13_105 ();
 sg13g2_decap_8 FILLER_13_112 ();
 sg13g2_decap_8 FILLER_13_119 ();
 sg13g2_decap_8 FILLER_13_126 ();
 sg13g2_decap_8 FILLER_13_133 ();
 sg13g2_decap_8 FILLER_13_140 ();
 sg13g2_decap_8 FILLER_13_147 ();
 sg13g2_decap_8 FILLER_13_154 ();
 sg13g2_decap_8 FILLER_13_161 ();
 sg13g2_decap_8 FILLER_13_168 ();
 sg13g2_decap_8 FILLER_13_175 ();
 sg13g2_decap_8 FILLER_13_182 ();
 sg13g2_decap_8 FILLER_13_189 ();
 sg13g2_decap_8 FILLER_13_196 ();
 sg13g2_decap_8 FILLER_13_203 ();
 sg13g2_decap_8 FILLER_13_210 ();
 sg13g2_decap_8 FILLER_13_217 ();
 sg13g2_decap_8 FILLER_13_224 ();
 sg13g2_decap_8 FILLER_13_231 ();
 sg13g2_decap_8 FILLER_13_238 ();
 sg13g2_decap_8 FILLER_13_245 ();
 sg13g2_decap_8 FILLER_13_252 ();
 sg13g2_decap_8 FILLER_13_259 ();
 sg13g2_fill_2 FILLER_13_266 ();
 sg13g2_fill_1 FILLER_13_304 ();
 sg13g2_decap_8 FILLER_13_369 ();
 sg13g2_decap_8 FILLER_13_376 ();
 sg13g2_decap_8 FILLER_13_383 ();
 sg13g2_decap_8 FILLER_13_390 ();
 sg13g2_decap_8 FILLER_13_397 ();
 sg13g2_decap_4 FILLER_13_404 ();
 sg13g2_fill_1 FILLER_13_408 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_decap_8 FILLER_14_42 ();
 sg13g2_decap_8 FILLER_14_49 ();
 sg13g2_decap_8 FILLER_14_56 ();
 sg13g2_decap_8 FILLER_14_63 ();
 sg13g2_decap_8 FILLER_14_70 ();
 sg13g2_decap_8 FILLER_14_77 ();
 sg13g2_decap_8 FILLER_14_84 ();
 sg13g2_decap_8 FILLER_14_91 ();
 sg13g2_decap_8 FILLER_14_98 ();
 sg13g2_decap_8 FILLER_14_105 ();
 sg13g2_decap_8 FILLER_14_112 ();
 sg13g2_decap_8 FILLER_14_119 ();
 sg13g2_decap_8 FILLER_14_126 ();
 sg13g2_decap_8 FILLER_14_133 ();
 sg13g2_decap_8 FILLER_14_140 ();
 sg13g2_decap_8 FILLER_14_147 ();
 sg13g2_decap_8 FILLER_14_154 ();
 sg13g2_decap_8 FILLER_14_161 ();
 sg13g2_decap_8 FILLER_14_168 ();
 sg13g2_decap_8 FILLER_14_175 ();
 sg13g2_decap_8 FILLER_14_182 ();
 sg13g2_decap_8 FILLER_14_189 ();
 sg13g2_decap_8 FILLER_14_196 ();
 sg13g2_decap_8 FILLER_14_203 ();
 sg13g2_decap_8 FILLER_14_210 ();
 sg13g2_decap_8 FILLER_14_217 ();
 sg13g2_decap_8 FILLER_14_224 ();
 sg13g2_decap_8 FILLER_14_231 ();
 sg13g2_decap_8 FILLER_14_238 ();
 sg13g2_decap_8 FILLER_14_245 ();
 sg13g2_decap_8 FILLER_14_252 ();
 sg13g2_decap_8 FILLER_14_259 ();
 sg13g2_decap_4 FILLER_14_266 ();
 sg13g2_fill_2 FILLER_14_286 ();
 sg13g2_fill_1 FILLER_14_288 ();
 sg13g2_fill_2 FILLER_14_299 ();
 sg13g2_fill_1 FILLER_14_301 ();
 sg13g2_fill_1 FILLER_14_326 ();
 sg13g2_decap_8 FILLER_14_370 ();
 sg13g2_decap_8 FILLER_14_377 ();
 sg13g2_decap_8 FILLER_14_384 ();
 sg13g2_decap_8 FILLER_14_391 ();
 sg13g2_decap_8 FILLER_14_398 ();
 sg13g2_decap_4 FILLER_14_405 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_8 FILLER_15_35 ();
 sg13g2_decap_8 FILLER_15_42 ();
 sg13g2_decap_8 FILLER_15_49 ();
 sg13g2_decap_8 FILLER_15_56 ();
 sg13g2_decap_8 FILLER_15_63 ();
 sg13g2_decap_8 FILLER_15_70 ();
 sg13g2_decap_8 FILLER_15_77 ();
 sg13g2_decap_8 FILLER_15_84 ();
 sg13g2_decap_8 FILLER_15_91 ();
 sg13g2_decap_8 FILLER_15_98 ();
 sg13g2_decap_8 FILLER_15_105 ();
 sg13g2_decap_8 FILLER_15_112 ();
 sg13g2_decap_8 FILLER_15_119 ();
 sg13g2_decap_8 FILLER_15_126 ();
 sg13g2_decap_8 FILLER_15_133 ();
 sg13g2_decap_8 FILLER_15_140 ();
 sg13g2_decap_8 FILLER_15_147 ();
 sg13g2_decap_8 FILLER_15_154 ();
 sg13g2_decap_8 FILLER_15_161 ();
 sg13g2_decap_8 FILLER_15_168 ();
 sg13g2_decap_8 FILLER_15_175 ();
 sg13g2_decap_8 FILLER_15_182 ();
 sg13g2_decap_8 FILLER_15_189 ();
 sg13g2_decap_8 FILLER_15_196 ();
 sg13g2_decap_8 FILLER_15_203 ();
 sg13g2_decap_8 FILLER_15_210 ();
 sg13g2_decap_8 FILLER_15_217 ();
 sg13g2_decap_8 FILLER_15_224 ();
 sg13g2_decap_8 FILLER_15_231 ();
 sg13g2_decap_8 FILLER_15_238 ();
 sg13g2_decap_8 FILLER_15_245 ();
 sg13g2_decap_8 FILLER_15_252 ();
 sg13g2_decap_8 FILLER_15_259 ();
 sg13g2_fill_1 FILLER_15_266 ();
 sg13g2_fill_2 FILLER_15_294 ();
 sg13g2_fill_1 FILLER_15_296 ();
 sg13g2_fill_2 FILLER_15_310 ();
 sg13g2_fill_1 FILLER_15_312 ();
 sg13g2_decap_4 FILLER_15_321 ();
 sg13g2_fill_2 FILLER_15_355 ();
 sg13g2_fill_1 FILLER_15_357 ();
 sg13g2_fill_2 FILLER_15_361 ();
 sg13g2_fill_1 FILLER_15_363 ();
 sg13g2_decap_8 FILLER_15_373 ();
 sg13g2_decap_8 FILLER_15_380 ();
 sg13g2_decap_8 FILLER_15_387 ();
 sg13g2_decap_8 FILLER_15_394 ();
 sg13g2_decap_8 FILLER_15_401 ();
 sg13g2_fill_1 FILLER_15_408 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_decap_8 FILLER_16_35 ();
 sg13g2_decap_8 FILLER_16_42 ();
 sg13g2_decap_8 FILLER_16_49 ();
 sg13g2_decap_8 FILLER_16_56 ();
 sg13g2_decap_8 FILLER_16_63 ();
 sg13g2_decap_8 FILLER_16_70 ();
 sg13g2_decap_8 FILLER_16_77 ();
 sg13g2_decap_8 FILLER_16_84 ();
 sg13g2_decap_8 FILLER_16_91 ();
 sg13g2_decap_8 FILLER_16_98 ();
 sg13g2_decap_8 FILLER_16_105 ();
 sg13g2_decap_8 FILLER_16_112 ();
 sg13g2_decap_8 FILLER_16_119 ();
 sg13g2_decap_8 FILLER_16_126 ();
 sg13g2_decap_4 FILLER_16_133 ();
 sg13g2_fill_2 FILLER_16_137 ();
 sg13g2_fill_2 FILLER_16_167 ();
 sg13g2_fill_1 FILLER_16_169 ();
 sg13g2_decap_8 FILLER_16_198 ();
 sg13g2_decap_8 FILLER_16_205 ();
 sg13g2_decap_8 FILLER_16_212 ();
 sg13g2_decap_8 FILLER_16_219 ();
 sg13g2_decap_8 FILLER_16_226 ();
 sg13g2_decap_8 FILLER_16_233 ();
 sg13g2_decap_8 FILLER_16_240 ();
 sg13g2_decap_8 FILLER_16_247 ();
 sg13g2_decap_8 FILLER_16_254 ();
 sg13g2_decap_8 FILLER_16_261 ();
 sg13g2_decap_8 FILLER_16_268 ();
 sg13g2_decap_8 FILLER_16_275 ();
 sg13g2_decap_4 FILLER_16_282 ();
 sg13g2_fill_2 FILLER_16_296 ();
 sg13g2_fill_2 FILLER_16_327 ();
 sg13g2_fill_1 FILLER_16_329 ();
 sg13g2_fill_2 FILLER_16_336 ();
 sg13g2_fill_1 FILLER_16_338 ();
 sg13g2_decap_8 FILLER_16_374 ();
 sg13g2_decap_8 FILLER_16_381 ();
 sg13g2_decap_8 FILLER_16_388 ();
 sg13g2_decap_8 FILLER_16_395 ();
 sg13g2_decap_8 FILLER_16_402 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_28 ();
 sg13g2_decap_8 FILLER_17_35 ();
 sg13g2_decap_8 FILLER_17_42 ();
 sg13g2_decap_8 FILLER_17_49 ();
 sg13g2_decap_8 FILLER_17_56 ();
 sg13g2_decap_8 FILLER_17_63 ();
 sg13g2_decap_8 FILLER_17_70 ();
 sg13g2_decap_8 FILLER_17_77 ();
 sg13g2_decap_8 FILLER_17_84 ();
 sg13g2_decap_8 FILLER_17_91 ();
 sg13g2_decap_8 FILLER_17_98 ();
 sg13g2_decap_8 FILLER_17_105 ();
 sg13g2_decap_8 FILLER_17_112 ();
 sg13g2_decap_8 FILLER_17_119 ();
 sg13g2_fill_1 FILLER_17_126 ();
 sg13g2_decap_8 FILLER_17_211 ();
 sg13g2_decap_8 FILLER_17_218 ();
 sg13g2_decap_8 FILLER_17_225 ();
 sg13g2_decap_8 FILLER_17_232 ();
 sg13g2_decap_8 FILLER_17_239 ();
 sg13g2_decap_8 FILLER_17_246 ();
 sg13g2_decap_8 FILLER_17_253 ();
 sg13g2_decap_8 FILLER_17_260 ();
 sg13g2_decap_8 FILLER_17_267 ();
 sg13g2_decap_8 FILLER_17_274 ();
 sg13g2_decap_8 FILLER_17_281 ();
 sg13g2_decap_8 FILLER_17_288 ();
 sg13g2_fill_1 FILLER_17_295 ();
 sg13g2_decap_8 FILLER_17_311 ();
 sg13g2_decap_4 FILLER_17_326 ();
 sg13g2_fill_1 FILLER_17_330 ();
 sg13g2_fill_2 FILLER_17_336 ();
 sg13g2_decap_8 FILLER_17_348 ();
 sg13g2_decap_8 FILLER_17_355 ();
 sg13g2_decap_8 FILLER_17_362 ();
 sg13g2_decap_8 FILLER_17_369 ();
 sg13g2_decap_8 FILLER_17_376 ();
 sg13g2_decap_8 FILLER_17_383 ();
 sg13g2_decap_8 FILLER_17_390 ();
 sg13g2_decap_8 FILLER_17_397 ();
 sg13g2_decap_4 FILLER_17_404 ();
 sg13g2_fill_1 FILLER_17_408 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_21 ();
 sg13g2_decap_8 FILLER_18_28 ();
 sg13g2_decap_8 FILLER_18_35 ();
 sg13g2_decap_8 FILLER_18_42 ();
 sg13g2_decap_8 FILLER_18_49 ();
 sg13g2_decap_8 FILLER_18_56 ();
 sg13g2_decap_8 FILLER_18_63 ();
 sg13g2_decap_8 FILLER_18_70 ();
 sg13g2_decap_8 FILLER_18_77 ();
 sg13g2_decap_8 FILLER_18_84 ();
 sg13g2_decap_8 FILLER_18_91 ();
 sg13g2_decap_8 FILLER_18_98 ();
 sg13g2_decap_8 FILLER_18_105 ();
 sg13g2_decap_8 FILLER_18_112 ();
 sg13g2_decap_8 FILLER_18_119 ();
 sg13g2_decap_4 FILLER_18_126 ();
 sg13g2_fill_2 FILLER_18_130 ();
 sg13g2_fill_1 FILLER_18_141 ();
 sg13g2_fill_2 FILLER_18_188 ();
 sg13g2_fill_1 FILLER_18_190 ();
 sg13g2_decap_8 FILLER_18_200 ();
 sg13g2_decap_8 FILLER_18_207 ();
 sg13g2_decap_8 FILLER_18_214 ();
 sg13g2_decap_8 FILLER_18_221 ();
 sg13g2_decap_8 FILLER_18_228 ();
 sg13g2_decap_8 FILLER_18_235 ();
 sg13g2_decap_8 FILLER_18_242 ();
 sg13g2_decap_8 FILLER_18_249 ();
 sg13g2_decap_8 FILLER_18_256 ();
 sg13g2_decap_8 FILLER_18_263 ();
 sg13g2_decap_8 FILLER_18_270 ();
 sg13g2_decap_8 FILLER_18_277 ();
 sg13g2_decap_8 FILLER_18_284 ();
 sg13g2_decap_4 FILLER_18_291 ();
 sg13g2_fill_2 FILLER_18_295 ();
 sg13g2_fill_2 FILLER_18_322 ();
 sg13g2_fill_1 FILLER_18_324 ();
 sg13g2_decap_4 FILLER_18_337 ();
 sg13g2_decap_8 FILLER_18_356 ();
 sg13g2_decap_8 FILLER_18_363 ();
 sg13g2_decap_8 FILLER_18_370 ();
 sg13g2_decap_8 FILLER_18_377 ();
 sg13g2_decap_8 FILLER_18_384 ();
 sg13g2_decap_8 FILLER_18_391 ();
 sg13g2_decap_8 FILLER_18_398 ();
 sg13g2_decap_4 FILLER_18_405 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_decap_8 FILLER_19_28 ();
 sg13g2_decap_8 FILLER_19_35 ();
 sg13g2_decap_8 FILLER_19_42 ();
 sg13g2_decap_8 FILLER_19_49 ();
 sg13g2_decap_8 FILLER_19_56 ();
 sg13g2_decap_8 FILLER_19_63 ();
 sg13g2_decap_8 FILLER_19_70 ();
 sg13g2_decap_8 FILLER_19_77 ();
 sg13g2_decap_8 FILLER_19_84 ();
 sg13g2_decap_8 FILLER_19_91 ();
 sg13g2_decap_8 FILLER_19_98 ();
 sg13g2_decap_8 FILLER_19_105 ();
 sg13g2_decap_8 FILLER_19_112 ();
 sg13g2_decap_8 FILLER_19_119 ();
 sg13g2_decap_8 FILLER_19_126 ();
 sg13g2_decap_8 FILLER_19_133 ();
 sg13g2_decap_4 FILLER_19_140 ();
 sg13g2_fill_1 FILLER_19_160 ();
 sg13g2_fill_1 FILLER_19_183 ();
 sg13g2_decap_8 FILLER_19_188 ();
 sg13g2_decap_8 FILLER_19_195 ();
 sg13g2_decap_8 FILLER_19_202 ();
 sg13g2_decap_8 FILLER_19_209 ();
 sg13g2_decap_8 FILLER_19_216 ();
 sg13g2_decap_8 FILLER_19_223 ();
 sg13g2_decap_8 FILLER_19_230 ();
 sg13g2_decap_8 FILLER_19_237 ();
 sg13g2_decap_8 FILLER_19_244 ();
 sg13g2_decap_8 FILLER_19_251 ();
 sg13g2_decap_8 FILLER_19_258 ();
 sg13g2_decap_8 FILLER_19_265 ();
 sg13g2_decap_8 FILLER_19_272 ();
 sg13g2_decap_8 FILLER_19_279 ();
 sg13g2_fill_2 FILLER_19_286 ();
 sg13g2_fill_1 FILLER_19_288 ();
 sg13g2_fill_2 FILLER_19_294 ();
 sg13g2_fill_2 FILLER_19_303 ();
 sg13g2_fill_1 FILLER_19_305 ();
 sg13g2_fill_2 FILLER_19_313 ();
 sg13g2_fill_2 FILLER_19_333 ();
 sg13g2_fill_1 FILLER_19_335 ();
 sg13g2_fill_2 FILLER_19_341 ();
 sg13g2_fill_1 FILLER_19_343 ();
 sg13g2_fill_2 FILLER_19_353 ();
 sg13g2_decap_8 FILLER_19_364 ();
 sg13g2_decap_8 FILLER_19_371 ();
 sg13g2_decap_8 FILLER_19_378 ();
 sg13g2_decap_8 FILLER_19_385 ();
 sg13g2_decap_8 FILLER_19_392 ();
 sg13g2_decap_8 FILLER_19_399 ();
 sg13g2_fill_2 FILLER_19_406 ();
 sg13g2_fill_1 FILLER_19_408 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_decap_8 FILLER_20_21 ();
 sg13g2_decap_8 FILLER_20_28 ();
 sg13g2_decap_8 FILLER_20_35 ();
 sg13g2_decap_8 FILLER_20_42 ();
 sg13g2_decap_8 FILLER_20_49 ();
 sg13g2_decap_8 FILLER_20_56 ();
 sg13g2_decap_8 FILLER_20_63 ();
 sg13g2_decap_8 FILLER_20_70 ();
 sg13g2_decap_8 FILLER_20_77 ();
 sg13g2_decap_8 FILLER_20_84 ();
 sg13g2_decap_8 FILLER_20_91 ();
 sg13g2_decap_8 FILLER_20_98 ();
 sg13g2_decap_8 FILLER_20_105 ();
 sg13g2_decap_8 FILLER_20_112 ();
 sg13g2_decap_8 FILLER_20_119 ();
 sg13g2_decap_4 FILLER_20_126 ();
 sg13g2_fill_1 FILLER_20_130 ();
 sg13g2_fill_1 FILLER_20_149 ();
 sg13g2_fill_1 FILLER_20_164 ();
 sg13g2_fill_2 FILLER_20_183 ();
 sg13g2_fill_1 FILLER_20_185 ();
 sg13g2_decap_8 FILLER_20_214 ();
 sg13g2_decap_8 FILLER_20_221 ();
 sg13g2_decap_8 FILLER_20_228 ();
 sg13g2_decap_8 FILLER_20_235 ();
 sg13g2_decap_8 FILLER_20_242 ();
 sg13g2_decap_8 FILLER_20_249 ();
 sg13g2_decap_8 FILLER_20_256 ();
 sg13g2_decap_8 FILLER_20_263 ();
 sg13g2_decap_8 FILLER_20_270 ();
 sg13g2_decap_8 FILLER_20_277 ();
 sg13g2_fill_2 FILLER_20_344 ();
 sg13g2_decap_8 FILLER_20_373 ();
 sg13g2_decap_8 FILLER_20_380 ();
 sg13g2_decap_8 FILLER_20_387 ();
 sg13g2_decap_8 FILLER_20_394 ();
 sg13g2_decap_8 FILLER_20_401 ();
 sg13g2_fill_1 FILLER_20_408 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_decap_8 FILLER_21_21 ();
 sg13g2_decap_8 FILLER_21_28 ();
 sg13g2_decap_8 FILLER_21_35 ();
 sg13g2_decap_8 FILLER_21_42 ();
 sg13g2_decap_8 FILLER_21_49 ();
 sg13g2_decap_8 FILLER_21_56 ();
 sg13g2_decap_8 FILLER_21_63 ();
 sg13g2_decap_8 FILLER_21_70 ();
 sg13g2_decap_8 FILLER_21_77 ();
 sg13g2_decap_8 FILLER_21_84 ();
 sg13g2_decap_8 FILLER_21_91 ();
 sg13g2_decap_8 FILLER_21_98 ();
 sg13g2_decap_8 FILLER_21_105 ();
 sg13g2_decap_8 FILLER_21_112 ();
 sg13g2_fill_2 FILLER_21_119 ();
 sg13g2_fill_1 FILLER_21_121 ();
 sg13g2_fill_1 FILLER_21_159 ();
 sg13g2_fill_2 FILLER_21_169 ();
 sg13g2_decap_8 FILLER_21_176 ();
 sg13g2_fill_2 FILLER_21_183 ();
 sg13g2_fill_1 FILLER_21_208 ();
 sg13g2_decap_8 FILLER_21_218 ();
 sg13g2_decap_8 FILLER_21_225 ();
 sg13g2_decap_8 FILLER_21_232 ();
 sg13g2_decap_8 FILLER_21_239 ();
 sg13g2_decap_8 FILLER_21_246 ();
 sg13g2_decap_8 FILLER_21_253 ();
 sg13g2_decap_8 FILLER_21_260 ();
 sg13g2_decap_4 FILLER_21_267 ();
 sg13g2_fill_1 FILLER_21_271 ();
 sg13g2_fill_2 FILLER_21_286 ();
 sg13g2_fill_1 FILLER_21_288 ();
 sg13g2_fill_1 FILLER_21_305 ();
 sg13g2_fill_2 FILLER_21_328 ();
 sg13g2_fill_1 FILLER_21_330 ();
 sg13g2_decap_8 FILLER_21_373 ();
 sg13g2_decap_8 FILLER_21_380 ();
 sg13g2_decap_8 FILLER_21_387 ();
 sg13g2_decap_8 FILLER_21_394 ();
 sg13g2_decap_8 FILLER_21_401 ();
 sg13g2_fill_1 FILLER_21_408 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_decap_8 FILLER_22_21 ();
 sg13g2_decap_8 FILLER_22_28 ();
 sg13g2_decap_8 FILLER_22_35 ();
 sg13g2_decap_8 FILLER_22_42 ();
 sg13g2_decap_8 FILLER_22_49 ();
 sg13g2_decap_8 FILLER_22_56 ();
 sg13g2_decap_8 FILLER_22_63 ();
 sg13g2_decap_8 FILLER_22_70 ();
 sg13g2_decap_8 FILLER_22_77 ();
 sg13g2_decap_8 FILLER_22_84 ();
 sg13g2_decap_8 FILLER_22_91 ();
 sg13g2_decap_8 FILLER_22_98 ();
 sg13g2_decap_8 FILLER_22_105 ();
 sg13g2_decap_8 FILLER_22_112 ();
 sg13g2_fill_2 FILLER_22_119 ();
 sg13g2_fill_2 FILLER_22_159 ();
 sg13g2_fill_2 FILLER_22_169 ();
 sg13g2_fill_1 FILLER_22_171 ();
 sg13g2_fill_1 FILLER_22_184 ();
 sg13g2_fill_1 FILLER_22_198 ();
 sg13g2_fill_1 FILLER_22_222 ();
 sg13g2_decap_8 FILLER_22_232 ();
 sg13g2_decap_8 FILLER_22_239 ();
 sg13g2_decap_8 FILLER_22_246 ();
 sg13g2_decap_8 FILLER_22_253 ();
 sg13g2_decap_4 FILLER_22_260 ();
 sg13g2_fill_1 FILLER_22_264 ();
 sg13g2_fill_2 FILLER_22_293 ();
 sg13g2_fill_2 FILLER_22_308 ();
 sg13g2_decap_8 FILLER_22_374 ();
 sg13g2_decap_8 FILLER_22_381 ();
 sg13g2_decap_8 FILLER_22_388 ();
 sg13g2_decap_8 FILLER_22_395 ();
 sg13g2_decap_8 FILLER_22_402 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_14 ();
 sg13g2_decap_8 FILLER_23_21 ();
 sg13g2_decap_8 FILLER_23_28 ();
 sg13g2_decap_8 FILLER_23_35 ();
 sg13g2_decap_8 FILLER_23_42 ();
 sg13g2_decap_8 FILLER_23_49 ();
 sg13g2_decap_8 FILLER_23_56 ();
 sg13g2_decap_8 FILLER_23_63 ();
 sg13g2_decap_8 FILLER_23_70 ();
 sg13g2_decap_8 FILLER_23_77 ();
 sg13g2_decap_8 FILLER_23_84 ();
 sg13g2_decap_8 FILLER_23_91 ();
 sg13g2_decap_8 FILLER_23_98 ();
 sg13g2_decap_8 FILLER_23_105 ();
 sg13g2_decap_8 FILLER_23_112 ();
 sg13g2_decap_8 FILLER_23_119 ();
 sg13g2_decap_4 FILLER_23_126 ();
 sg13g2_fill_1 FILLER_23_130 ();
 sg13g2_fill_2 FILLER_23_144 ();
 sg13g2_decap_8 FILLER_23_181 ();
 sg13g2_fill_2 FILLER_23_188 ();
 sg13g2_fill_1 FILLER_23_190 ();
 sg13g2_decap_4 FILLER_23_203 ();
 sg13g2_fill_1 FILLER_23_207 ();
 sg13g2_decap_8 FILLER_23_236 ();
 sg13g2_decap_8 FILLER_23_243 ();
 sg13g2_decap_8 FILLER_23_250 ();
 sg13g2_decap_8 FILLER_23_257 ();
 sg13g2_decap_8 FILLER_23_264 ();
 sg13g2_decap_4 FILLER_23_271 ();
 sg13g2_fill_2 FILLER_23_283 ();
 sg13g2_fill_1 FILLER_23_285 ();
 sg13g2_fill_1 FILLER_23_300 ();
 sg13g2_decap_8 FILLER_23_356 ();
 sg13g2_decap_8 FILLER_23_363 ();
 sg13g2_decap_8 FILLER_23_370 ();
 sg13g2_decap_8 FILLER_23_377 ();
 sg13g2_decap_8 FILLER_23_384 ();
 sg13g2_decap_8 FILLER_23_391 ();
 sg13g2_decap_8 FILLER_23_398 ();
 sg13g2_decap_4 FILLER_23_405 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_14 ();
 sg13g2_decap_8 FILLER_24_21 ();
 sg13g2_decap_8 FILLER_24_28 ();
 sg13g2_decap_8 FILLER_24_35 ();
 sg13g2_decap_8 FILLER_24_42 ();
 sg13g2_decap_8 FILLER_24_49 ();
 sg13g2_decap_8 FILLER_24_56 ();
 sg13g2_decap_8 FILLER_24_63 ();
 sg13g2_decap_8 FILLER_24_70 ();
 sg13g2_decap_8 FILLER_24_77 ();
 sg13g2_decap_8 FILLER_24_84 ();
 sg13g2_decap_8 FILLER_24_91 ();
 sg13g2_decap_8 FILLER_24_98 ();
 sg13g2_decap_8 FILLER_24_105 ();
 sg13g2_decap_8 FILLER_24_112 ();
 sg13g2_decap_8 FILLER_24_119 ();
 sg13g2_decap_8 FILLER_24_126 ();
 sg13g2_fill_2 FILLER_24_133 ();
 sg13g2_fill_1 FILLER_24_135 ();
 sg13g2_fill_2 FILLER_24_141 ();
 sg13g2_fill_1 FILLER_24_143 ();
 sg13g2_fill_1 FILLER_24_156 ();
 sg13g2_decap_4 FILLER_24_162 ();
 sg13g2_fill_2 FILLER_24_166 ();
 sg13g2_fill_1 FILLER_24_174 ();
 sg13g2_fill_2 FILLER_24_193 ();
 sg13g2_decap_8 FILLER_24_238 ();
 sg13g2_decap_8 FILLER_24_245 ();
 sg13g2_decap_8 FILLER_24_252 ();
 sg13g2_decap_8 FILLER_24_259 ();
 sg13g2_decap_8 FILLER_24_266 ();
 sg13g2_decap_4 FILLER_24_273 ();
 sg13g2_fill_2 FILLER_24_288 ();
 sg13g2_fill_2 FILLER_24_298 ();
 sg13g2_decap_4 FILLER_24_326 ();
 sg13g2_fill_1 FILLER_24_330 ();
 sg13g2_decap_8 FILLER_24_348 ();
 sg13g2_decap_8 FILLER_24_355 ();
 sg13g2_decap_8 FILLER_24_362 ();
 sg13g2_decap_8 FILLER_24_369 ();
 sg13g2_decap_8 FILLER_24_376 ();
 sg13g2_decap_8 FILLER_24_383 ();
 sg13g2_decap_8 FILLER_24_390 ();
 sg13g2_decap_8 FILLER_24_397 ();
 sg13g2_decap_4 FILLER_24_404 ();
 sg13g2_fill_1 FILLER_24_408 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_decap_8 FILLER_25_14 ();
 sg13g2_decap_8 FILLER_25_21 ();
 sg13g2_decap_8 FILLER_25_28 ();
 sg13g2_decap_8 FILLER_25_35 ();
 sg13g2_decap_8 FILLER_25_42 ();
 sg13g2_decap_8 FILLER_25_49 ();
 sg13g2_decap_8 FILLER_25_56 ();
 sg13g2_decap_8 FILLER_25_63 ();
 sg13g2_decap_8 FILLER_25_70 ();
 sg13g2_decap_8 FILLER_25_77 ();
 sg13g2_decap_8 FILLER_25_84 ();
 sg13g2_decap_8 FILLER_25_91 ();
 sg13g2_decap_8 FILLER_25_98 ();
 sg13g2_decap_8 FILLER_25_105 ();
 sg13g2_decap_8 FILLER_25_112 ();
 sg13g2_decap_8 FILLER_25_119 ();
 sg13g2_decap_8 FILLER_25_126 ();
 sg13g2_decap_8 FILLER_25_133 ();
 sg13g2_decap_8 FILLER_25_159 ();
 sg13g2_fill_2 FILLER_25_166 ();
 sg13g2_decap_4 FILLER_25_191 ();
 sg13g2_fill_2 FILLER_25_195 ();
 sg13g2_fill_1 FILLER_25_205 ();
 sg13g2_decap_4 FILLER_25_219 ();
 sg13g2_decap_8 FILLER_25_232 ();
 sg13g2_decap_8 FILLER_25_239 ();
 sg13g2_decap_8 FILLER_25_246 ();
 sg13g2_decap_8 FILLER_25_253 ();
 sg13g2_decap_8 FILLER_25_260 ();
 sg13g2_decap_8 FILLER_25_267 ();
 sg13g2_decap_8 FILLER_25_274 ();
 sg13g2_decap_8 FILLER_25_281 ();
 sg13g2_fill_2 FILLER_25_288 ();
 sg13g2_decap_8 FILLER_25_294 ();
 sg13g2_decap_8 FILLER_25_301 ();
 sg13g2_decap_4 FILLER_25_308 ();
 sg13g2_fill_1 FILLER_25_312 ();
 sg13g2_decap_8 FILLER_25_349 ();
 sg13g2_decap_8 FILLER_25_356 ();
 sg13g2_decap_8 FILLER_25_363 ();
 sg13g2_decap_8 FILLER_25_370 ();
 sg13g2_decap_8 FILLER_25_377 ();
 sg13g2_decap_8 FILLER_25_384 ();
 sg13g2_decap_8 FILLER_25_391 ();
 sg13g2_decap_8 FILLER_25_398 ();
 sg13g2_decap_4 FILLER_25_405 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_14 ();
 sg13g2_decap_8 FILLER_26_21 ();
 sg13g2_decap_8 FILLER_26_28 ();
 sg13g2_decap_8 FILLER_26_35 ();
 sg13g2_decap_8 FILLER_26_42 ();
 sg13g2_decap_8 FILLER_26_49 ();
 sg13g2_decap_8 FILLER_26_56 ();
 sg13g2_decap_8 FILLER_26_63 ();
 sg13g2_decap_8 FILLER_26_70 ();
 sg13g2_decap_8 FILLER_26_77 ();
 sg13g2_decap_8 FILLER_26_84 ();
 sg13g2_decap_8 FILLER_26_91 ();
 sg13g2_decap_8 FILLER_26_98 ();
 sg13g2_decap_8 FILLER_26_105 ();
 sg13g2_decap_8 FILLER_26_112 ();
 sg13g2_decap_8 FILLER_26_119 ();
 sg13g2_decap_4 FILLER_26_131 ();
 sg13g2_fill_1 FILLER_26_150 ();
 sg13g2_decap_8 FILLER_26_164 ();
 sg13g2_decap_4 FILLER_26_171 ();
 sg13g2_fill_1 FILLER_26_188 ();
 sg13g2_fill_2 FILLER_26_202 ();
 sg13g2_decap_8 FILLER_26_213 ();
 sg13g2_fill_2 FILLER_26_220 ();
 sg13g2_decap_8 FILLER_26_231 ();
 sg13g2_decap_8 FILLER_26_238 ();
 sg13g2_decap_8 FILLER_26_245 ();
 sg13g2_decap_8 FILLER_26_252 ();
 sg13g2_decap_8 FILLER_26_259 ();
 sg13g2_decap_8 FILLER_26_266 ();
 sg13g2_fill_1 FILLER_26_273 ();
 sg13g2_fill_2 FILLER_26_303 ();
 sg13g2_decap_8 FILLER_26_333 ();
 sg13g2_fill_1 FILLER_26_340 ();
 sg13g2_decap_8 FILLER_26_354 ();
 sg13g2_decap_8 FILLER_26_361 ();
 sg13g2_decap_8 FILLER_26_368 ();
 sg13g2_decap_8 FILLER_26_375 ();
 sg13g2_decap_8 FILLER_26_382 ();
 sg13g2_decap_8 FILLER_26_389 ();
 sg13g2_decap_8 FILLER_26_396 ();
 sg13g2_decap_4 FILLER_26_403 ();
 sg13g2_fill_2 FILLER_26_407 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_14 ();
 sg13g2_decap_8 FILLER_27_21 ();
 sg13g2_decap_8 FILLER_27_28 ();
 sg13g2_decap_8 FILLER_27_35 ();
 sg13g2_decap_8 FILLER_27_42 ();
 sg13g2_decap_8 FILLER_27_49 ();
 sg13g2_decap_8 FILLER_27_56 ();
 sg13g2_decap_8 FILLER_27_63 ();
 sg13g2_decap_8 FILLER_27_70 ();
 sg13g2_decap_8 FILLER_27_77 ();
 sg13g2_decap_8 FILLER_27_84 ();
 sg13g2_decap_8 FILLER_27_91 ();
 sg13g2_decap_8 FILLER_27_98 ();
 sg13g2_decap_8 FILLER_27_105 ();
 sg13g2_decap_8 FILLER_27_112 ();
 sg13g2_decap_4 FILLER_27_165 ();
 sg13g2_fill_2 FILLER_27_169 ();
 sg13g2_fill_1 FILLER_27_206 ();
 sg13g2_decap_8 FILLER_27_235 ();
 sg13g2_decap_8 FILLER_27_242 ();
 sg13g2_decap_8 FILLER_27_249 ();
 sg13g2_decap_4 FILLER_27_256 ();
 sg13g2_fill_2 FILLER_27_260 ();
 sg13g2_fill_2 FILLER_27_301 ();
 sg13g2_fill_1 FILLER_27_344 ();
 sg13g2_decap_8 FILLER_27_371 ();
 sg13g2_decap_8 FILLER_27_378 ();
 sg13g2_decap_8 FILLER_27_385 ();
 sg13g2_decap_8 FILLER_27_392 ();
 sg13g2_decap_8 FILLER_27_399 ();
 sg13g2_fill_2 FILLER_27_406 ();
 sg13g2_fill_1 FILLER_27_408 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_decap_8 FILLER_28_14 ();
 sg13g2_decap_8 FILLER_28_21 ();
 sg13g2_decap_8 FILLER_28_28 ();
 sg13g2_decap_8 FILLER_28_35 ();
 sg13g2_decap_8 FILLER_28_42 ();
 sg13g2_decap_8 FILLER_28_49 ();
 sg13g2_decap_8 FILLER_28_56 ();
 sg13g2_decap_8 FILLER_28_63 ();
 sg13g2_decap_8 FILLER_28_70 ();
 sg13g2_decap_8 FILLER_28_77 ();
 sg13g2_decap_8 FILLER_28_84 ();
 sg13g2_decap_8 FILLER_28_91 ();
 sg13g2_decap_8 FILLER_28_98 ();
 sg13g2_decap_8 FILLER_28_105 ();
 sg13g2_decap_8 FILLER_28_112 ();
 sg13g2_decap_4 FILLER_28_119 ();
 sg13g2_fill_1 FILLER_28_123 ();
 sg13g2_decap_4 FILLER_28_152 ();
 sg13g2_fill_1 FILLER_28_156 ();
 sg13g2_decap_4 FILLER_28_173 ();
 sg13g2_fill_2 FILLER_28_177 ();
 sg13g2_decap_4 FILLER_28_191 ();
 sg13g2_fill_2 FILLER_28_225 ();
 sg13g2_decap_8 FILLER_28_240 ();
 sg13g2_decap_8 FILLER_28_247 ();
 sg13g2_decap_8 FILLER_28_254 ();
 sg13g2_decap_8 FILLER_28_261 ();
 sg13g2_decap_8 FILLER_28_268 ();
 sg13g2_fill_1 FILLER_28_288 ();
 sg13g2_fill_2 FILLER_28_325 ();
 sg13g2_decap_4 FILLER_28_354 ();
 sg13g2_fill_2 FILLER_28_358 ();
 sg13g2_decap_8 FILLER_28_373 ();
 sg13g2_decap_8 FILLER_28_380 ();
 sg13g2_decap_8 FILLER_28_387 ();
 sg13g2_decap_8 FILLER_28_394 ();
 sg13g2_decap_8 FILLER_28_401 ();
 sg13g2_fill_1 FILLER_28_408 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_decap_8 FILLER_29_14 ();
 sg13g2_decap_8 FILLER_29_21 ();
 sg13g2_decap_8 FILLER_29_28 ();
 sg13g2_decap_8 FILLER_29_35 ();
 sg13g2_decap_8 FILLER_29_42 ();
 sg13g2_decap_8 FILLER_29_49 ();
 sg13g2_decap_8 FILLER_29_56 ();
 sg13g2_decap_8 FILLER_29_63 ();
 sg13g2_decap_8 FILLER_29_70 ();
 sg13g2_decap_8 FILLER_29_77 ();
 sg13g2_decap_8 FILLER_29_84 ();
 sg13g2_decap_8 FILLER_29_91 ();
 sg13g2_decap_8 FILLER_29_98 ();
 sg13g2_decap_8 FILLER_29_105 ();
 sg13g2_decap_8 FILLER_29_112 ();
 sg13g2_fill_2 FILLER_29_119 ();
 sg13g2_fill_2 FILLER_29_131 ();
 sg13g2_fill_1 FILLER_29_146 ();
 sg13g2_fill_2 FILLER_29_151 ();
 sg13g2_fill_1 FILLER_29_153 ();
 sg13g2_decap_8 FILLER_29_170 ();
 sg13g2_decap_4 FILLER_29_177 ();
 sg13g2_decap_8 FILLER_29_189 ();
 sg13g2_decap_8 FILLER_29_196 ();
 sg13g2_decap_8 FILLER_29_203 ();
 sg13g2_fill_1 FILLER_29_210 ();
 sg13g2_decap_8 FILLER_29_215 ();
 sg13g2_decap_8 FILLER_29_222 ();
 sg13g2_decap_8 FILLER_29_229 ();
 sg13g2_decap_8 FILLER_29_236 ();
 sg13g2_decap_8 FILLER_29_243 ();
 sg13g2_fill_2 FILLER_29_250 ();
 sg13g2_fill_1 FILLER_29_252 ();
 sg13g2_decap_8 FILLER_29_266 ();
 sg13g2_decap_8 FILLER_29_273 ();
 sg13g2_fill_1 FILLER_29_280 ();
 sg13g2_decap_8 FILLER_29_302 ();
 sg13g2_decap_8 FILLER_29_309 ();
 sg13g2_decap_8 FILLER_29_316 ();
 sg13g2_decap_8 FILLER_29_323 ();
 sg13g2_fill_1 FILLER_29_348 ();
 sg13g2_decap_8 FILLER_29_390 ();
 sg13g2_decap_8 FILLER_29_397 ();
 sg13g2_decap_4 FILLER_29_404 ();
 sg13g2_fill_1 FILLER_29_408 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_14 ();
 sg13g2_decap_8 FILLER_30_21 ();
 sg13g2_decap_8 FILLER_30_28 ();
 sg13g2_decap_8 FILLER_30_35 ();
 sg13g2_decap_8 FILLER_30_42 ();
 sg13g2_decap_8 FILLER_30_49 ();
 sg13g2_decap_8 FILLER_30_56 ();
 sg13g2_decap_8 FILLER_30_63 ();
 sg13g2_decap_8 FILLER_30_70 ();
 sg13g2_decap_8 FILLER_30_77 ();
 sg13g2_decap_8 FILLER_30_84 ();
 sg13g2_decap_8 FILLER_30_91 ();
 sg13g2_decap_8 FILLER_30_98 ();
 sg13g2_decap_8 FILLER_30_105 ();
 sg13g2_decap_4 FILLER_30_112 ();
 sg13g2_fill_1 FILLER_30_125 ();
 sg13g2_fill_2 FILLER_30_149 ();
 sg13g2_decap_8 FILLER_30_173 ();
 sg13g2_decap_8 FILLER_30_200 ();
 sg13g2_decap_8 FILLER_30_207 ();
 sg13g2_decap_8 FILLER_30_214 ();
 sg13g2_fill_1 FILLER_30_221 ();
 sg13g2_decap_8 FILLER_30_231 ();
 sg13g2_fill_2 FILLER_30_238 ();
 sg13g2_decap_8 FILLER_30_253 ();
 sg13g2_decap_8 FILLER_30_260 ();
 sg13g2_decap_8 FILLER_30_267 ();
 sg13g2_decap_8 FILLER_30_274 ();
 sg13g2_decap_8 FILLER_30_294 ();
 sg13g2_decap_8 FILLER_30_301 ();
 sg13g2_decap_8 FILLER_30_308 ();
 sg13g2_decap_8 FILLER_30_315 ();
 sg13g2_decap_8 FILLER_30_322 ();
 sg13g2_decap_8 FILLER_30_329 ();
 sg13g2_decap_8 FILLER_30_336 ();
 sg13g2_fill_1 FILLER_30_348 ();
 sg13g2_decap_8 FILLER_30_359 ();
 sg13g2_decap_8 FILLER_30_366 ();
 sg13g2_decap_8 FILLER_30_377 ();
 sg13g2_decap_8 FILLER_30_384 ();
 sg13g2_decap_8 FILLER_30_391 ();
 sg13g2_decap_8 FILLER_30_398 ();
 sg13g2_decap_4 FILLER_30_405 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_decap_8 FILLER_31_14 ();
 sg13g2_decap_8 FILLER_31_21 ();
 sg13g2_decap_8 FILLER_31_28 ();
 sg13g2_decap_8 FILLER_31_35 ();
 sg13g2_decap_8 FILLER_31_42 ();
 sg13g2_decap_8 FILLER_31_49 ();
 sg13g2_decap_8 FILLER_31_56 ();
 sg13g2_decap_8 FILLER_31_63 ();
 sg13g2_decap_8 FILLER_31_70 ();
 sg13g2_decap_8 FILLER_31_77 ();
 sg13g2_decap_8 FILLER_31_84 ();
 sg13g2_decap_8 FILLER_31_91 ();
 sg13g2_decap_8 FILLER_31_98 ();
 sg13g2_decap_4 FILLER_31_105 ();
 sg13g2_fill_2 FILLER_31_156 ();
 sg13g2_decap_8 FILLER_31_254 ();
 sg13g2_decap_4 FILLER_31_261 ();
 sg13g2_decap_4 FILLER_31_298 ();
 sg13g2_fill_2 FILLER_31_302 ();
 sg13g2_decap_8 FILLER_31_308 ();
 sg13g2_decap_4 FILLER_31_315 ();
 sg13g2_fill_2 FILLER_31_340 ();
 sg13g2_decap_4 FILLER_31_360 ();
 sg13g2_fill_1 FILLER_31_377 ();
 sg13g2_decap_8 FILLER_31_391 ();
 sg13g2_decap_8 FILLER_31_398 ();
 sg13g2_decap_4 FILLER_31_405 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_decap_8 FILLER_32_14 ();
 sg13g2_decap_8 FILLER_32_21 ();
 sg13g2_decap_8 FILLER_32_28 ();
 sg13g2_decap_8 FILLER_32_35 ();
 sg13g2_decap_8 FILLER_32_42 ();
 sg13g2_decap_8 FILLER_32_49 ();
 sg13g2_decap_8 FILLER_32_56 ();
 sg13g2_decap_8 FILLER_32_63 ();
 sg13g2_decap_8 FILLER_32_70 ();
 sg13g2_decap_8 FILLER_32_77 ();
 sg13g2_decap_8 FILLER_32_84 ();
 sg13g2_decap_8 FILLER_32_91 ();
 sg13g2_decap_8 FILLER_32_98 ();
 sg13g2_decap_4 FILLER_32_105 ();
 sg13g2_fill_1 FILLER_32_136 ();
 sg13g2_fill_1 FILLER_32_163 ();
 sg13g2_decap_4 FILLER_32_182 ();
 sg13g2_fill_2 FILLER_32_186 ();
 sg13g2_fill_2 FILLER_32_196 ();
 sg13g2_fill_2 FILLER_32_224 ();
 sg13g2_fill_1 FILLER_32_226 ();
 sg13g2_decap_4 FILLER_32_255 ();
 sg13g2_decap_4 FILLER_32_272 ();
 sg13g2_decap_4 FILLER_32_338 ();
 sg13g2_fill_2 FILLER_32_342 ();
 sg13g2_fill_2 FILLER_32_383 ();
 sg13g2_fill_1 FILLER_32_385 ();
 sg13g2_decap_8 FILLER_32_399 ();
 sg13g2_fill_2 FILLER_32_406 ();
 sg13g2_fill_1 FILLER_32_408 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_decap_8 FILLER_33_14 ();
 sg13g2_decap_8 FILLER_33_21 ();
 sg13g2_decap_8 FILLER_33_28 ();
 sg13g2_decap_8 FILLER_33_35 ();
 sg13g2_decap_8 FILLER_33_42 ();
 sg13g2_decap_8 FILLER_33_49 ();
 sg13g2_decap_8 FILLER_33_56 ();
 sg13g2_decap_8 FILLER_33_63 ();
 sg13g2_decap_8 FILLER_33_70 ();
 sg13g2_decap_8 FILLER_33_77 ();
 sg13g2_decap_8 FILLER_33_84 ();
 sg13g2_decap_8 FILLER_33_91 ();
 sg13g2_decap_8 FILLER_33_98 ();
 sg13g2_decap_8 FILLER_33_105 ();
 sg13g2_decap_4 FILLER_33_112 ();
 sg13g2_fill_1 FILLER_33_125 ();
 sg13g2_fill_2 FILLER_33_150 ();
 sg13g2_fill_2 FILLER_33_157 ();
 sg13g2_fill_1 FILLER_33_172 ();
 sg13g2_fill_2 FILLER_33_178 ();
 sg13g2_decap_4 FILLER_33_216 ();
 sg13g2_fill_2 FILLER_33_338 ();
 sg13g2_fill_1 FILLER_33_340 ();
 sg13g2_decap_8 FILLER_33_353 ();
 sg13g2_decap_8 FILLER_33_360 ();
 sg13g2_decap_8 FILLER_33_381 ();
 sg13g2_decap_8 FILLER_33_388 ();
 sg13g2_decap_8 FILLER_33_395 ();
 sg13g2_decap_8 FILLER_33_402 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_8 FILLER_34_14 ();
 sg13g2_decap_8 FILLER_34_21 ();
 sg13g2_decap_8 FILLER_34_28 ();
 sg13g2_decap_8 FILLER_34_35 ();
 sg13g2_decap_8 FILLER_34_42 ();
 sg13g2_decap_8 FILLER_34_49 ();
 sg13g2_decap_8 FILLER_34_56 ();
 sg13g2_decap_8 FILLER_34_63 ();
 sg13g2_decap_8 FILLER_34_70 ();
 sg13g2_decap_8 FILLER_34_77 ();
 sg13g2_decap_8 FILLER_34_84 ();
 sg13g2_decap_8 FILLER_34_91 ();
 sg13g2_decap_8 FILLER_34_98 ();
 sg13g2_decap_8 FILLER_34_105 ();
 sg13g2_decap_8 FILLER_34_112 ();
 sg13g2_fill_2 FILLER_34_119 ();
 sg13g2_fill_2 FILLER_34_126 ();
 sg13g2_fill_1 FILLER_34_128 ();
 sg13g2_decap_4 FILLER_34_148 ();
 sg13g2_fill_1 FILLER_34_152 ();
 sg13g2_decap_4 FILLER_34_170 ();
 sg13g2_fill_2 FILLER_34_174 ();
 sg13g2_fill_2 FILLER_34_185 ();
 sg13g2_fill_2 FILLER_34_190 ();
 sg13g2_fill_1 FILLER_34_192 ();
 sg13g2_fill_1 FILLER_34_207 ();
 sg13g2_fill_1 FILLER_34_217 ();
 sg13g2_fill_2 FILLER_34_223 ();
 sg13g2_fill_1 FILLER_34_225 ();
 sg13g2_fill_1 FILLER_34_231 ();
 sg13g2_fill_1 FILLER_34_241 ();
 sg13g2_decap_8 FILLER_34_260 ();
 sg13g2_decap_8 FILLER_34_267 ();
 sg13g2_decap_4 FILLER_34_274 ();
 sg13g2_fill_2 FILLER_34_278 ();
 sg13g2_fill_2 FILLER_34_346 ();
 sg13g2_fill_1 FILLER_34_348 ();
 sg13g2_decap_8 FILLER_34_354 ();
 sg13g2_decap_4 FILLER_34_361 ();
 sg13g2_decap_8 FILLER_34_379 ();
 sg13g2_decap_8 FILLER_34_386 ();
 sg13g2_decap_8 FILLER_34_393 ();
 sg13g2_decap_8 FILLER_34_400 ();
 sg13g2_fill_2 FILLER_34_407 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_decap_8 FILLER_35_21 ();
 sg13g2_decap_8 FILLER_35_28 ();
 sg13g2_decap_8 FILLER_35_35 ();
 sg13g2_decap_8 FILLER_35_42 ();
 sg13g2_decap_8 FILLER_35_49 ();
 sg13g2_decap_8 FILLER_35_56 ();
 sg13g2_decap_8 FILLER_35_63 ();
 sg13g2_decap_8 FILLER_35_70 ();
 sg13g2_decap_8 FILLER_35_77 ();
 sg13g2_decap_8 FILLER_35_84 ();
 sg13g2_decap_8 FILLER_35_91 ();
 sg13g2_decap_8 FILLER_35_98 ();
 sg13g2_decap_8 FILLER_35_105 ();
 sg13g2_decap_8 FILLER_35_112 ();
 sg13g2_decap_4 FILLER_35_119 ();
 sg13g2_fill_2 FILLER_35_149 ();
 sg13g2_decap_8 FILLER_35_165 ();
 sg13g2_decap_8 FILLER_35_186 ();
 sg13g2_decap_8 FILLER_35_193 ();
 sg13g2_fill_1 FILLER_35_200 ();
 sg13g2_decap_8 FILLER_35_205 ();
 sg13g2_fill_2 FILLER_35_212 ();
 sg13g2_fill_2 FILLER_35_218 ();
 sg13g2_fill_1 FILLER_35_220 ();
 sg13g2_decap_4 FILLER_35_249 ();
 sg13g2_fill_2 FILLER_35_253 ();
 sg13g2_fill_2 FILLER_35_304 ();
 sg13g2_fill_2 FILLER_35_340 ();
 sg13g2_fill_1 FILLER_35_382 ();
 sg13g2_decap_8 FILLER_35_388 ();
 sg13g2_decap_8 FILLER_35_395 ();
 sg13g2_decap_8 FILLER_35_402 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_8 FILLER_36_21 ();
 sg13g2_decap_8 FILLER_36_28 ();
 sg13g2_decap_8 FILLER_36_35 ();
 sg13g2_decap_8 FILLER_36_42 ();
 sg13g2_decap_8 FILLER_36_49 ();
 sg13g2_decap_8 FILLER_36_56 ();
 sg13g2_decap_8 FILLER_36_63 ();
 sg13g2_decap_8 FILLER_36_70 ();
 sg13g2_decap_8 FILLER_36_77 ();
 sg13g2_decap_8 FILLER_36_84 ();
 sg13g2_decap_8 FILLER_36_91 ();
 sg13g2_decap_8 FILLER_36_98 ();
 sg13g2_decap_8 FILLER_36_105 ();
 sg13g2_fill_1 FILLER_36_112 ();
 sg13g2_fill_2 FILLER_36_140 ();
 sg13g2_fill_1 FILLER_36_157 ();
 sg13g2_fill_1 FILLER_36_171 ();
 sg13g2_fill_2 FILLER_36_205 ();
 sg13g2_fill_1 FILLER_36_207 ();
 sg13g2_decap_4 FILLER_36_252 ();
 sg13g2_fill_2 FILLER_36_256 ();
 sg13g2_fill_2 FILLER_36_286 ();
 sg13g2_fill_1 FILLER_36_288 ();
 sg13g2_fill_2 FILLER_36_333 ();
 sg13g2_decap_8 FILLER_36_400 ();
 sg13g2_fill_2 FILLER_36_407 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_decap_8 FILLER_37_28 ();
 sg13g2_decap_8 FILLER_37_35 ();
 sg13g2_decap_8 FILLER_37_42 ();
 sg13g2_decap_8 FILLER_37_49 ();
 sg13g2_decap_8 FILLER_37_56 ();
 sg13g2_decap_8 FILLER_37_63 ();
 sg13g2_decap_8 FILLER_37_70 ();
 sg13g2_decap_8 FILLER_37_77 ();
 sg13g2_decap_8 FILLER_37_84 ();
 sg13g2_decap_8 FILLER_37_91 ();
 sg13g2_decap_8 FILLER_37_98 ();
 sg13g2_decap_8 FILLER_37_105 ();
 sg13g2_decap_4 FILLER_37_112 ();
 sg13g2_fill_1 FILLER_37_143 ();
 sg13g2_decap_4 FILLER_37_153 ();
 sg13g2_decap_8 FILLER_37_171 ();
 sg13g2_decap_8 FILLER_37_182 ();
 sg13g2_fill_2 FILLER_37_189 ();
 sg13g2_fill_2 FILLER_37_200 ();
 sg13g2_decap_8 FILLER_37_247 ();
 sg13g2_decap_8 FILLER_37_254 ();
 sg13g2_decap_4 FILLER_37_261 ();
 sg13g2_fill_1 FILLER_37_265 ();
 sg13g2_fill_1 FILLER_37_272 ();
 sg13g2_fill_2 FILLER_37_291 ();
 sg13g2_fill_1 FILLER_37_293 ();
 sg13g2_fill_1 FILLER_37_330 ();
 sg13g2_fill_2 FILLER_37_349 ();
 sg13g2_fill_1 FILLER_37_351 ();
 sg13g2_decap_4 FILLER_37_357 ();
 sg13g2_fill_2 FILLER_37_365 ();
 sg13g2_decap_8 FILLER_37_390 ();
 sg13g2_decap_8 FILLER_37_397 ();
 sg13g2_decap_4 FILLER_37_404 ();
 sg13g2_fill_1 FILLER_37_408 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_decap_8 FILLER_38_35 ();
 sg13g2_decap_8 FILLER_38_42 ();
 sg13g2_decap_8 FILLER_38_49 ();
 sg13g2_decap_8 FILLER_38_56 ();
 sg13g2_decap_8 FILLER_38_63 ();
 sg13g2_decap_8 FILLER_38_70 ();
 sg13g2_decap_8 FILLER_38_77 ();
 sg13g2_decap_8 FILLER_38_84 ();
 sg13g2_decap_8 FILLER_38_91 ();
 sg13g2_decap_8 FILLER_38_98 ();
 sg13g2_decap_8 FILLER_38_105 ();
 sg13g2_decap_8 FILLER_38_112 ();
 sg13g2_decap_8 FILLER_38_119 ();
 sg13g2_fill_2 FILLER_38_126 ();
 sg13g2_fill_2 FILLER_38_146 ();
 sg13g2_fill_2 FILLER_38_166 ();
 sg13g2_decap_4 FILLER_38_187 ();
 sg13g2_fill_1 FILLER_38_224 ();
 sg13g2_fill_2 FILLER_38_231 ();
 sg13g2_fill_2 FILLER_38_249 ();
 sg13g2_fill_1 FILLER_38_251 ();
 sg13g2_fill_2 FILLER_38_283 ();
 sg13g2_decap_8 FILLER_38_348 ();
 sg13g2_fill_1 FILLER_38_355 ();
 sg13g2_decap_4 FILLER_38_360 ();
 sg13g2_fill_1 FILLER_38_364 ();
 sg13g2_fill_2 FILLER_38_369 ();
 sg13g2_fill_1 FILLER_38_371 ();
 sg13g2_fill_2 FILLER_38_382 ();
 sg13g2_fill_1 FILLER_38_384 ();
 sg13g2_decap_4 FILLER_38_403 ();
 sg13g2_fill_2 FILLER_38_407 ();
 sg13g2_decap_8 FILLER_39_0 ();
 sg13g2_decap_8 FILLER_39_7 ();
 sg13g2_decap_8 FILLER_39_14 ();
 sg13g2_decap_8 FILLER_39_21 ();
 sg13g2_decap_8 FILLER_39_28 ();
 sg13g2_decap_8 FILLER_39_35 ();
 sg13g2_decap_8 FILLER_39_42 ();
 sg13g2_decap_8 FILLER_39_49 ();
 sg13g2_decap_8 FILLER_39_56 ();
 sg13g2_decap_8 FILLER_39_63 ();
 sg13g2_decap_8 FILLER_39_70 ();
 sg13g2_decap_8 FILLER_39_77 ();
 sg13g2_decap_8 FILLER_39_84 ();
 sg13g2_decap_8 FILLER_39_91 ();
 sg13g2_decap_8 FILLER_39_98 ();
 sg13g2_decap_8 FILLER_39_105 ();
 sg13g2_decap_8 FILLER_39_112 ();
 sg13g2_fill_2 FILLER_39_119 ();
 sg13g2_decap_8 FILLER_39_125 ();
 sg13g2_fill_1 FILLER_39_199 ();
 sg13g2_decap_8 FILLER_39_222 ();
 sg13g2_decap_4 FILLER_39_233 ();
 sg13g2_decap_8 FILLER_39_241 ();
 sg13g2_decap_8 FILLER_39_248 ();
 sg13g2_decap_8 FILLER_39_255 ();
 sg13g2_fill_1 FILLER_39_262 ();
 sg13g2_fill_2 FILLER_39_272 ();
 sg13g2_fill_1 FILLER_39_274 ();
 sg13g2_decap_8 FILLER_39_284 ();
 sg13g2_fill_2 FILLER_39_291 ();
 sg13g2_decap_8 FILLER_39_302 ();
 sg13g2_decap_8 FILLER_39_309 ();
 sg13g2_decap_8 FILLER_39_316 ();
 sg13g2_fill_1 FILLER_39_323 ();
 sg13g2_decap_8 FILLER_39_328 ();
 sg13g2_decap_8 FILLER_39_335 ();
 sg13g2_fill_2 FILLER_39_342 ();
 sg13g2_decap_8 FILLER_39_373 ();
 sg13g2_fill_2 FILLER_39_380 ();
 sg13g2_fill_1 FILLER_39_382 ();
 sg13g2_decap_8 FILLER_39_388 ();
 sg13g2_decap_8 FILLER_39_395 ();
 sg13g2_decap_8 FILLER_39_402 ();
 sg13g2_decap_8 FILLER_40_0 ();
 sg13g2_decap_8 FILLER_40_7 ();
 sg13g2_decap_8 FILLER_40_14 ();
 sg13g2_decap_8 FILLER_40_21 ();
 sg13g2_decap_8 FILLER_40_28 ();
 sg13g2_decap_8 FILLER_40_35 ();
 sg13g2_decap_8 FILLER_40_42 ();
 sg13g2_decap_8 FILLER_40_49 ();
 sg13g2_decap_8 FILLER_40_56 ();
 sg13g2_decap_8 FILLER_40_63 ();
 sg13g2_decap_8 FILLER_40_70 ();
 sg13g2_decap_8 FILLER_40_77 ();
 sg13g2_decap_8 FILLER_40_84 ();
 sg13g2_decap_8 FILLER_40_91 ();
 sg13g2_fill_1 FILLER_40_98 ();
 sg13g2_fill_2 FILLER_40_136 ();
 sg13g2_fill_1 FILLER_40_138 ();
 sg13g2_fill_2 FILLER_40_160 ();
 sg13g2_decap_4 FILLER_40_207 ();
 sg13g2_fill_1 FILLER_40_211 ();
 sg13g2_decap_4 FILLER_40_217 ();
 sg13g2_decap_8 FILLER_40_254 ();
 sg13g2_fill_2 FILLER_40_261 ();
 sg13g2_fill_1 FILLER_40_263 ();
 sg13g2_fill_2 FILLER_40_279 ();
 sg13g2_fill_1 FILLER_40_281 ();
 sg13g2_fill_2 FILLER_40_292 ();
 sg13g2_fill_2 FILLER_40_312 ();
 sg13g2_fill_2 FILLER_40_319 ();
 sg13g2_fill_1 FILLER_40_321 ();
 sg13g2_decap_4 FILLER_40_330 ();
 sg13g2_fill_1 FILLER_40_379 ();
 sg13g2_decap_8 FILLER_40_384 ();
 sg13g2_decap_8 FILLER_40_391 ();
 sg13g2_decap_8 FILLER_40_398 ();
 sg13g2_decap_4 FILLER_40_405 ();
 sg13g2_decap_8 FILLER_41_0 ();
 sg13g2_decap_8 FILLER_41_7 ();
 sg13g2_decap_8 FILLER_41_14 ();
 sg13g2_decap_8 FILLER_41_21 ();
 sg13g2_decap_8 FILLER_41_28 ();
 sg13g2_decap_8 FILLER_41_35 ();
 sg13g2_decap_8 FILLER_41_42 ();
 sg13g2_decap_8 FILLER_41_49 ();
 sg13g2_decap_8 FILLER_41_56 ();
 sg13g2_decap_8 FILLER_41_63 ();
 sg13g2_decap_8 FILLER_41_70 ();
 sg13g2_decap_8 FILLER_41_77 ();
 sg13g2_decap_8 FILLER_41_84 ();
 sg13g2_decap_8 FILLER_41_91 ();
 sg13g2_fill_2 FILLER_41_98 ();
 sg13g2_fill_2 FILLER_41_132 ();
 sg13g2_fill_2 FILLER_41_229 ();
 sg13g2_decap_8 FILLER_41_249 ();
 sg13g2_decap_4 FILLER_41_256 ();
 sg13g2_fill_2 FILLER_41_260 ();
 sg13g2_fill_2 FILLER_41_275 ();
 sg13g2_fill_1 FILLER_41_277 ();
 sg13g2_fill_2 FILLER_41_316 ();
 sg13g2_fill_2 FILLER_41_341 ();
 sg13g2_fill_1 FILLER_41_343 ();
 sg13g2_fill_1 FILLER_41_349 ();
 sg13g2_decap_8 FILLER_41_354 ();
 sg13g2_fill_2 FILLER_41_361 ();
 sg13g2_fill_1 FILLER_41_382 ();
 sg13g2_decap_8 FILLER_41_393 ();
 sg13g2_decap_8 FILLER_41_400 ();
 sg13g2_fill_2 FILLER_41_407 ();
 sg13g2_decap_8 FILLER_42_0 ();
 sg13g2_decap_8 FILLER_42_7 ();
 sg13g2_decap_8 FILLER_42_14 ();
 sg13g2_decap_8 FILLER_42_21 ();
 sg13g2_decap_8 FILLER_42_28 ();
 sg13g2_decap_8 FILLER_42_35 ();
 sg13g2_decap_8 FILLER_42_42 ();
 sg13g2_decap_8 FILLER_42_49 ();
 sg13g2_decap_8 FILLER_42_56 ();
 sg13g2_decap_8 FILLER_42_63 ();
 sg13g2_decap_8 FILLER_42_70 ();
 sg13g2_decap_8 FILLER_42_77 ();
 sg13g2_decap_8 FILLER_42_84 ();
 sg13g2_decap_8 FILLER_42_91 ();
 sg13g2_decap_8 FILLER_42_98 ();
 sg13g2_fill_2 FILLER_42_105 ();
 sg13g2_decap_8 FILLER_42_135 ();
 sg13g2_fill_2 FILLER_42_142 ();
 sg13g2_fill_2 FILLER_42_148 ();
 sg13g2_fill_1 FILLER_42_150 ();
 sg13g2_fill_1 FILLER_42_164 ();
 sg13g2_fill_2 FILLER_42_191 ();
 sg13g2_fill_2 FILLER_42_206 ();
 sg13g2_fill_1 FILLER_42_208 ();
 sg13g2_fill_2 FILLER_42_228 ();
 sg13g2_fill_1 FILLER_42_230 ();
 sg13g2_fill_1 FILLER_42_248 ();
 sg13g2_fill_2 FILLER_42_262 ();
 sg13g2_fill_1 FILLER_42_264 ();
 sg13g2_fill_1 FILLER_42_288 ();
 sg13g2_fill_2 FILLER_42_329 ();
 sg13g2_fill_2 FILLER_42_368 ();
 sg13g2_fill_1 FILLER_42_370 ();
 sg13g2_decap_4 FILLER_42_384 ();
 sg13g2_decap_8 FILLER_42_402 ();
 sg13g2_decap_8 FILLER_43_0 ();
 sg13g2_decap_8 FILLER_43_7 ();
 sg13g2_decap_8 FILLER_43_14 ();
 sg13g2_decap_8 FILLER_43_21 ();
 sg13g2_decap_8 FILLER_43_28 ();
 sg13g2_decap_8 FILLER_43_35 ();
 sg13g2_decap_8 FILLER_43_42 ();
 sg13g2_decap_8 FILLER_43_49 ();
 sg13g2_decap_8 FILLER_43_56 ();
 sg13g2_decap_8 FILLER_43_63 ();
 sg13g2_decap_8 FILLER_43_70 ();
 sg13g2_decap_8 FILLER_43_77 ();
 sg13g2_decap_8 FILLER_43_84 ();
 sg13g2_decap_8 FILLER_43_91 ();
 sg13g2_decap_8 FILLER_43_98 ();
 sg13g2_decap_8 FILLER_43_105 ();
 sg13g2_fill_2 FILLER_43_112 ();
 sg13g2_fill_1 FILLER_43_114 ();
 sg13g2_decap_4 FILLER_43_134 ();
 sg13g2_fill_2 FILLER_43_138 ();
 sg13g2_decap_8 FILLER_43_167 ();
 sg13g2_decap_8 FILLER_43_174 ();
 sg13g2_fill_2 FILLER_43_213 ();
 sg13g2_fill_1 FILLER_43_215 ();
 sg13g2_decap_4 FILLER_43_238 ();
 sg13g2_fill_2 FILLER_43_242 ();
 sg13g2_fill_2 FILLER_43_288 ();
 sg13g2_decap_4 FILLER_43_306 ();
 sg13g2_fill_2 FILLER_43_310 ();
 sg13g2_fill_2 FILLER_43_319 ();
 sg13g2_fill_1 FILLER_43_321 ();
 sg13g2_fill_2 FILLER_43_327 ();
 sg13g2_fill_1 FILLER_43_345 ();
 sg13g2_fill_1 FILLER_43_366 ();
 sg13g2_decap_4 FILLER_43_373 ();
 sg13g2_fill_1 FILLER_43_377 ();
 sg13g2_fill_2 FILLER_43_406 ();
 sg13g2_fill_1 FILLER_43_408 ();
 sg13g2_decap_8 FILLER_44_0 ();
 sg13g2_decap_8 FILLER_44_7 ();
 sg13g2_decap_8 FILLER_44_14 ();
 sg13g2_decap_8 FILLER_44_21 ();
 sg13g2_decap_8 FILLER_44_28 ();
 sg13g2_decap_8 FILLER_44_35 ();
 sg13g2_decap_8 FILLER_44_42 ();
 sg13g2_decap_8 FILLER_44_49 ();
 sg13g2_decap_8 FILLER_44_56 ();
 sg13g2_decap_8 FILLER_44_63 ();
 sg13g2_decap_8 FILLER_44_70 ();
 sg13g2_decap_8 FILLER_44_77 ();
 sg13g2_decap_8 FILLER_44_84 ();
 sg13g2_decap_8 FILLER_44_91 ();
 sg13g2_decap_8 FILLER_44_98 ();
 sg13g2_fill_1 FILLER_44_105 ();
 sg13g2_fill_1 FILLER_44_129 ();
 sg13g2_fill_1 FILLER_44_166 ();
 sg13g2_fill_1 FILLER_44_177 ();
 sg13g2_fill_1 FILLER_44_183 ();
 sg13g2_fill_2 FILLER_44_207 ();
 sg13g2_fill_1 FILLER_44_209 ();
 sg13g2_decap_8 FILLER_44_243 ();
 sg13g2_decap_8 FILLER_44_250 ();
 sg13g2_decap_4 FILLER_44_257 ();
 sg13g2_fill_1 FILLER_44_261 ();
 sg13g2_decap_4 FILLER_44_268 ();
 sg13g2_fill_2 FILLER_44_281 ();
 sg13g2_fill_1 FILLER_44_283 ();
 sg13g2_decap_4 FILLER_44_298 ();
 sg13g2_decap_8 FILLER_44_306 ();
 sg13g2_decap_8 FILLER_44_313 ();
 sg13g2_decap_8 FILLER_44_320 ();
 sg13g2_fill_2 FILLER_44_327 ();
 sg13g2_fill_1 FILLER_44_329 ();
 sg13g2_fill_2 FILLER_44_334 ();
 sg13g2_fill_1 FILLER_44_336 ();
 sg13g2_decap_8 FILLER_44_351 ();
 sg13g2_fill_1 FILLER_44_361 ();
 sg13g2_decap_8 FILLER_44_367 ();
 sg13g2_fill_2 FILLER_44_374 ();
 sg13g2_fill_1 FILLER_44_376 ();
 sg13g2_decap_8 FILLER_44_380 ();
 sg13g2_fill_1 FILLER_44_387 ();
 sg13g2_decap_8 FILLER_44_402 ();
 sg13g2_decap_8 FILLER_45_0 ();
 sg13g2_decap_8 FILLER_45_7 ();
 sg13g2_decap_8 FILLER_45_14 ();
 sg13g2_decap_8 FILLER_45_21 ();
 sg13g2_decap_8 FILLER_45_28 ();
 sg13g2_decap_8 FILLER_45_35 ();
 sg13g2_decap_8 FILLER_45_42 ();
 sg13g2_decap_8 FILLER_45_49 ();
 sg13g2_decap_8 FILLER_45_56 ();
 sg13g2_decap_8 FILLER_45_63 ();
 sg13g2_decap_8 FILLER_45_70 ();
 sg13g2_decap_8 FILLER_45_77 ();
 sg13g2_decap_8 FILLER_45_84 ();
 sg13g2_decap_4 FILLER_45_91 ();
 sg13g2_fill_1 FILLER_45_95 ();
 sg13g2_fill_2 FILLER_45_155 ();
 sg13g2_decap_4 FILLER_45_211 ();
 sg13g2_fill_2 FILLER_45_215 ();
 sg13g2_decap_8 FILLER_45_221 ();
 sg13g2_decap_8 FILLER_45_232 ();
 sg13g2_fill_1 FILLER_45_239 ();
 sg13g2_decap_8 FILLER_45_244 ();
 sg13g2_decap_4 FILLER_45_251 ();
 sg13g2_fill_2 FILLER_45_255 ();
 sg13g2_fill_2 FILLER_45_262 ();
 sg13g2_decap_8 FILLER_45_280 ();
 sg13g2_decap_8 FILLER_45_287 ();
 sg13g2_fill_2 FILLER_45_294 ();
 sg13g2_decap_8 FILLER_45_301 ();
 sg13g2_decap_8 FILLER_45_308 ();
 sg13g2_decap_8 FILLER_45_315 ();
 sg13g2_decap_8 FILLER_45_322 ();
 sg13g2_decap_8 FILLER_45_329 ();
 sg13g2_fill_2 FILLER_45_341 ();
 sg13g2_decap_4 FILLER_45_365 ();
 sg13g2_fill_2 FILLER_45_369 ();
 sg13g2_decap_4 FILLER_45_376 ();
 sg13g2_fill_1 FILLER_45_408 ();
 sg13g2_decap_8 FILLER_46_0 ();
 sg13g2_decap_8 FILLER_46_7 ();
 sg13g2_decap_8 FILLER_46_14 ();
 sg13g2_decap_8 FILLER_46_21 ();
 sg13g2_decap_8 FILLER_46_28 ();
 sg13g2_decap_8 FILLER_46_35 ();
 sg13g2_decap_8 FILLER_46_42 ();
 sg13g2_decap_8 FILLER_46_49 ();
 sg13g2_decap_8 FILLER_46_56 ();
 sg13g2_decap_8 FILLER_46_63 ();
 sg13g2_decap_8 FILLER_46_70 ();
 sg13g2_decap_8 FILLER_46_77 ();
 sg13g2_decap_8 FILLER_46_84 ();
 sg13g2_decap_8 FILLER_46_91 ();
 sg13g2_decap_8 FILLER_46_98 ();
 sg13g2_decap_8 FILLER_46_105 ();
 sg13g2_fill_1 FILLER_46_112 ();
 sg13g2_fill_1 FILLER_46_164 ();
 sg13g2_fill_2 FILLER_46_212 ();
 sg13g2_fill_1 FILLER_46_242 ();
 sg13g2_fill_1 FILLER_46_261 ();
 sg13g2_fill_2 FILLER_46_288 ();
 sg13g2_decap_8 FILLER_46_303 ();
 sg13g2_fill_2 FILLER_46_310 ();
 sg13g2_fill_2 FILLER_46_343 ();
 sg13g2_fill_1 FILLER_46_345 ();
 sg13g2_fill_2 FILLER_46_363 ();
 sg13g2_decap_8 FILLER_46_383 ();
 sg13g2_decap_8 FILLER_46_390 ();
 sg13g2_decap_8 FILLER_46_397 ();
 sg13g2_decap_4 FILLER_46_404 ();
 sg13g2_fill_1 FILLER_46_408 ();
 sg13g2_decap_8 FILLER_47_0 ();
 sg13g2_decap_8 FILLER_47_7 ();
 sg13g2_decap_8 FILLER_47_14 ();
 sg13g2_decap_8 FILLER_47_21 ();
 sg13g2_decap_8 FILLER_47_28 ();
 sg13g2_decap_8 FILLER_47_35 ();
 sg13g2_decap_8 FILLER_47_42 ();
 sg13g2_decap_8 FILLER_47_49 ();
 sg13g2_decap_8 FILLER_47_56 ();
 sg13g2_decap_8 FILLER_47_63 ();
 sg13g2_decap_8 FILLER_47_70 ();
 sg13g2_decap_8 FILLER_47_77 ();
 sg13g2_decap_8 FILLER_47_84 ();
 sg13g2_decap_8 FILLER_47_91 ();
 sg13g2_decap_8 FILLER_47_98 ();
 sg13g2_decap_8 FILLER_47_105 ();
 sg13g2_decap_8 FILLER_47_112 ();
 sg13g2_decap_8 FILLER_47_123 ();
 sg13g2_decap_8 FILLER_47_130 ();
 sg13g2_fill_1 FILLER_47_137 ();
 sg13g2_fill_2 FILLER_47_153 ();
 sg13g2_fill_2 FILLER_47_160 ();
 sg13g2_fill_1 FILLER_47_162 ();
 sg13g2_decap_4 FILLER_47_167 ();
 sg13g2_fill_1 FILLER_47_171 ();
 sg13g2_fill_2 FILLER_47_176 ();
 sg13g2_decap_8 FILLER_47_201 ();
 sg13g2_decap_4 FILLER_47_208 ();
 sg13g2_fill_1 FILLER_47_212 ();
 sg13g2_decap_4 FILLER_47_218 ();
 sg13g2_fill_1 FILLER_47_240 ();
 sg13g2_fill_2 FILLER_47_304 ();
 sg13g2_fill_2 FILLER_47_341 ();
 sg13g2_fill_1 FILLER_47_374 ();
 sg13g2_decap_4 FILLER_47_403 ();
 sg13g2_fill_2 FILLER_47_407 ();
 sg13g2_decap_8 FILLER_48_0 ();
 sg13g2_decap_8 FILLER_48_7 ();
 sg13g2_decap_8 FILLER_48_14 ();
 sg13g2_decap_8 FILLER_48_21 ();
 sg13g2_decap_8 FILLER_48_28 ();
 sg13g2_decap_8 FILLER_48_35 ();
 sg13g2_decap_8 FILLER_48_42 ();
 sg13g2_decap_8 FILLER_48_49 ();
 sg13g2_decap_8 FILLER_48_56 ();
 sg13g2_decap_8 FILLER_48_63 ();
 sg13g2_decap_8 FILLER_48_70 ();
 sg13g2_decap_8 FILLER_48_77 ();
 sg13g2_decap_8 FILLER_48_84 ();
 sg13g2_decap_8 FILLER_48_91 ();
 sg13g2_decap_8 FILLER_48_98 ();
 sg13g2_decap_8 FILLER_48_105 ();
 sg13g2_fill_1 FILLER_48_112 ();
 sg13g2_decap_8 FILLER_48_132 ();
 sg13g2_fill_2 FILLER_48_139 ();
 sg13g2_fill_1 FILLER_48_141 ();
 sg13g2_decap_4 FILLER_48_146 ();
 sg13g2_fill_2 FILLER_48_150 ();
 sg13g2_decap_8 FILLER_48_161 ();
 sg13g2_decap_8 FILLER_48_168 ();
 sg13g2_decap_8 FILLER_48_175 ();
 sg13g2_decap_4 FILLER_48_182 ();
 sg13g2_fill_2 FILLER_48_186 ();
 sg13g2_decap_8 FILLER_48_201 ();
 sg13g2_fill_1 FILLER_48_224 ();
 sg13g2_fill_1 FILLER_48_233 ();
 sg13g2_decap_8 FILLER_48_247 ();
 sg13g2_decap_8 FILLER_48_254 ();
 sg13g2_fill_2 FILLER_48_261 ();
 sg13g2_fill_1 FILLER_48_263 ();
 sg13g2_fill_2 FILLER_48_281 ();
 sg13g2_fill_1 FILLER_48_283 ();
 sg13g2_fill_2 FILLER_48_304 ();
 sg13g2_fill_1 FILLER_48_306 ();
 sg13g2_decap_8 FILLER_48_344 ();
 sg13g2_fill_2 FILLER_48_351 ();
 sg13g2_fill_1 FILLER_48_353 ();
 sg13g2_fill_2 FILLER_48_364 ();
 sg13g2_decap_8 FILLER_49_0 ();
 sg13g2_decap_8 FILLER_49_7 ();
 sg13g2_decap_8 FILLER_49_14 ();
 sg13g2_decap_8 FILLER_49_21 ();
 sg13g2_decap_8 FILLER_49_28 ();
 sg13g2_decap_8 FILLER_49_35 ();
 sg13g2_decap_8 FILLER_49_42 ();
 sg13g2_decap_8 FILLER_49_49 ();
 sg13g2_decap_8 FILLER_49_56 ();
 sg13g2_decap_8 FILLER_49_63 ();
 sg13g2_decap_8 FILLER_49_70 ();
 sg13g2_decap_8 FILLER_49_77 ();
 sg13g2_decap_8 FILLER_49_84 ();
 sg13g2_decap_8 FILLER_49_91 ();
 sg13g2_decap_4 FILLER_49_98 ();
 sg13g2_fill_1 FILLER_49_102 ();
 sg13g2_fill_2 FILLER_49_130 ();
 sg13g2_fill_1 FILLER_49_132 ();
 sg13g2_fill_2 FILLER_49_143 ();
 sg13g2_fill_1 FILLER_49_145 ();
 sg13g2_decap_8 FILLER_49_164 ();
 sg13g2_decap_8 FILLER_49_171 ();
 sg13g2_fill_2 FILLER_49_178 ();
 sg13g2_fill_2 FILLER_49_185 ();
 sg13g2_decap_4 FILLER_49_197 ();
 sg13g2_fill_1 FILLER_49_201 ();
 sg13g2_decap_8 FILLER_49_242 ();
 sg13g2_decap_8 FILLER_49_249 ();
 sg13g2_decap_8 FILLER_49_256 ();
 sg13g2_fill_2 FILLER_49_273 ();
 sg13g2_fill_2 FILLER_49_285 ();
 sg13g2_fill_1 FILLER_49_287 ();
 sg13g2_fill_1 FILLER_49_293 ();
 sg13g2_decap_8 FILLER_49_299 ();
 sg13g2_decap_4 FILLER_49_306 ();
 sg13g2_fill_1 FILLER_49_310 ();
 sg13g2_decap_8 FILLER_49_324 ();
 sg13g2_decap_8 FILLER_49_331 ();
 sg13g2_decap_8 FILLER_49_338 ();
 sg13g2_decap_4 FILLER_49_345 ();
 sg13g2_fill_2 FILLER_49_359 ();
 sg13g2_fill_1 FILLER_49_361 ();
 sg13g2_fill_2 FILLER_49_406 ();
 sg13g2_fill_1 FILLER_49_408 ();
 sg13g2_decap_8 FILLER_50_0 ();
 sg13g2_decap_8 FILLER_50_7 ();
 sg13g2_decap_8 FILLER_50_14 ();
 sg13g2_decap_8 FILLER_50_21 ();
 sg13g2_decap_8 FILLER_50_28 ();
 sg13g2_decap_8 FILLER_50_35 ();
 sg13g2_decap_8 FILLER_50_42 ();
 sg13g2_decap_8 FILLER_50_49 ();
 sg13g2_decap_8 FILLER_50_56 ();
 sg13g2_decap_8 FILLER_50_63 ();
 sg13g2_decap_8 FILLER_50_70 ();
 sg13g2_decap_8 FILLER_50_77 ();
 sg13g2_decap_8 FILLER_50_84 ();
 sg13g2_decap_4 FILLER_50_91 ();
 sg13g2_fill_2 FILLER_50_95 ();
 sg13g2_fill_2 FILLER_50_124 ();
 sg13g2_fill_1 FILLER_50_126 ();
 sg13g2_fill_2 FILLER_50_160 ();
 sg13g2_fill_1 FILLER_50_162 ();
 sg13g2_decap_4 FILLER_50_193 ();
 sg13g2_fill_2 FILLER_50_197 ();
 sg13g2_decap_8 FILLER_50_224 ();
 sg13g2_decap_8 FILLER_50_231 ();
 sg13g2_decap_8 FILLER_50_238 ();
 sg13g2_decap_8 FILLER_50_245 ();
 sg13g2_decap_8 FILLER_50_252 ();
 sg13g2_decap_4 FILLER_50_259 ();
 sg13g2_fill_1 FILLER_50_263 ();
 sg13g2_fill_2 FILLER_50_290 ();
 sg13g2_decap_8 FILLER_50_298 ();
 sg13g2_decap_8 FILLER_50_305 ();
 sg13g2_fill_2 FILLER_50_312 ();
 sg13g2_fill_1 FILLER_50_314 ();
 sg13g2_decap_8 FILLER_50_325 ();
 sg13g2_fill_2 FILLER_50_338 ();
 sg13g2_fill_2 FILLER_50_375 ();
 sg13g2_decap_8 FILLER_51_0 ();
 sg13g2_decap_8 FILLER_51_7 ();
 sg13g2_decap_8 FILLER_51_14 ();
 sg13g2_decap_8 FILLER_51_21 ();
 sg13g2_decap_8 FILLER_51_28 ();
 sg13g2_decap_8 FILLER_51_35 ();
 sg13g2_decap_8 FILLER_51_42 ();
 sg13g2_decap_8 FILLER_51_49 ();
 sg13g2_decap_8 FILLER_51_56 ();
 sg13g2_decap_8 FILLER_51_63 ();
 sg13g2_decap_8 FILLER_51_70 ();
 sg13g2_decap_8 FILLER_51_77 ();
 sg13g2_decap_8 FILLER_51_84 ();
 sg13g2_decap_8 FILLER_51_91 ();
 sg13g2_decap_8 FILLER_51_98 ();
 sg13g2_fill_1 FILLER_51_105 ();
 sg13g2_fill_1 FILLER_51_130 ();
 sg13g2_fill_2 FILLER_51_145 ();
 sg13g2_fill_2 FILLER_51_163 ();
 sg13g2_fill_2 FILLER_51_219 ();
 sg13g2_decap_4 FILLER_51_304 ();
 sg13g2_fill_1 FILLER_51_308 ();
 sg13g2_fill_2 FILLER_51_338 ();
 sg13g2_fill_1 FILLER_51_340 ();
 sg13g2_fill_1 FILLER_51_359 ();
 sg13g2_decap_4 FILLER_51_385 ();
 sg13g2_fill_2 FILLER_51_389 ();
 sg13g2_decap_4 FILLER_51_404 ();
 sg13g2_fill_1 FILLER_51_408 ();
 sg13g2_decap_8 FILLER_52_0 ();
 sg13g2_decap_8 FILLER_52_7 ();
 sg13g2_decap_8 FILLER_52_14 ();
 sg13g2_decap_8 FILLER_52_21 ();
 sg13g2_decap_8 FILLER_52_28 ();
 sg13g2_decap_8 FILLER_52_35 ();
 sg13g2_decap_8 FILLER_52_42 ();
 sg13g2_decap_8 FILLER_52_49 ();
 sg13g2_decap_8 FILLER_52_56 ();
 sg13g2_decap_8 FILLER_52_63 ();
 sg13g2_decap_8 FILLER_52_70 ();
 sg13g2_decap_8 FILLER_52_77 ();
 sg13g2_decap_8 FILLER_52_84 ();
 sg13g2_decap_8 FILLER_52_91 ();
 sg13g2_decap_4 FILLER_52_98 ();
 sg13g2_decap_8 FILLER_52_184 ();
 sg13g2_fill_2 FILLER_52_191 ();
 sg13g2_fill_1 FILLER_52_193 ();
 sg13g2_decap_8 FILLER_52_213 ();
 sg13g2_decap_4 FILLER_52_220 ();
 sg13g2_decap_8 FILLER_52_227 ();
 sg13g2_fill_2 FILLER_52_234 ();
 sg13g2_fill_1 FILLER_52_236 ();
 sg13g2_decap_8 FILLER_52_249 ();
 sg13g2_fill_2 FILLER_52_256 ();
 sg13g2_fill_1 FILLER_52_258 ();
 sg13g2_fill_1 FILLER_52_273 ();
 sg13g2_fill_1 FILLER_52_294 ();
 sg13g2_fill_2 FILLER_52_310 ();
 sg13g2_fill_1 FILLER_52_317 ();
 sg13g2_fill_2 FILLER_52_349 ();
 sg13g2_fill_1 FILLER_52_356 ();
 sg13g2_fill_2 FILLER_52_399 ();
 sg13g2_fill_1 FILLER_52_401 ();
 sg13g2_fill_2 FILLER_52_407 ();
 sg13g2_decap_8 FILLER_53_0 ();
 sg13g2_decap_8 FILLER_53_7 ();
 sg13g2_decap_8 FILLER_53_14 ();
 sg13g2_decap_8 FILLER_53_21 ();
 sg13g2_decap_8 FILLER_53_28 ();
 sg13g2_decap_8 FILLER_53_35 ();
 sg13g2_decap_8 FILLER_53_42 ();
 sg13g2_decap_8 FILLER_53_49 ();
 sg13g2_decap_8 FILLER_53_56 ();
 sg13g2_decap_8 FILLER_53_63 ();
 sg13g2_decap_8 FILLER_53_70 ();
 sg13g2_decap_8 FILLER_53_77 ();
 sg13g2_decap_8 FILLER_53_84 ();
 sg13g2_decap_4 FILLER_53_91 ();
 sg13g2_fill_1 FILLER_53_95 ();
 sg13g2_fill_2 FILLER_53_133 ();
 sg13g2_decap_4 FILLER_53_149 ();
 sg13g2_fill_1 FILLER_53_153 ();
 sg13g2_decap_4 FILLER_53_171 ();
 sg13g2_fill_2 FILLER_53_175 ();
 sg13g2_decap_8 FILLER_53_181 ();
 sg13g2_fill_2 FILLER_53_188 ();
 sg13g2_decap_8 FILLER_53_208 ();
 sg13g2_fill_1 FILLER_53_215 ();
 sg13g2_fill_2 FILLER_53_220 ();
 sg13g2_decap_4 FILLER_53_246 ();
 sg13g2_decap_4 FILLER_53_259 ();
 sg13g2_fill_2 FILLER_53_263 ();
 sg13g2_fill_2 FILLER_53_284 ();
 sg13g2_fill_2 FILLER_53_292 ();
 sg13g2_fill_1 FILLER_53_294 ();
 sg13g2_decap_8 FILLER_53_300 ();
 sg13g2_decap_8 FILLER_53_307 ();
 sg13g2_decap_8 FILLER_53_314 ();
 sg13g2_fill_1 FILLER_53_321 ();
 sg13g2_decap_8 FILLER_53_334 ();
 sg13g2_fill_1 FILLER_53_341 ();
 sg13g2_decap_8 FILLER_53_346 ();
 sg13g2_decap_8 FILLER_53_353 ();
 sg13g2_decap_8 FILLER_53_360 ();
 sg13g2_decap_4 FILLER_53_367 ();
 sg13g2_fill_2 FILLER_53_371 ();
 sg13g2_fill_2 FILLER_53_392 ();
 sg13g2_fill_1 FILLER_53_394 ();
 sg13g2_fill_2 FILLER_53_407 ();
 sg13g2_decap_8 FILLER_54_0 ();
 sg13g2_decap_8 FILLER_54_7 ();
 sg13g2_decap_8 FILLER_54_14 ();
 sg13g2_decap_8 FILLER_54_21 ();
 sg13g2_decap_8 FILLER_54_28 ();
 sg13g2_decap_8 FILLER_54_35 ();
 sg13g2_decap_8 FILLER_54_42 ();
 sg13g2_decap_8 FILLER_54_49 ();
 sg13g2_decap_8 FILLER_54_56 ();
 sg13g2_decap_8 FILLER_54_63 ();
 sg13g2_decap_8 FILLER_54_70 ();
 sg13g2_decap_8 FILLER_54_77 ();
 sg13g2_decap_8 FILLER_54_84 ();
 sg13g2_decap_8 FILLER_54_91 ();
 sg13g2_decap_8 FILLER_54_98 ();
 sg13g2_decap_8 FILLER_54_105 ();
 sg13g2_decap_4 FILLER_54_117 ();
 sg13g2_fill_1 FILLER_54_162 ();
 sg13g2_fill_1 FILLER_54_183 ();
 sg13g2_decap_4 FILLER_54_191 ();
 sg13g2_fill_1 FILLER_54_195 ();
 sg13g2_fill_2 FILLER_54_212 ();
 sg13g2_fill_1 FILLER_54_261 ();
 sg13g2_decap_8 FILLER_54_274 ();
 sg13g2_decap_8 FILLER_54_281 ();
 sg13g2_decap_8 FILLER_54_288 ();
 sg13g2_decap_4 FILLER_54_295 ();
 sg13g2_decap_8 FILLER_54_309 ();
 sg13g2_fill_1 FILLER_54_322 ();
 sg13g2_fill_1 FILLER_54_330 ();
 sg13g2_decap_8 FILLER_54_340 ();
 sg13g2_decap_8 FILLER_54_347 ();
 sg13g2_decap_4 FILLER_54_354 ();
 sg13g2_fill_2 FILLER_54_368 ();
 sg13g2_fill_1 FILLER_54_370 ();
 sg13g2_fill_2 FILLER_54_381 ();
 sg13g2_fill_1 FILLER_54_383 ();
 sg13g2_fill_2 FILLER_54_407 ();
 sg13g2_decap_8 FILLER_55_0 ();
 sg13g2_decap_8 FILLER_55_7 ();
 sg13g2_decap_8 FILLER_55_14 ();
 sg13g2_decap_8 FILLER_55_21 ();
 sg13g2_decap_8 FILLER_55_28 ();
 sg13g2_decap_8 FILLER_55_35 ();
 sg13g2_decap_8 FILLER_55_42 ();
 sg13g2_decap_8 FILLER_55_49 ();
 sg13g2_decap_8 FILLER_55_56 ();
 sg13g2_decap_8 FILLER_55_63 ();
 sg13g2_decap_8 FILLER_55_70 ();
 sg13g2_decap_8 FILLER_55_77 ();
 sg13g2_decap_8 FILLER_55_84 ();
 sg13g2_decap_8 FILLER_55_91 ();
 sg13g2_decap_8 FILLER_55_98 ();
 sg13g2_decap_8 FILLER_55_105 ();
 sg13g2_decap_8 FILLER_55_112 ();
 sg13g2_fill_1 FILLER_55_119 ();
 sg13g2_fill_2 FILLER_55_125 ();
 sg13g2_fill_2 FILLER_55_194 ();
 sg13g2_decap_4 FILLER_55_265 ();
 sg13g2_fill_2 FILLER_55_269 ();
 sg13g2_decap_8 FILLER_55_275 ();
 sg13g2_decap_4 FILLER_55_282 ();
 sg13g2_fill_2 FILLER_55_286 ();
 sg13g2_decap_4 FILLER_55_293 ();
 sg13g2_fill_2 FILLER_55_302 ();
 sg13g2_decap_4 FILLER_55_309 ();
 sg13g2_fill_2 FILLER_55_313 ();
 sg13g2_decap_8 FILLER_55_324 ();
 sg13g2_decap_8 FILLER_55_331 ();
 sg13g2_decap_4 FILLER_55_343 ();
 sg13g2_fill_1 FILLER_55_367 ();
 sg13g2_fill_2 FILLER_55_381 ();
 sg13g2_decap_8 FILLER_56_0 ();
 sg13g2_decap_8 FILLER_56_7 ();
 sg13g2_decap_8 FILLER_56_14 ();
 sg13g2_decap_8 FILLER_56_21 ();
 sg13g2_decap_8 FILLER_56_28 ();
 sg13g2_decap_8 FILLER_56_35 ();
 sg13g2_decap_8 FILLER_56_42 ();
 sg13g2_decap_8 FILLER_56_49 ();
 sg13g2_decap_8 FILLER_56_56 ();
 sg13g2_decap_8 FILLER_56_63 ();
 sg13g2_decap_8 FILLER_56_70 ();
 sg13g2_decap_8 FILLER_56_77 ();
 sg13g2_decap_8 FILLER_56_84 ();
 sg13g2_decap_8 FILLER_56_91 ();
 sg13g2_decap_8 FILLER_56_98 ();
 sg13g2_decap_8 FILLER_56_105 ();
 sg13g2_decap_8 FILLER_56_112 ();
 sg13g2_decap_4 FILLER_56_119 ();
 sg13g2_fill_2 FILLER_56_123 ();
 sg13g2_fill_1 FILLER_56_142 ();
 sg13g2_fill_2 FILLER_56_175 ();
 sg13g2_decap_8 FILLER_56_198 ();
 sg13g2_decap_8 FILLER_56_205 ();
 sg13g2_fill_2 FILLER_56_212 ();
 sg13g2_decap_4 FILLER_56_219 ();
 sg13g2_fill_2 FILLER_56_236 ();
 sg13g2_decap_4 FILLER_56_256 ();
 sg13g2_fill_1 FILLER_56_315 ();
 sg13g2_decap_4 FILLER_56_325 ();
 sg13g2_fill_2 FILLER_56_329 ();
 sg13g2_fill_2 FILLER_56_344 ();
 sg13g2_fill_1 FILLER_56_346 ();
 sg13g2_decap_4 FILLER_56_371 ();
 sg13g2_fill_2 FILLER_56_375 ();
 sg13g2_decap_8 FILLER_56_401 ();
 sg13g2_fill_1 FILLER_56_408 ();
 sg13g2_decap_8 FILLER_57_0 ();
 sg13g2_decap_8 FILLER_57_7 ();
 sg13g2_decap_8 FILLER_57_14 ();
 sg13g2_decap_8 FILLER_57_21 ();
 sg13g2_decap_8 FILLER_57_28 ();
 sg13g2_decap_8 FILLER_57_35 ();
 sg13g2_decap_8 FILLER_57_42 ();
 sg13g2_decap_8 FILLER_57_49 ();
 sg13g2_decap_8 FILLER_57_56 ();
 sg13g2_decap_8 FILLER_57_63 ();
 sg13g2_decap_8 FILLER_57_70 ();
 sg13g2_decap_8 FILLER_57_77 ();
 sg13g2_decap_8 FILLER_57_84 ();
 sg13g2_decap_4 FILLER_57_91 ();
 sg13g2_fill_2 FILLER_57_95 ();
 sg13g2_fill_2 FILLER_57_128 ();
 sg13g2_fill_1 FILLER_57_130 ();
 sg13g2_fill_2 FILLER_57_136 ();
 sg13g2_fill_1 FILLER_57_138 ();
 sg13g2_decap_8 FILLER_57_147 ();
 sg13g2_fill_2 FILLER_57_170 ();
 sg13g2_decap_4 FILLER_57_190 ();
 sg13g2_fill_2 FILLER_57_215 ();
 sg13g2_fill_2 FILLER_57_249 ();
 sg13g2_decap_8 FILLER_57_256 ();
 sg13g2_fill_1 FILLER_57_263 ();
 sg13g2_decap_8 FILLER_57_267 ();
 sg13g2_decap_8 FILLER_57_274 ();
 sg13g2_decap_8 FILLER_57_281 ();
 sg13g2_decap_8 FILLER_57_315 ();
 sg13g2_fill_1 FILLER_57_322 ();
 sg13g2_decap_8 FILLER_57_370 ();
 sg13g2_decap_8 FILLER_57_377 ();
 sg13g2_decap_8 FILLER_57_384 ();
 sg13g2_decap_8 FILLER_57_391 ();
 sg13g2_decap_8 FILLER_57_398 ();
 sg13g2_decap_4 FILLER_57_405 ();
 sg13g2_decap_8 FILLER_58_0 ();
 sg13g2_decap_8 FILLER_58_7 ();
 sg13g2_decap_8 FILLER_58_14 ();
 sg13g2_decap_8 FILLER_58_21 ();
 sg13g2_decap_8 FILLER_58_28 ();
 sg13g2_decap_8 FILLER_58_35 ();
 sg13g2_decap_8 FILLER_58_42 ();
 sg13g2_decap_8 FILLER_58_49 ();
 sg13g2_decap_8 FILLER_58_56 ();
 sg13g2_decap_8 FILLER_58_63 ();
 sg13g2_decap_8 FILLER_58_70 ();
 sg13g2_decap_8 FILLER_58_77 ();
 sg13g2_decap_8 FILLER_58_84 ();
 sg13g2_decap_4 FILLER_58_91 ();
 sg13g2_fill_2 FILLER_58_146 ();
 sg13g2_decap_8 FILLER_58_155 ();
 sg13g2_decap_8 FILLER_58_162 ();
 sg13g2_fill_2 FILLER_58_169 ();
 sg13g2_fill_1 FILLER_58_171 ();
 sg13g2_decap_4 FILLER_58_177 ();
 sg13g2_decap_8 FILLER_58_184 ();
 sg13g2_decap_8 FILLER_58_191 ();
 sg13g2_decap_4 FILLER_58_198 ();
 sg13g2_fill_1 FILLER_58_237 ();
 sg13g2_decap_4 FILLER_58_260 ();
 sg13g2_decap_8 FILLER_58_267 ();
 sg13g2_fill_1 FILLER_58_327 ();
 sg13g2_fill_1 FILLER_58_332 ();
 sg13g2_decap_4 FILLER_58_339 ();
 sg13g2_fill_1 FILLER_58_343 ();
 sg13g2_decap_8 FILLER_58_357 ();
 sg13g2_decap_8 FILLER_58_364 ();
 sg13g2_decap_8 FILLER_58_371 ();
 sg13g2_decap_8 FILLER_58_378 ();
 sg13g2_fill_2 FILLER_58_385 ();
 sg13g2_decap_8 FILLER_58_400 ();
 sg13g2_fill_2 FILLER_58_407 ();
 sg13g2_decap_8 FILLER_59_0 ();
 sg13g2_decap_8 FILLER_59_7 ();
 sg13g2_decap_8 FILLER_59_14 ();
 sg13g2_decap_8 FILLER_59_21 ();
 sg13g2_decap_8 FILLER_59_28 ();
 sg13g2_decap_8 FILLER_59_35 ();
 sg13g2_decap_8 FILLER_59_42 ();
 sg13g2_decap_8 FILLER_59_49 ();
 sg13g2_decap_8 FILLER_59_56 ();
 sg13g2_decap_8 FILLER_59_63 ();
 sg13g2_decap_8 FILLER_59_70 ();
 sg13g2_decap_8 FILLER_59_77 ();
 sg13g2_decap_8 FILLER_59_84 ();
 sg13g2_decap_8 FILLER_59_91 ();
 sg13g2_fill_1 FILLER_59_98 ();
 sg13g2_fill_2 FILLER_59_104 ();
 sg13g2_fill_1 FILLER_59_106 ();
 sg13g2_fill_2 FILLER_59_148 ();
 sg13g2_fill_2 FILLER_59_188 ();
 sg13g2_fill_1 FILLER_59_190 ();
 sg13g2_decap_8 FILLER_59_194 ();
 sg13g2_decap_8 FILLER_59_201 ();
 sg13g2_decap_4 FILLER_59_208 ();
 sg13g2_fill_1 FILLER_59_212 ();
 sg13g2_fill_1 FILLER_59_226 ();
 sg13g2_fill_2 FILLER_59_273 ();
 sg13g2_fill_1 FILLER_59_275 ();
 sg13g2_fill_1 FILLER_59_296 ();
 sg13g2_decap_8 FILLER_59_329 ();
 sg13g2_decap_8 FILLER_59_336 ();
 sg13g2_decap_4 FILLER_59_363 ();
 sg13g2_decap_8 FILLER_59_401 ();
 sg13g2_fill_1 FILLER_59_408 ();
 sg13g2_decap_8 FILLER_60_0 ();
 sg13g2_decap_8 FILLER_60_7 ();
 sg13g2_decap_8 FILLER_60_14 ();
 sg13g2_decap_8 FILLER_60_21 ();
 sg13g2_decap_8 FILLER_60_28 ();
 sg13g2_decap_8 FILLER_60_35 ();
 sg13g2_decap_8 FILLER_60_42 ();
 sg13g2_decap_8 FILLER_60_49 ();
 sg13g2_decap_8 FILLER_60_56 ();
 sg13g2_decap_8 FILLER_60_63 ();
 sg13g2_decap_8 FILLER_60_70 ();
 sg13g2_decap_8 FILLER_60_77 ();
 sg13g2_decap_8 FILLER_60_84 ();
 sg13g2_decap_8 FILLER_60_91 ();
 sg13g2_decap_8 FILLER_60_98 ();
 sg13g2_fill_2 FILLER_60_105 ();
 sg13g2_fill_1 FILLER_60_107 ();
 sg13g2_decap_4 FILLER_60_203 ();
 sg13g2_fill_1 FILLER_60_207 ();
 sg13g2_decap_8 FILLER_60_220 ();
 sg13g2_fill_1 FILLER_60_280 ();
 sg13g2_decap_4 FILLER_60_295 ();
 sg13g2_fill_2 FILLER_60_299 ();
 sg13g2_fill_1 FILLER_60_318 ();
 sg13g2_decap_8 FILLER_60_322 ();
 sg13g2_decap_8 FILLER_60_329 ();
 sg13g2_fill_2 FILLER_60_336 ();
 sg13g2_fill_1 FILLER_60_338 ();
 sg13g2_decap_8 FILLER_60_343 ();
 sg13g2_fill_2 FILLER_60_350 ();
 sg13g2_decap_4 FILLER_60_362 ();
 sg13g2_fill_1 FILLER_60_366 ();
 sg13g2_decap_4 FILLER_60_388 ();
 sg13g2_decap_4 FILLER_60_403 ();
 sg13g2_fill_2 FILLER_60_407 ();
 sg13g2_decap_8 FILLER_61_0 ();
 sg13g2_decap_8 FILLER_61_7 ();
 sg13g2_decap_8 FILLER_61_14 ();
 sg13g2_decap_8 FILLER_61_21 ();
 sg13g2_decap_8 FILLER_61_28 ();
 sg13g2_decap_8 FILLER_61_35 ();
 sg13g2_decap_8 FILLER_61_42 ();
 sg13g2_decap_8 FILLER_61_49 ();
 sg13g2_decap_8 FILLER_61_56 ();
 sg13g2_decap_8 FILLER_61_63 ();
 sg13g2_decap_8 FILLER_61_70 ();
 sg13g2_decap_8 FILLER_61_77 ();
 sg13g2_decap_8 FILLER_61_84 ();
 sg13g2_decap_4 FILLER_61_91 ();
 sg13g2_fill_2 FILLER_61_123 ();
 sg13g2_fill_1 FILLER_61_125 ();
 sg13g2_fill_2 FILLER_61_130 ();
 sg13g2_fill_1 FILLER_61_132 ();
 sg13g2_fill_1 FILLER_61_167 ();
 sg13g2_fill_1 FILLER_61_194 ();
 sg13g2_decap_4 FILLER_61_259 ();
 sg13g2_fill_1 FILLER_61_263 ();
 sg13g2_decap_4 FILLER_61_301 ();
 sg13g2_fill_1 FILLER_61_305 ();
 sg13g2_decap_8 FILLER_61_309 ();
 sg13g2_decap_8 FILLER_61_316 ();
 sg13g2_decap_8 FILLER_61_323 ();
 sg13g2_fill_2 FILLER_61_348 ();
 sg13g2_fill_1 FILLER_61_350 ();
 sg13g2_decap_8 FILLER_61_361 ();
 sg13g2_fill_2 FILLER_61_368 ();
 sg13g2_fill_1 FILLER_61_370 ();
 sg13g2_decap_4 FILLER_61_381 ();
 sg13g2_fill_1 FILLER_61_408 ();
 sg13g2_decap_8 FILLER_62_0 ();
 sg13g2_decap_8 FILLER_62_7 ();
 sg13g2_decap_8 FILLER_62_14 ();
 sg13g2_decap_8 FILLER_62_21 ();
 sg13g2_decap_8 FILLER_62_28 ();
 sg13g2_decap_8 FILLER_62_35 ();
 sg13g2_decap_8 FILLER_62_42 ();
 sg13g2_decap_8 FILLER_62_49 ();
 sg13g2_decap_8 FILLER_62_56 ();
 sg13g2_decap_8 FILLER_62_63 ();
 sg13g2_decap_8 FILLER_62_70 ();
 sg13g2_decap_8 FILLER_62_77 ();
 sg13g2_decap_8 FILLER_62_84 ();
 sg13g2_decap_8 FILLER_62_91 ();
 sg13g2_fill_1 FILLER_62_98 ();
 sg13g2_decap_8 FILLER_62_152 ();
 sg13g2_decap_8 FILLER_62_159 ();
 sg13g2_fill_2 FILLER_62_166 ();
 sg13g2_fill_2 FILLER_62_219 ();
 sg13g2_decap_8 FILLER_62_260 ();
 sg13g2_fill_1 FILLER_62_267 ();
 sg13g2_fill_1 FILLER_62_281 ();
 sg13g2_decap_4 FILLER_62_309 ();
 sg13g2_decap_4 FILLER_62_317 ();
 sg13g2_decap_4 FILLER_62_360 ();
 sg13g2_fill_1 FILLER_62_364 ();
 sg13g2_fill_2 FILLER_62_406 ();
 sg13g2_fill_1 FILLER_62_408 ();
 sg13g2_decap_8 FILLER_63_0 ();
 sg13g2_decap_8 FILLER_63_7 ();
 sg13g2_decap_8 FILLER_63_14 ();
 sg13g2_decap_8 FILLER_63_21 ();
 sg13g2_decap_8 FILLER_63_28 ();
 sg13g2_decap_8 FILLER_63_35 ();
 sg13g2_decap_8 FILLER_63_42 ();
 sg13g2_decap_8 FILLER_63_49 ();
 sg13g2_decap_8 FILLER_63_56 ();
 sg13g2_decap_8 FILLER_63_63 ();
 sg13g2_decap_8 FILLER_63_70 ();
 sg13g2_decap_8 FILLER_63_77 ();
 sg13g2_decap_8 FILLER_63_84 ();
 sg13g2_decap_8 FILLER_63_91 ();
 sg13g2_fill_2 FILLER_63_135 ();
 sg13g2_decap_8 FILLER_63_146 ();
 sg13g2_fill_2 FILLER_63_153 ();
 sg13g2_fill_1 FILLER_63_155 ();
 sg13g2_fill_2 FILLER_63_243 ();
 sg13g2_fill_1 FILLER_63_245 ();
 sg13g2_decap_8 FILLER_63_260 ();
 sg13g2_fill_2 FILLER_63_271 ();
 sg13g2_fill_1 FILLER_63_273 ();
 sg13g2_fill_1 FILLER_63_279 ();
 sg13g2_fill_2 FILLER_63_300 ();
 sg13g2_fill_2 FILLER_63_307 ();
 sg13g2_fill_1 FILLER_63_309 ();
 sg13g2_fill_2 FILLER_63_352 ();
 sg13g2_fill_1 FILLER_63_354 ();
 sg13g2_decap_8 FILLER_64_0 ();
 sg13g2_decap_8 FILLER_64_7 ();
 sg13g2_decap_8 FILLER_64_14 ();
 sg13g2_decap_8 FILLER_64_21 ();
 sg13g2_decap_8 FILLER_64_28 ();
 sg13g2_decap_8 FILLER_64_35 ();
 sg13g2_decap_8 FILLER_64_42 ();
 sg13g2_decap_8 FILLER_64_49 ();
 sg13g2_decap_8 FILLER_64_56 ();
 sg13g2_decap_8 FILLER_64_63 ();
 sg13g2_decap_8 FILLER_64_70 ();
 sg13g2_decap_8 FILLER_64_77 ();
 sg13g2_decap_8 FILLER_64_84 ();
 sg13g2_decap_8 FILLER_64_91 ();
 sg13g2_decap_8 FILLER_64_98 ();
 sg13g2_fill_2 FILLER_64_105 ();
 sg13g2_fill_1 FILLER_64_135 ();
 sg13g2_fill_2 FILLER_64_151 ();
 sg13g2_fill_1 FILLER_64_153 ();
 sg13g2_fill_2 FILLER_64_161 ();
 sg13g2_fill_1 FILLER_64_163 ();
 sg13g2_fill_2 FILLER_64_201 ();
 sg13g2_fill_1 FILLER_64_203 ();
 sg13g2_fill_1 FILLER_64_232 ();
 sg13g2_fill_2 FILLER_64_242 ();
 sg13g2_fill_1 FILLER_64_276 ();
 sg13g2_fill_2 FILLER_64_304 ();
 sg13g2_fill_2 FILLER_64_340 ();
 sg13g2_decap_4 FILLER_64_379 ();
 sg13g2_decap_8 FILLER_65_0 ();
 sg13g2_decap_8 FILLER_65_7 ();
 sg13g2_decap_8 FILLER_65_14 ();
 sg13g2_decap_8 FILLER_65_21 ();
 sg13g2_decap_8 FILLER_65_28 ();
 sg13g2_decap_8 FILLER_65_35 ();
 sg13g2_decap_8 FILLER_65_42 ();
 sg13g2_decap_8 FILLER_65_49 ();
 sg13g2_decap_8 FILLER_65_56 ();
 sg13g2_decap_8 FILLER_65_63 ();
 sg13g2_decap_8 FILLER_65_70 ();
 sg13g2_decap_8 FILLER_65_77 ();
 sg13g2_decap_4 FILLER_65_84 ();
 sg13g2_fill_2 FILLER_65_145 ();
 sg13g2_fill_1 FILLER_65_147 ();
 sg13g2_decap_8 FILLER_65_166 ();
 sg13g2_decap_8 FILLER_65_173 ();
 sg13g2_decap_4 FILLER_65_180 ();
 sg13g2_fill_2 FILLER_65_184 ();
 sg13g2_decap_4 FILLER_65_227 ();
 sg13g2_decap_4 FILLER_65_248 ();
 sg13g2_decap_4 FILLER_65_257 ();
 sg13g2_fill_1 FILLER_65_261 ();
 sg13g2_decap_4 FILLER_65_265 ();
 sg13g2_fill_2 FILLER_65_269 ();
 sg13g2_fill_1 FILLER_65_282 ();
 sg13g2_decap_4 FILLER_65_296 ();
 sg13g2_decap_8 FILLER_65_328 ();
 sg13g2_decap_8 FILLER_65_335 ();
 sg13g2_fill_2 FILLER_65_342 ();
 sg13g2_fill_1 FILLER_65_344 ();
 sg13g2_decap_4 FILLER_65_359 ();
 sg13g2_fill_2 FILLER_65_372 ();
 sg13g2_fill_2 FILLER_65_392 ();
 sg13g2_fill_1 FILLER_65_394 ();
 sg13g2_decap_8 FILLER_66_0 ();
 sg13g2_decap_8 FILLER_66_7 ();
 sg13g2_decap_8 FILLER_66_14 ();
 sg13g2_decap_8 FILLER_66_21 ();
 sg13g2_decap_8 FILLER_66_28 ();
 sg13g2_decap_8 FILLER_66_35 ();
 sg13g2_decap_8 FILLER_66_42 ();
 sg13g2_decap_8 FILLER_66_49 ();
 sg13g2_decap_8 FILLER_66_56 ();
 sg13g2_decap_8 FILLER_66_63 ();
 sg13g2_decap_8 FILLER_66_70 ();
 sg13g2_decap_8 FILLER_66_77 ();
 sg13g2_decap_8 FILLER_66_84 ();
 sg13g2_fill_2 FILLER_66_91 ();
 sg13g2_fill_2 FILLER_66_106 ();
 sg13g2_fill_1 FILLER_66_108 ();
 sg13g2_fill_2 FILLER_66_123 ();
 sg13g2_fill_1 FILLER_66_154 ();
 sg13g2_decap_8 FILLER_66_168 ();
 sg13g2_decap_8 FILLER_66_175 ();
 sg13g2_decap_8 FILLER_66_182 ();
 sg13g2_decap_4 FILLER_66_211 ();
 sg13g2_fill_2 FILLER_66_215 ();
 sg13g2_fill_2 FILLER_66_222 ();
 sg13g2_fill_1 FILLER_66_224 ();
 sg13g2_fill_2 FILLER_66_265 ();
 sg13g2_decap_4 FILLER_66_280 ();
 sg13g2_fill_2 FILLER_66_284 ();
 sg13g2_decap_8 FILLER_66_292 ();
 sg13g2_decap_4 FILLER_66_299 ();
 sg13g2_fill_2 FILLER_66_303 ();
 sg13g2_decap_8 FILLER_66_328 ();
 sg13g2_decap_4 FILLER_66_335 ();
 sg13g2_decap_8 FILLER_66_354 ();
 sg13g2_decap_8 FILLER_66_361 ();
 sg13g2_decap_8 FILLER_66_368 ();
 sg13g2_decap_8 FILLER_66_375 ();
 sg13g2_fill_1 FILLER_66_408 ();
 sg13g2_decap_8 FILLER_67_0 ();
 sg13g2_decap_8 FILLER_67_7 ();
 sg13g2_decap_8 FILLER_67_14 ();
 sg13g2_decap_8 FILLER_67_21 ();
 sg13g2_decap_8 FILLER_67_28 ();
 sg13g2_decap_8 FILLER_67_35 ();
 sg13g2_decap_8 FILLER_67_42 ();
 sg13g2_decap_8 FILLER_67_49 ();
 sg13g2_decap_8 FILLER_67_56 ();
 sg13g2_decap_8 FILLER_67_63 ();
 sg13g2_decap_8 FILLER_67_70 ();
 sg13g2_decap_8 FILLER_67_77 ();
 sg13g2_decap_8 FILLER_67_84 ();
 sg13g2_decap_4 FILLER_67_91 ();
 sg13g2_fill_1 FILLER_67_95 ();
 sg13g2_fill_1 FILLER_67_125 ();
 sg13g2_decap_8 FILLER_67_130 ();
 sg13g2_fill_1 FILLER_67_137 ();
 sg13g2_fill_2 FILLER_67_172 ();
 sg13g2_decap_8 FILLER_67_202 ();
 sg13g2_decap_8 FILLER_67_209 ();
 sg13g2_fill_2 FILLER_67_216 ();
 sg13g2_decap_4 FILLER_67_231 ();
 sg13g2_fill_1 FILLER_67_272 ();
 sg13g2_decap_4 FILLER_67_285 ();
 sg13g2_fill_1 FILLER_67_289 ();
 sg13g2_decap_4 FILLER_67_294 ();
 sg13g2_fill_1 FILLER_67_298 ();
 sg13g2_decap_8 FILLER_67_304 ();
 sg13g2_fill_2 FILLER_67_311 ();
 sg13g2_fill_2 FILLER_67_347 ();
 sg13g2_fill_1 FILLER_67_349 ();
 sg13g2_fill_2 FILLER_67_386 ();
 sg13g2_fill_1 FILLER_67_388 ();
 sg13g2_fill_2 FILLER_67_406 ();
 sg13g2_fill_1 FILLER_67_408 ();
 sg13g2_decap_8 FILLER_68_0 ();
 sg13g2_decap_8 FILLER_68_7 ();
 sg13g2_decap_8 FILLER_68_14 ();
 sg13g2_decap_8 FILLER_68_21 ();
 sg13g2_decap_8 FILLER_68_28 ();
 sg13g2_decap_8 FILLER_68_35 ();
 sg13g2_decap_8 FILLER_68_42 ();
 sg13g2_decap_8 FILLER_68_49 ();
 sg13g2_decap_8 FILLER_68_56 ();
 sg13g2_decap_8 FILLER_68_63 ();
 sg13g2_decap_8 FILLER_68_70 ();
 sg13g2_decap_8 FILLER_68_77 ();
 sg13g2_fill_2 FILLER_68_84 ();
 sg13g2_decap_8 FILLER_68_128 ();
 sg13g2_decap_8 FILLER_68_135 ();
 sg13g2_decap_8 FILLER_68_142 ();
 sg13g2_fill_1 FILLER_68_149 ();
 sg13g2_decap_8 FILLER_68_182 ();
 sg13g2_fill_2 FILLER_68_189 ();
 sg13g2_decap_8 FILLER_68_202 ();
 sg13g2_decap_4 FILLER_68_236 ();
 sg13g2_fill_2 FILLER_68_274 ();
 sg13g2_fill_1 FILLER_68_276 ();
 sg13g2_fill_1 FILLER_68_316 ();
 sg13g2_fill_1 FILLER_68_322 ();
 sg13g2_fill_2 FILLER_68_342 ();
 sg13g2_fill_2 FILLER_68_406 ();
 sg13g2_fill_1 FILLER_68_408 ();
 sg13g2_decap_8 FILLER_69_0 ();
 sg13g2_decap_8 FILLER_69_7 ();
 sg13g2_decap_8 FILLER_69_14 ();
 sg13g2_decap_8 FILLER_69_21 ();
 sg13g2_decap_8 FILLER_69_28 ();
 sg13g2_decap_8 FILLER_69_35 ();
 sg13g2_decap_8 FILLER_69_42 ();
 sg13g2_decap_8 FILLER_69_49 ();
 sg13g2_decap_8 FILLER_69_56 ();
 sg13g2_decap_8 FILLER_69_63 ();
 sg13g2_decap_8 FILLER_69_70 ();
 sg13g2_decap_8 FILLER_69_77 ();
 sg13g2_decap_8 FILLER_69_84 ();
 sg13g2_decap_4 FILLER_69_91 ();
 sg13g2_decap_4 FILLER_69_104 ();
 sg13g2_fill_2 FILLER_69_126 ();
 sg13g2_fill_1 FILLER_69_137 ();
 sg13g2_fill_2 FILLER_69_152 ();
 sg13g2_fill_1 FILLER_69_172 ();
 sg13g2_fill_1 FILLER_69_186 ();
 sg13g2_fill_2 FILLER_69_235 ();
 sg13g2_fill_2 FILLER_69_256 ();
 sg13g2_fill_2 FILLER_69_305 ();
 sg13g2_fill_1 FILLER_69_340 ();
 sg13g2_decap_8 FILLER_70_0 ();
 sg13g2_decap_8 FILLER_70_7 ();
 sg13g2_decap_8 FILLER_70_14 ();
 sg13g2_decap_8 FILLER_70_21 ();
 sg13g2_decap_8 FILLER_70_28 ();
 sg13g2_decap_8 FILLER_70_35 ();
 sg13g2_decap_8 FILLER_70_42 ();
 sg13g2_decap_8 FILLER_70_49 ();
 sg13g2_decap_8 FILLER_70_56 ();
 sg13g2_decap_8 FILLER_70_63 ();
 sg13g2_decap_8 FILLER_70_70 ();
 sg13g2_decap_8 FILLER_70_77 ();
 sg13g2_decap_8 FILLER_70_84 ();
 sg13g2_decap_8 FILLER_70_91 ();
 sg13g2_decap_4 FILLER_70_98 ();
 sg13g2_fill_2 FILLER_70_107 ();
 sg13g2_fill_1 FILLER_70_109 ();
 sg13g2_fill_2 FILLER_70_118 ();
 sg13g2_fill_2 FILLER_70_126 ();
 sg13g2_fill_1 FILLER_70_163 ();
 sg13g2_fill_2 FILLER_70_168 ();
 sg13g2_fill_2 FILLER_70_190 ();
 sg13g2_fill_1 FILLER_70_195 ();
 sg13g2_fill_2 FILLER_70_207 ();
 sg13g2_decap_4 FILLER_70_218 ();
 sg13g2_decap_4 FILLER_70_241 ();
 sg13g2_fill_2 FILLER_70_245 ();
 sg13g2_fill_2 FILLER_70_251 ();
 sg13g2_fill_1 FILLER_70_253 ();
 sg13g2_fill_1 FILLER_70_289 ();
 sg13g2_decap_8 FILLER_70_333 ();
 sg13g2_fill_2 FILLER_70_350 ();
 sg13g2_fill_1 FILLER_70_352 ();
 sg13g2_fill_2 FILLER_70_388 ();
 sg13g2_decap_8 FILLER_71_0 ();
 sg13g2_decap_8 FILLER_71_7 ();
 sg13g2_decap_8 FILLER_71_14 ();
 sg13g2_decap_8 FILLER_71_21 ();
 sg13g2_decap_8 FILLER_71_28 ();
 sg13g2_decap_8 FILLER_71_35 ();
 sg13g2_decap_8 FILLER_71_42 ();
 sg13g2_decap_8 FILLER_71_49 ();
 sg13g2_decap_8 FILLER_71_56 ();
 sg13g2_decap_8 FILLER_71_63 ();
 sg13g2_decap_8 FILLER_71_70 ();
 sg13g2_decap_8 FILLER_71_77 ();
 sg13g2_decap_8 FILLER_71_84 ();
 sg13g2_decap_8 FILLER_71_91 ();
 sg13g2_decap_8 FILLER_71_98 ();
 sg13g2_fill_2 FILLER_71_105 ();
 sg13g2_decap_8 FILLER_71_124 ();
 sg13g2_fill_2 FILLER_71_131 ();
 sg13g2_fill_1 FILLER_71_133 ();
 sg13g2_fill_1 FILLER_71_144 ();
 sg13g2_fill_1 FILLER_71_157 ();
 sg13g2_fill_2 FILLER_71_230 ();
 sg13g2_decap_8 FILLER_71_241 ();
 sg13g2_decap_4 FILLER_71_252 ();
 sg13g2_decap_4 FILLER_71_303 ();
 sg13g2_fill_2 FILLER_71_316 ();
 sg13g2_fill_1 FILLER_71_318 ();
 sg13g2_decap_8 FILLER_71_327 ();
 sg13g2_fill_2 FILLER_71_342 ();
 sg13g2_decap_8 FILLER_72_0 ();
 sg13g2_decap_8 FILLER_72_7 ();
 sg13g2_decap_8 FILLER_72_14 ();
 sg13g2_decap_8 FILLER_72_21 ();
 sg13g2_decap_8 FILLER_72_28 ();
 sg13g2_decap_8 FILLER_72_35 ();
 sg13g2_decap_8 FILLER_72_42 ();
 sg13g2_decap_8 FILLER_72_49 ();
 sg13g2_decap_8 FILLER_72_56 ();
 sg13g2_decap_8 FILLER_72_63 ();
 sg13g2_decap_8 FILLER_72_70 ();
 sg13g2_decap_8 FILLER_72_77 ();
 sg13g2_decap_4 FILLER_72_84 ();
 sg13g2_fill_2 FILLER_72_88 ();
 sg13g2_fill_2 FILLER_72_178 ();
 sg13g2_fill_2 FILLER_72_184 ();
 sg13g2_fill_1 FILLER_72_189 ();
 sg13g2_decap_8 FILLER_72_196 ();
 sg13g2_fill_2 FILLER_72_203 ();
 sg13g2_fill_1 FILLER_72_259 ();
 sg13g2_decap_8 FILLER_72_273 ();
 sg13g2_fill_2 FILLER_72_280 ();
 sg13g2_fill_1 FILLER_72_282 ();
 sg13g2_decap_4 FILLER_72_296 ();
 sg13g2_decap_8 FILLER_72_309 ();
 sg13g2_fill_1 FILLER_72_337 ();
 sg13g2_fill_2 FILLER_72_406 ();
 sg13g2_fill_1 FILLER_72_408 ();
 sg13g2_decap_8 FILLER_73_0 ();
 sg13g2_decap_8 FILLER_73_7 ();
 sg13g2_decap_8 FILLER_73_14 ();
 sg13g2_decap_8 FILLER_73_21 ();
 sg13g2_decap_8 FILLER_73_28 ();
 sg13g2_decap_8 FILLER_73_35 ();
 sg13g2_decap_8 FILLER_73_42 ();
 sg13g2_decap_8 FILLER_73_49 ();
 sg13g2_decap_8 FILLER_73_56 ();
 sg13g2_decap_8 FILLER_73_63 ();
 sg13g2_decap_8 FILLER_73_70 ();
 sg13g2_decap_8 FILLER_73_77 ();
 sg13g2_decap_4 FILLER_73_84 ();
 sg13g2_fill_1 FILLER_73_88 ();
 sg13g2_decap_4 FILLER_73_143 ();
 sg13g2_fill_2 FILLER_73_188 ();
 sg13g2_decap_8 FILLER_73_198 ();
 sg13g2_fill_1 FILLER_73_205 ();
 sg13g2_fill_1 FILLER_73_277 ();
 sg13g2_fill_2 FILLER_73_291 ();
 sg13g2_fill_1 FILLER_73_293 ();
 sg13g2_decap_8 FILLER_73_394 ();
 sg13g2_decap_8 FILLER_73_401 ();
 sg13g2_fill_1 FILLER_73_408 ();
 sg13g2_decap_8 FILLER_74_0 ();
 sg13g2_decap_8 FILLER_74_7 ();
 sg13g2_decap_8 FILLER_74_14 ();
 sg13g2_decap_8 FILLER_74_21 ();
 sg13g2_decap_8 FILLER_74_28 ();
 sg13g2_decap_8 FILLER_74_35 ();
 sg13g2_decap_8 FILLER_74_42 ();
 sg13g2_decap_8 FILLER_74_49 ();
 sg13g2_decap_8 FILLER_74_56 ();
 sg13g2_decap_8 FILLER_74_63 ();
 sg13g2_decap_8 FILLER_74_70 ();
 sg13g2_decap_8 FILLER_74_77 ();
 sg13g2_decap_8 FILLER_74_84 ();
 sg13g2_decap_8 FILLER_74_91 ();
 sg13g2_decap_4 FILLER_74_98 ();
 sg13g2_fill_1 FILLER_74_111 ();
 sg13g2_fill_1 FILLER_74_133 ();
 sg13g2_decap_4 FILLER_74_143 ();
 sg13g2_fill_1 FILLER_74_147 ();
 sg13g2_fill_2 FILLER_74_152 ();
 sg13g2_fill_2 FILLER_74_180 ();
 sg13g2_fill_1 FILLER_74_182 ();
 sg13g2_decap_8 FILLER_74_219 ();
 sg13g2_fill_2 FILLER_74_226 ();
 sg13g2_fill_1 FILLER_74_228 ();
 sg13g2_decap_8 FILLER_74_278 ();
 sg13g2_fill_2 FILLER_74_285 ();
 sg13g2_decap_8 FILLER_74_359 ();
 sg13g2_decap_8 FILLER_74_366 ();
 sg13g2_decap_8 FILLER_74_373 ();
 sg13g2_fill_1 FILLER_74_380 ();
 sg13g2_fill_1 FILLER_74_408 ();
 sg13g2_decap_8 FILLER_75_0 ();
 sg13g2_decap_8 FILLER_75_7 ();
 sg13g2_decap_8 FILLER_75_14 ();
 sg13g2_decap_8 FILLER_75_21 ();
 sg13g2_decap_8 FILLER_75_28 ();
 sg13g2_decap_8 FILLER_75_35 ();
 sg13g2_decap_8 FILLER_75_42 ();
 sg13g2_decap_8 FILLER_75_49 ();
 sg13g2_decap_8 FILLER_75_56 ();
 sg13g2_decap_8 FILLER_75_63 ();
 sg13g2_decap_8 FILLER_75_70 ();
 sg13g2_decap_8 FILLER_75_77 ();
 sg13g2_decap_8 FILLER_75_84 ();
 sg13g2_decap_8 FILLER_75_91 ();
 sg13g2_fill_1 FILLER_75_98 ();
 sg13g2_fill_1 FILLER_75_112 ();
 sg13g2_fill_2 FILLER_75_127 ();
 sg13g2_fill_1 FILLER_75_142 ();
 sg13g2_decap_4 FILLER_75_169 ();
 sg13g2_fill_2 FILLER_75_173 ();
 sg13g2_decap_8 FILLER_75_215 ();
 sg13g2_decap_8 FILLER_75_222 ();
 sg13g2_decap_8 FILLER_75_265 ();
 sg13g2_fill_1 FILLER_75_285 ();
 sg13g2_decap_8 FILLER_75_295 ();
 sg13g2_decap_8 FILLER_75_302 ();
 sg13g2_fill_1 FILLER_75_309 ();
 sg13g2_fill_1 FILLER_75_379 ();
 sg13g2_fill_2 FILLER_75_407 ();
 sg13g2_decap_8 FILLER_76_0 ();
 sg13g2_decap_8 FILLER_76_7 ();
 sg13g2_decap_8 FILLER_76_14 ();
 sg13g2_decap_8 FILLER_76_21 ();
 sg13g2_decap_8 FILLER_76_28 ();
 sg13g2_decap_8 FILLER_76_35 ();
 sg13g2_decap_8 FILLER_76_42 ();
 sg13g2_decap_8 FILLER_76_49 ();
 sg13g2_decap_8 FILLER_76_56 ();
 sg13g2_decap_8 FILLER_76_63 ();
 sg13g2_decap_8 FILLER_76_70 ();
 sg13g2_decap_8 FILLER_76_77 ();
 sg13g2_decap_8 FILLER_76_84 ();
 sg13g2_decap_8 FILLER_76_91 ();
 sg13g2_fill_1 FILLER_76_98 ();
 sg13g2_decap_4 FILLER_76_169 ();
 sg13g2_fill_1 FILLER_76_173 ();
 sg13g2_decap_8 FILLER_76_208 ();
 sg13g2_decap_8 FILLER_76_215 ();
 sg13g2_fill_2 FILLER_76_222 ();
 sg13g2_decap_4 FILLER_76_250 ();
 sg13g2_decap_4 FILLER_76_307 ();
 sg13g2_fill_2 FILLER_76_311 ();
 sg13g2_fill_2 FILLER_76_350 ();
 sg13g2_decap_8 FILLER_76_356 ();
 sg13g2_decap_8 FILLER_76_363 ();
 sg13g2_fill_1 FILLER_76_383 ();
 sg13g2_fill_2 FILLER_76_406 ();
 sg13g2_fill_1 FILLER_76_408 ();
 sg13g2_decap_8 FILLER_77_0 ();
 sg13g2_decap_8 FILLER_77_7 ();
 sg13g2_decap_8 FILLER_77_14 ();
 sg13g2_decap_8 FILLER_77_21 ();
 sg13g2_decap_8 FILLER_77_28 ();
 sg13g2_decap_8 FILLER_77_35 ();
 sg13g2_decap_8 FILLER_77_42 ();
 sg13g2_decap_8 FILLER_77_49 ();
 sg13g2_decap_8 FILLER_77_56 ();
 sg13g2_decap_8 FILLER_77_63 ();
 sg13g2_decap_8 FILLER_77_70 ();
 sg13g2_decap_8 FILLER_77_77 ();
 sg13g2_decap_8 FILLER_77_84 ();
 sg13g2_decap_4 FILLER_77_91 ();
 sg13g2_decap_4 FILLER_77_114 ();
 sg13g2_decap_8 FILLER_77_236 ();
 sg13g2_fill_1 FILLER_77_270 ();
 sg13g2_decap_4 FILLER_77_284 ();
 sg13g2_fill_2 FILLER_77_288 ();
 sg13g2_fill_2 FILLER_77_307 ();
 sg13g2_fill_1 FILLER_77_309 ();
 sg13g2_fill_2 FILLER_77_340 ();
 sg13g2_fill_1 FILLER_77_397 ();
 sg13g2_decap_8 FILLER_77_402 ();
 sg13g2_decap_8 FILLER_78_0 ();
 sg13g2_decap_8 FILLER_78_7 ();
 sg13g2_decap_8 FILLER_78_14 ();
 sg13g2_decap_8 FILLER_78_21 ();
 sg13g2_decap_8 FILLER_78_28 ();
 sg13g2_decap_8 FILLER_78_35 ();
 sg13g2_decap_8 FILLER_78_42 ();
 sg13g2_decap_8 FILLER_78_49 ();
 sg13g2_decap_8 FILLER_78_56 ();
 sg13g2_decap_8 FILLER_78_63 ();
 sg13g2_decap_8 FILLER_78_70 ();
 sg13g2_decap_8 FILLER_78_77 ();
 sg13g2_decap_8 FILLER_78_84 ();
 sg13g2_decap_8 FILLER_78_91 ();
 sg13g2_fill_2 FILLER_78_98 ();
 sg13g2_fill_2 FILLER_78_104 ();
 sg13g2_decap_8 FILLER_78_170 ();
 sg13g2_fill_2 FILLER_78_177 ();
 sg13g2_fill_1 FILLER_78_179 ();
 sg13g2_decap_4 FILLER_78_189 ();
 sg13g2_fill_2 FILLER_78_193 ();
 sg13g2_fill_2 FILLER_78_345 ();
 sg13g2_fill_1 FILLER_78_369 ();
 sg13g2_decap_8 FILLER_78_397 ();
 sg13g2_decap_4 FILLER_78_404 ();
 sg13g2_fill_1 FILLER_78_408 ();
 sg13g2_decap_8 FILLER_79_0 ();
 sg13g2_decap_8 FILLER_79_7 ();
 sg13g2_decap_8 FILLER_79_14 ();
 sg13g2_decap_8 FILLER_79_21 ();
 sg13g2_decap_8 FILLER_79_28 ();
 sg13g2_decap_8 FILLER_79_35 ();
 sg13g2_decap_8 FILLER_79_42 ();
 sg13g2_decap_8 FILLER_79_49 ();
 sg13g2_decap_8 FILLER_79_56 ();
 sg13g2_decap_8 FILLER_79_63 ();
 sg13g2_decap_8 FILLER_79_70 ();
 sg13g2_decap_8 FILLER_79_77 ();
 sg13g2_decap_8 FILLER_79_84 ();
 sg13g2_decap_8 FILLER_79_91 ();
 sg13g2_decap_8 FILLER_79_98 ();
 sg13g2_fill_2 FILLER_79_132 ();
 sg13g2_decap_4 FILLER_79_160 ();
 sg13g2_fill_1 FILLER_79_164 ();
 sg13g2_fill_2 FILLER_79_192 ();
 sg13g2_fill_1 FILLER_79_194 ();
 sg13g2_fill_2 FILLER_79_204 ();
 sg13g2_fill_2 FILLER_79_264 ();
 sg13g2_fill_2 FILLER_79_293 ();
 sg13g2_fill_1 FILLER_79_295 ();
 sg13g2_fill_1 FILLER_79_323 ();
 sg13g2_fill_1 FILLER_79_356 ();
 sg13g2_decap_8 FILLER_79_397 ();
 sg13g2_decap_4 FILLER_79_404 ();
 sg13g2_fill_1 FILLER_79_408 ();
 sg13g2_decap_8 FILLER_80_0 ();
 sg13g2_decap_8 FILLER_80_7 ();
 sg13g2_decap_8 FILLER_80_14 ();
 sg13g2_decap_8 FILLER_80_21 ();
 sg13g2_decap_8 FILLER_80_28 ();
 sg13g2_decap_8 FILLER_80_35 ();
 sg13g2_decap_8 FILLER_80_42 ();
 sg13g2_decap_8 FILLER_80_49 ();
 sg13g2_decap_4 FILLER_80_60 ();
 sg13g2_decap_4 FILLER_80_68 ();
 sg13g2_decap_4 FILLER_80_76 ();
 sg13g2_decap_4 FILLER_80_84 ();
 sg13g2_decap_4 FILLER_80_92 ();
 sg13g2_fill_2 FILLER_80_100 ();
 sg13g2_decap_4 FILLER_80_140 ();
 sg13g2_decap_4 FILLER_80_148 ();
 sg13g2_decap_4 FILLER_80_156 ();
 sg13g2_decap_8 FILLER_80_164 ();
 sg13g2_decap_8 FILLER_80_171 ();
 sg13g2_fill_2 FILLER_80_178 ();
 sg13g2_fill_1 FILLER_80_180 ();
 sg13g2_decap_8 FILLER_80_190 ();
 sg13g2_decap_8 FILLER_80_197 ();
 sg13g2_decap_8 FILLER_80_204 ();
 sg13g2_fill_1 FILLER_80_211 ();
 sg13g2_decap_8 FILLER_80_234 ();
 sg13g2_decap_4 FILLER_80_241 ();
 sg13g2_fill_2 FILLER_80_245 ();
 sg13g2_fill_2 FILLER_80_285 ();
 sg13g2_fill_1 FILLER_80_287 ();
 sg13g2_fill_1 FILLER_80_339 ();
 sg13g2_fill_2 FILLER_80_367 ();
 assign uio_oe[0] = net38;
 assign uio_oe[1] = net39;
 assign uio_oe[2] = net20;
 assign uio_oe[3] = net21;
 assign uio_oe[4] = net22;
 assign uio_oe[5] = net23;
 assign uio_oe[6] = net24;
 assign uio_oe[7] = net25;
 assign uio_out[2] = net26;
 assign uio_out[3] = net27;
 assign uio_out[4] = net28;
 assign uio_out[5] = net29;
 assign uio_out[6] = net30;
 assign uio_out[7] = net31;
endmodule
