module tt_um_dranoel06_SAP1 (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire clknet_0_clk;
 wire \cpu0.a_reg[0] ;
 wire \cpu0.a_reg[1] ;
 wire \cpu0.a_reg[2] ;
 wire \cpu0.a_reg[3] ;
 wire \cpu0.a_reg[4] ;
 wire \cpu0.a_reg[5] ;
 wire \cpu0.a_reg[6] ;
 wire \cpu0.a_reg[7] ;
 wire \cpu0.b_reg[0] ;
 wire \cpu0.b_reg[1] ;
 wire \cpu0.b_reg[2] ;
 wire \cpu0.b_reg[3] ;
 wire \cpu0.b_reg[4] ;
 wire \cpu0.b_reg[5] ;
 wire \cpu0.b_reg[6] ;
 wire \cpu0.b_reg[7] ;
 wire \cpu0.ir[0] ;
 wire \cpu0.ir[1] ;
 wire \cpu0.ir[2] ;
 wire \cpu0.ir[3] ;
 wire \cpu0.ir[4] ;
 wire \cpu0.ir[5] ;
 wire \cpu0.ir[6] ;
 wire \cpu0.ir[7] ;
 wire \cpu0.mar[0] ;
 wire \cpu0.mar[1] ;
 wire \cpu0.mar[2] ;
 wire \cpu0.mar[3] ;
 wire \cpu0.pc[0] ;
 wire \cpu0.pc[1] ;
 wire \cpu0.pc[2] ;
 wire \cpu0.pc[3] ;
 wire \cpu0.ram[0][0] ;
 wire \cpu0.ram[0][1] ;
 wire \cpu0.ram[0][2] ;
 wire \cpu0.ram[0][3] ;
 wire \cpu0.ram[0][4] ;
 wire \cpu0.ram[0][5] ;
 wire \cpu0.ram[0][6] ;
 wire \cpu0.ram[0][7] ;
 wire \cpu0.ram[10][0] ;
 wire \cpu0.ram[10][1] ;
 wire \cpu0.ram[10][2] ;
 wire \cpu0.ram[10][3] ;
 wire \cpu0.ram[10][4] ;
 wire \cpu0.ram[10][5] ;
 wire \cpu0.ram[10][6] ;
 wire \cpu0.ram[10][7] ;
 wire \cpu0.ram[11][0] ;
 wire \cpu0.ram[11][1] ;
 wire \cpu0.ram[11][2] ;
 wire \cpu0.ram[11][3] ;
 wire \cpu0.ram[11][4] ;
 wire \cpu0.ram[11][5] ;
 wire \cpu0.ram[11][6] ;
 wire \cpu0.ram[11][7] ;
 wire \cpu0.ram[12][0] ;
 wire \cpu0.ram[12][1] ;
 wire \cpu0.ram[12][2] ;
 wire \cpu0.ram[12][3] ;
 wire \cpu0.ram[12][4] ;
 wire \cpu0.ram[12][5] ;
 wire \cpu0.ram[12][6] ;
 wire \cpu0.ram[12][7] ;
 wire \cpu0.ram[13][0] ;
 wire \cpu0.ram[13][1] ;
 wire \cpu0.ram[13][2] ;
 wire \cpu0.ram[13][3] ;
 wire \cpu0.ram[13][4] ;
 wire \cpu0.ram[13][5] ;
 wire \cpu0.ram[13][6] ;
 wire \cpu0.ram[13][7] ;
 wire \cpu0.ram[14][0] ;
 wire \cpu0.ram[14][1] ;
 wire \cpu0.ram[14][2] ;
 wire \cpu0.ram[14][3] ;
 wire \cpu0.ram[14][4] ;
 wire \cpu0.ram[14][5] ;
 wire \cpu0.ram[14][6] ;
 wire \cpu0.ram[14][7] ;
 wire \cpu0.ram[15][0] ;
 wire \cpu0.ram[15][1] ;
 wire \cpu0.ram[15][2] ;
 wire \cpu0.ram[15][3] ;
 wire \cpu0.ram[15][4] ;
 wire \cpu0.ram[15][5] ;
 wire \cpu0.ram[15][6] ;
 wire \cpu0.ram[15][7] ;
 wire \cpu0.ram[1][0] ;
 wire \cpu0.ram[1][1] ;
 wire \cpu0.ram[1][2] ;
 wire \cpu0.ram[1][3] ;
 wire \cpu0.ram[1][4] ;
 wire \cpu0.ram[1][5] ;
 wire \cpu0.ram[1][6] ;
 wire \cpu0.ram[1][7] ;
 wire \cpu0.ram[2][0] ;
 wire \cpu0.ram[2][1] ;
 wire \cpu0.ram[2][2] ;
 wire \cpu0.ram[2][3] ;
 wire \cpu0.ram[2][4] ;
 wire \cpu0.ram[2][5] ;
 wire \cpu0.ram[2][6] ;
 wire \cpu0.ram[2][7] ;
 wire \cpu0.ram[3][0] ;
 wire \cpu0.ram[3][1] ;
 wire \cpu0.ram[3][2] ;
 wire \cpu0.ram[3][3] ;
 wire \cpu0.ram[3][4] ;
 wire \cpu0.ram[3][5] ;
 wire \cpu0.ram[3][6] ;
 wire \cpu0.ram[3][7] ;
 wire \cpu0.ram[4][0] ;
 wire \cpu0.ram[4][1] ;
 wire \cpu0.ram[4][2] ;
 wire \cpu0.ram[4][3] ;
 wire \cpu0.ram[4][4] ;
 wire \cpu0.ram[4][5] ;
 wire \cpu0.ram[4][6] ;
 wire \cpu0.ram[4][7] ;
 wire \cpu0.ram[5][0] ;
 wire \cpu0.ram[5][1] ;
 wire \cpu0.ram[5][2] ;
 wire \cpu0.ram[5][3] ;
 wire \cpu0.ram[5][4] ;
 wire \cpu0.ram[5][5] ;
 wire \cpu0.ram[5][6] ;
 wire \cpu0.ram[5][7] ;
 wire \cpu0.ram[6][0] ;
 wire \cpu0.ram[6][1] ;
 wire \cpu0.ram[6][2] ;
 wire \cpu0.ram[6][3] ;
 wire \cpu0.ram[6][4] ;
 wire \cpu0.ram[6][5] ;
 wire \cpu0.ram[6][6] ;
 wire \cpu0.ram[6][7] ;
 wire \cpu0.ram[7][0] ;
 wire \cpu0.ram[7][1] ;
 wire \cpu0.ram[7][2] ;
 wire \cpu0.ram[7][3] ;
 wire \cpu0.ram[7][4] ;
 wire \cpu0.ram[7][5] ;
 wire \cpu0.ram[7][6] ;
 wire \cpu0.ram[7][7] ;
 wire \cpu0.ram[8][0] ;
 wire \cpu0.ram[8][1] ;
 wire \cpu0.ram[8][2] ;
 wire \cpu0.ram[8][3] ;
 wire \cpu0.ram[8][4] ;
 wire \cpu0.ram[8][5] ;
 wire \cpu0.ram[8][6] ;
 wire \cpu0.ram[8][7] ;
 wire \cpu0.ram[9][0] ;
 wire \cpu0.ram[9][1] ;
 wire \cpu0.ram[9][2] ;
 wire \cpu0.ram[9][3] ;
 wire \cpu0.ram[9][4] ;
 wire \cpu0.ram[9][5] ;
 wire \cpu0.ram[9][6] ;
 wire \cpu0.ram[9][7] ;
 wire \cpu0.step[0] ;
 wire \cpu0.step[1] ;
 wire \cpu0.step[2] ;
 wire \cpu0.zero_flag ;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire clknet_5_0__leaf_clk;
 wire clknet_5_1__leaf_clk;
 wire clknet_5_2__leaf_clk;
 wire clknet_5_3__leaf_clk;
 wire clknet_5_4__leaf_clk;
 wire clknet_5_5__leaf_clk;
 wire clknet_5_6__leaf_clk;
 wire clknet_5_7__leaf_clk;
 wire clknet_5_8__leaf_clk;
 wire clknet_5_9__leaf_clk;
 wire clknet_5_10__leaf_clk;
 wire clknet_5_11__leaf_clk;
 wire clknet_5_12__leaf_clk;
 wire clknet_5_13__leaf_clk;
 wire clknet_5_14__leaf_clk;
 wire clknet_5_15__leaf_clk;
 wire clknet_5_16__leaf_clk;
 wire clknet_5_17__leaf_clk;
 wire clknet_5_18__leaf_clk;
 wire clknet_5_19__leaf_clk;
 wire clknet_5_20__leaf_clk;
 wire clknet_5_21__leaf_clk;
 wire clknet_5_22__leaf_clk;
 wire clknet_5_23__leaf_clk;
 wire clknet_5_24__leaf_clk;
 wire clknet_5_25__leaf_clk;
 wire clknet_5_26__leaf_clk;
 wire clknet_5_27__leaf_clk;
 wire clknet_5_28__leaf_clk;
 wire clknet_5_29__leaf_clk;
 wire clknet_5_30__leaf_clk;
 wire clknet_5_31__leaf_clk;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;

 sg13g2_inv_1 _0764_ (.Y(_0180_),
    .A(net463));
 sg13g2_inv_1 _0765_ (.Y(_0181_),
    .A(\cpu0.ir[1] ));
 sg13g2_inv_1 _0766_ (.Y(_0182_),
    .A(\cpu0.b_reg[4] ));
 sg13g2_inv_2 _0767_ (.Y(_0183_),
    .A(net193));
 sg13g2_inv_2 _0768_ (.Y(_0184_),
    .A(net175));
 sg13g2_inv_1 _0769_ (.Y(_0185_),
    .A(\cpu0.ram[4][0] ));
 sg13g2_inv_2 _0770_ (.Y(_0186_),
    .A(net169));
 sg13g2_inv_1 _0771_ (.Y(_0187_),
    .A(net281));
 sg13g2_inv_1 _0772_ (.Y(_0188_),
    .A(net167));
 sg13g2_inv_1 _0773_ (.Y(_0189_),
    .A(\cpu0.ram[4][2] ));
 sg13g2_inv_1 _0774_ (.Y(_0190_),
    .A(\cpu0.ram[12][2] ));
 sg13g2_inv_1 _0775_ (.Y(_0191_),
    .A(net285));
 sg13g2_inv_1 _0776_ (.Y(_0192_),
    .A(net275));
 sg13g2_inv_1 _0777_ (.Y(_0193_),
    .A(net280));
 sg13g2_inv_1 _0778_ (.Y(_0194_),
    .A(\cpu0.ram[15][5] ));
 sg13g2_inv_1 _0779_ (.Y(_0195_),
    .A(\cpu0.ram[9][6] ));
 sg13g2_inv_1 _0780_ (.Y(_0196_),
    .A(net282));
 sg13g2_inv_1 _0781_ (.Y(_0197_),
    .A(net277));
 sg13g2_inv_1 _0782_ (.Y(_0198_),
    .A(\cpu0.ram[15][7] ));
 sg13g2_nor2b_2 _0783_ (.A(\cpu0.ir[7] ),
    .B_N(\cpu0.ir[6] ),
    .Y(_0199_));
 sg13g2_nor2_1 _0784_ (.A(net166),
    .B(net464),
    .Y(_0200_));
 sg13g2_nand2_1 _0785_ (.Y(_0201_),
    .A(net459),
    .B(net192));
 sg13g2_nand2b_2 _0786_ (.Y(_0202_),
    .B(\cpu0.ir[4] ),
    .A_N(\cpu0.ir[5] ));
 sg13g2_nor4_2 _0787_ (.A(net166),
    .B(\cpu0.step[0] ),
    .C(_0201_),
    .Y(_0203_),
    .D(_0202_));
 sg13g2_nand2_1 _0788_ (.Y(_0204_),
    .A(_0199_),
    .B(_0203_));
 sg13g2_a21oi_2 _0789_ (.B1(net13),
    .Y(_0205_),
    .A2(_0203_),
    .A1(_0199_));
 sg13g2_nor2_1 _0790_ (.A(net13),
    .B(_0204_),
    .Y(_0206_));
 sg13g2_mux2_1 _0791_ (.A0(net9),
    .A1(\cpu0.mar[0] ),
    .S(net157),
    .X(_0207_));
 sg13g2_nor2b_2 _0792_ (.A(_0205_),
    .B_N(_0207_),
    .Y(_0208_));
 sg13g2_nor2b_1 _0793_ (.A(net158),
    .B_N(net10),
    .Y(_0209_));
 sg13g2_a21oi_2 _0794_ (.B1(_0209_),
    .Y(_0210_),
    .A2(net157),
    .A1(\cpu0.mar[1] ));
 sg13g2_a21o_2 _0795_ (.A2(net157),
    .A1(\cpu0.mar[1] ),
    .B1(_0209_),
    .X(_0211_));
 sg13g2_nand2_1 _0796_ (.Y(_0212_),
    .A(_0208_),
    .B(_0210_));
 sg13g2_mux2_1 _0797_ (.A0(net11),
    .A1(\cpu0.mar[2] ),
    .S(net158),
    .X(_0213_));
 sg13g2_mux2_1 _0798_ (.A0(net12),
    .A1(\cpu0.mar[3] ),
    .S(net158),
    .X(_0214_));
 sg13g2_nand2b_1 _0799_ (.Y(_0215_),
    .B(_0213_),
    .A_N(_0214_));
 sg13g2_or2_1 _0800_ (.X(_0216_),
    .B(_0215_),
    .A(_0212_));
 sg13g2_nor2b_1 _0801_ (.A(net459),
    .B_N(net464),
    .Y(_0217_));
 sg13g2_nor2_2 _0802_ (.A(net459),
    .B(net191),
    .Y(_0218_));
 sg13g2_nand2_1 _0803_ (.Y(_0219_),
    .A(net192),
    .B(_0217_));
 sg13g2_nor2b_1 _0804_ (.A(net166),
    .B_N(net464),
    .Y(_0220_));
 sg13g2_nor2_2 _0805_ (.A(net166),
    .B(_0219_),
    .Y(_0221_));
 sg13g2_or2_1 _0806_ (.X(_0222_),
    .B(_0219_),
    .A(net166));
 sg13g2_mux4_1 _0807_ (.S0(net178),
    .A0(\cpu0.ram[0][0] ),
    .A1(\cpu0.ram[1][0] ),
    .A2(\cpu0.ram[2][0] ),
    .A3(\cpu0.ram[3][0] ),
    .S1(net171),
    .X(_0223_));
 sg13g2_a21oi_1 _0808_ (.A1(net182),
    .A2(\cpu0.ram[5][0] ),
    .Y(_0224_),
    .B1(net174));
 sg13g2_o21ai_1 _0809_ (.B1(_0224_),
    .Y(_0225_),
    .A1(net182),
    .A2(_0185_));
 sg13g2_nor2b_1 _0810_ (.A(net183),
    .B_N(\cpu0.ram[6][0] ),
    .Y(_0226_));
 sg13g2_a21oi_1 _0811_ (.A1(net183),
    .A2(\cpu0.ram[7][0] ),
    .Y(_0227_),
    .B1(_0226_));
 sg13g2_a21oi_1 _0812_ (.A1(net173),
    .A2(_0227_),
    .Y(_0228_),
    .B1(_0186_));
 sg13g2_a221oi_1 _0813_ (.B2(_0228_),
    .C1(net168),
    .B1(_0225_),
    .A1(net163),
    .Y(_0229_),
    .A2(_0223_));
 sg13g2_nor2b_1 _0814_ (.A(net180),
    .B_N(\cpu0.ram[8][0] ),
    .Y(_0230_));
 sg13g2_a21oi_1 _0815_ (.A1(net180),
    .A2(\cpu0.ram[9][0] ),
    .Y(_0231_),
    .B1(_0230_));
 sg13g2_nand2b_1 _0816_ (.Y(_0232_),
    .B(\cpu0.ram[10][0] ),
    .A_N(net180));
 sg13g2_a21oi_1 _0817_ (.A1(net179),
    .A2(\cpu0.ram[11][0] ),
    .Y(_0233_),
    .B1(net165));
 sg13g2_a221oi_1 _0818_ (.B2(_0233_),
    .C1(net169),
    .B1(_0232_),
    .A1(net165),
    .Y(_0234_),
    .A2(_0231_));
 sg13g2_mux2_1 _0819_ (.A0(\cpu0.ram[12][0] ),
    .A1(\cpu0.ram[13][0] ),
    .S(net188),
    .X(_0235_));
 sg13g2_o21ai_1 _0820_ (.B1(net175),
    .Y(_0236_),
    .A1(net186),
    .A2(_0187_));
 sg13g2_a21oi_1 _0821_ (.A1(net186),
    .A2(\cpu0.ram[15][0] ),
    .Y(_0237_),
    .B1(_0236_));
 sg13g2_o21ai_1 _0822_ (.B1(net170),
    .Y(_0238_),
    .A1(net175),
    .A2(_0235_));
 sg13g2_o21ai_1 _0823_ (.B1(_0003_),
    .Y(_0239_),
    .A1(_0237_),
    .A2(_0238_));
 sg13g2_nor2_2 _0824_ (.A(\cpu0.ir[7] ),
    .B(net286),
    .Y(_0240_));
 sg13g2_nor2b_1 _0825_ (.A(\cpu0.ir[4] ),
    .B_N(\cpu0.ir[5] ),
    .Y(_0241_));
 sg13g2_and3_2 _0826_ (.X(_0242_),
    .A(\cpu0.ir[5] ),
    .B(\cpu0.ir[4] ),
    .C(_0199_));
 sg13g2_a21oi_1 _0827_ (.A1(_0240_),
    .A2(_0241_),
    .Y(_0243_),
    .B1(_0242_));
 sg13g2_nand2b_1 _0828_ (.Y(_0244_),
    .B(\cpu0.ir[7] ),
    .A_N(\cpu0.ir[6] ));
 sg13g2_o21ai_1 _0829_ (.B1(_0243_),
    .Y(_0245_),
    .A1(_0202_),
    .A2(_0244_));
 sg13g2_inv_1 _0830_ (.Y(_0246_),
    .A(_0245_));
 sg13g2_nand4_1 _0831_ (.B(net192),
    .C(_0200_),
    .A(net467),
    .Y(_0247_),
    .D(_0245_));
 sg13g2_nor2b_2 _0832_ (.A(net466),
    .B_N(net166),
    .Y(_0248_));
 sg13g2_nand2_2 _0833_ (.Y(_0249_),
    .A(_0218_),
    .B(_0248_));
 sg13g2_nand2_1 _0834_ (.Y(_0250_),
    .A(_0203_),
    .B(_0240_));
 sg13g2_and3_2 _0835_ (.X(_0251_),
    .A(_0247_),
    .B(net162),
    .C(_0250_));
 sg13g2_nand3_1 _0836_ (.B(net162),
    .C(_0250_),
    .A(net156),
    .Y(_0252_));
 sg13g2_o21ai_1 _0837_ (.B1(net155),
    .Y(_0253_),
    .A1(_0234_),
    .A2(_0239_));
 sg13g2_and2_1 _0838_ (.A(net456),
    .B(net464),
    .X(_0254_));
 sg13g2_and2_1 _0839_ (.A(_0218_),
    .B(_0254_),
    .X(_0255_));
 sg13g2_nand2_1 _0840_ (.Y(_0256_),
    .A(_0218_),
    .B(_0254_));
 sg13g2_nand4_1 _0841_ (.B(\cpu0.ir[4] ),
    .C(_0240_),
    .A(net413),
    .Y(_0257_),
    .D(_0255_));
 sg13g2_nand2_2 _0842_ (.Y(_0258_),
    .A(_0204_),
    .B(net161));
 sg13g2_nand2_2 _0843_ (.Y(_0259_),
    .A(\cpu0.step[2] ),
    .B(_0248_));
 sg13g2_nor2_1 _0844_ (.A(_0243_),
    .B(_0259_),
    .Y(_0260_));
 sg13g2_nor3_2 _0845_ (.A(net191),
    .B(_0243_),
    .C(_0259_),
    .Y(_0261_));
 sg13g2_inv_1 _0846_ (.Y(_0262_),
    .A(_0261_));
 sg13g2_nor2b_1 _0847_ (.A(\cpu0.a_reg[0] ),
    .B_N(\cpu0.b_reg[0] ),
    .Y(_0263_));
 sg13g2_xor2_1 _0848_ (.B(net347),
    .A(net292),
    .X(_0264_));
 sg13g2_o21ai_1 _0849_ (.B1(_0246_),
    .Y(_0265_),
    .A1(\cpu0.ir[7] ),
    .A2(_0202_));
 sg13g2_inv_1 _0850_ (.Y(_0266_),
    .A(_0265_));
 sg13g2_nand3_1 _0851_ (.B(net166),
    .C(_0217_),
    .A(\cpu0.zero_flag ),
    .Y(_0267_));
 sg13g2_nor2_1 _0852_ (.A(_0244_),
    .B(_0267_),
    .Y(_0268_));
 sg13g2_nor3_1 _0853_ (.A(\cpu0.ir[5] ),
    .B(\cpu0.ir[4] ),
    .C(_0256_),
    .Y(_0269_));
 sg13g2_o21ai_1 _0854_ (.B1(_0269_),
    .Y(_0270_),
    .A1(_0199_),
    .A2(_0268_));
 sg13g2_and3_2 _0855_ (.X(_0271_),
    .A(_0199_),
    .B(_0241_),
    .C(_0255_));
 sg13g2_a21oi_1 _0856_ (.A1(_0255_),
    .A2(_0265_),
    .Y(_0272_),
    .B1(_0271_));
 sg13g2_nand2_2 _0857_ (.Y(_0273_),
    .A(_0270_),
    .B(_0272_));
 sg13g2_a21o_1 _0858_ (.A2(_0273_),
    .A1(\cpu0.ir[0] ),
    .B1(_0221_),
    .X(_0274_));
 sg13g2_a221oi_1 _0859_ (.B2(_0264_),
    .C1(_0274_),
    .B1(_0261_),
    .A1(\cpu0.a_reg[0] ),
    .Y(_0275_),
    .A2(_0258_));
 sg13g2_o21ai_1 _0860_ (.B1(_0275_),
    .Y(_0276_),
    .A1(_0229_),
    .A2(_0253_));
 sg13g2_o21ai_1 _0861_ (.B1(_0276_),
    .Y(_0277_),
    .A1(\cpu0.pc[0] ),
    .A2(_0222_));
 sg13g2_nor2_1 _0862_ (.A(net1),
    .B(net159),
    .Y(_0278_));
 sg13g2_a21oi_2 _0863_ (.B1(_0278_),
    .Y(_0279_),
    .A2(_0277_),
    .A1(net159));
 sg13g2_mux2_1 _0864_ (.A0(net146),
    .A1(net364),
    .S(_0216_),
    .X(_0004_));
 sg13g2_nor2_1 _0865_ (.A(net2),
    .B(net159),
    .Y(_0280_));
 sg13g2_a21oi_1 _0866_ (.A1(\cpu0.a_reg[1] ),
    .A2(_0258_),
    .Y(_0281_),
    .B1(_0273_));
 sg13g2_nand3b_1 _0867_ (.B(\cpu0.step[0] ),
    .C(\cpu0.step[2] ),
    .Y(_0282_),
    .A_N(net166));
 sg13g2_nor3_1 _0868_ (.A(_0202_),
    .B(_0244_),
    .C(_0282_),
    .Y(_0283_));
 sg13g2_nor2_2 _0869_ (.A(_0242_),
    .B(_0283_),
    .Y(_0284_));
 sg13g2_a21o_2 _0870_ (.A2(_0259_),
    .A1(_0242_),
    .B1(net191),
    .X(_0285_));
 sg13g2_nor2_1 _0871_ (.A(_0284_),
    .B(_0285_),
    .Y(_0286_));
 sg13g2_o21ai_1 _0872_ (.B1(\cpu0.b_reg[0] ),
    .Y(_0287_),
    .A1(_0284_),
    .A2(_0285_));
 sg13g2_xor2_1 _0873_ (.B(_0287_),
    .A(\cpu0.b_reg[1] ),
    .X(_0288_));
 sg13g2_nand2_1 _0874_ (.Y(_0289_),
    .A(\cpu0.a_reg[1] ),
    .B(_0288_));
 sg13g2_xnor2_1 _0875_ (.Y(_0290_),
    .A(\cpu0.a_reg[1] ),
    .B(_0288_));
 sg13g2_a21oi_1 _0876_ (.A1(_0263_),
    .A2(_0290_),
    .Y(_0291_),
    .B1(_0262_));
 sg13g2_o21ai_1 _0877_ (.B1(_0291_),
    .Y(_0292_),
    .A1(_0263_),
    .A2(_0290_));
 sg13g2_a22oi_1 _0878_ (.Y(_0293_),
    .B1(_0281_),
    .B2(_0292_),
    .A2(_0273_),
    .A1(_0181_));
 sg13g2_mux4_1 _0879_ (.S0(net179),
    .A0(\cpu0.ram[8][1] ),
    .A1(\cpu0.ram[9][1] ),
    .A2(\cpu0.ram[10][1] ),
    .A3(\cpu0.ram[11][1] ),
    .S1(net172),
    .X(_0294_));
 sg13g2_nor2b_1 _0880_ (.A(net186),
    .B_N(\cpu0.ram[12][1] ),
    .Y(_0295_));
 sg13g2_a21oi_1 _0881_ (.A1(net186),
    .A2(\cpu0.ram[13][1] ),
    .Y(_0296_),
    .B1(_0295_));
 sg13g2_mux2_1 _0882_ (.A0(\cpu0.ram[14][1] ),
    .A1(\cpu0.ram[15][1] ),
    .S(net184),
    .X(_0297_));
 sg13g2_a21oi_1 _0883_ (.A1(net174),
    .A2(_0297_),
    .Y(_0298_),
    .B1(net164));
 sg13g2_o21ai_1 _0884_ (.B1(_0298_),
    .Y(_0299_),
    .A1(net175),
    .A2(_0296_));
 sg13g2_o21ai_1 _0885_ (.B1(_0299_),
    .Y(_0300_),
    .A1(net169),
    .A2(_0294_));
 sg13g2_mux2_1 _0886_ (.A0(\cpu0.ram[4][1] ),
    .A1(\cpu0.ram[5][1] ),
    .S(net178),
    .X(_0301_));
 sg13g2_mux2_1 _0887_ (.A0(\cpu0.ram[6][1] ),
    .A1(\cpu0.ram[7][1] ),
    .S(net182),
    .X(_0302_));
 sg13g2_mux2_1 _0888_ (.A0(\cpu0.ram[2][1] ),
    .A1(\cpu0.ram[3][1] ),
    .S(net178),
    .X(_0303_));
 sg13g2_mux2_1 _0889_ (.A0(\cpu0.ram[0][1] ),
    .A1(\cpu0.ram[1][1] ),
    .S(net178),
    .X(_0304_));
 sg13g2_mux4_1 _0890_ (.S0(net171),
    .A0(_0301_),
    .A1(_0302_),
    .A2(_0304_),
    .A3(_0303_),
    .S1(net163),
    .X(_0305_));
 sg13g2_o21ai_1 _0891_ (.B1(net155),
    .Y(_0306_),
    .A1(net168),
    .A2(_0305_));
 sg13g2_a21oi_1 _0892_ (.A1(net167),
    .A2(_0300_),
    .Y(_0307_),
    .B1(_0306_));
 sg13g2_or3_1 _0893_ (.A(_0221_),
    .B(_0293_),
    .C(_0307_),
    .X(_0308_));
 sg13g2_o21ai_1 _0894_ (.B1(_0308_),
    .Y(_0309_),
    .A1(\cpu0.pc[1] ),
    .A2(_0222_));
 sg13g2_a21oi_1 _0895_ (.A1(net159),
    .A2(_0309_),
    .Y(_0310_),
    .B1(_0280_));
 sg13g2_mux2_1 _0896_ (.A0(net142),
    .A1(net383),
    .S(_0216_),
    .X(_0005_));
 sg13g2_nor2_1 _0897_ (.A(net3),
    .B(net159),
    .Y(_0311_));
 sg13g2_o21ai_1 _0898_ (.B1(_0289_),
    .Y(_0312_),
    .A1(_0263_),
    .A2(_0290_));
 sg13g2_or2_1 _0899_ (.X(_0313_),
    .B(\cpu0.b_reg[0] ),
    .A(\cpu0.b_reg[1] ));
 sg13g2_o21ai_1 _0900_ (.B1(_0313_),
    .Y(_0314_),
    .A1(_0284_),
    .A2(_0285_));
 sg13g2_xor2_1 _0901_ (.B(_0314_),
    .A(\cpu0.b_reg[2] ),
    .X(_0315_));
 sg13g2_nand2_1 _0902_ (.Y(_0316_),
    .A(\cpu0.a_reg[2] ),
    .B(_0315_));
 sg13g2_xnor2_1 _0903_ (.Y(_0317_),
    .A(\cpu0.a_reg[2] ),
    .B(_0315_));
 sg13g2_nand2b_1 _0904_ (.Y(_0318_),
    .B(_0312_),
    .A_N(_0317_));
 sg13g2_xnor2_1 _0905_ (.Y(_0319_),
    .A(_0312_),
    .B(_0317_));
 sg13g2_a221oi_1 _0906_ (.B2(_0319_),
    .C1(_0273_),
    .B1(_0261_),
    .A1(\cpu0.a_reg[2] ),
    .Y(_0320_),
    .A2(_0258_));
 sg13g2_a21oi_1 _0907_ (.A1(_0270_),
    .A2(_0272_),
    .Y(_0321_),
    .B1(\cpu0.ir[2] ));
 sg13g2_nor3_1 _0908_ (.A(net155),
    .B(_0320_),
    .C(_0321_),
    .Y(_0322_));
 sg13g2_mux4_1 _0909_ (.S0(net179),
    .A0(\cpu0.ram[8][2] ),
    .A1(\cpu0.ram[9][2] ),
    .A2(\cpu0.ram[10][2] ),
    .A3(\cpu0.ram[11][2] ),
    .S1(net172),
    .X(_0323_));
 sg13g2_a21oi_1 _0910_ (.A1(net189),
    .A2(\cpu0.ram[13][2] ),
    .Y(_0324_),
    .B1(net176));
 sg13g2_o21ai_1 _0911_ (.B1(_0324_),
    .Y(_0325_),
    .A1(net189),
    .A2(_0190_));
 sg13g2_nor2b_1 _0912_ (.A(net184),
    .B_N(\cpu0.ram[14][2] ),
    .Y(_0326_));
 sg13g2_a21oi_1 _0913_ (.A1(net184),
    .A2(\cpu0.ram[15][2] ),
    .Y(_0327_),
    .B1(_0326_));
 sg13g2_a21oi_1 _0914_ (.A1(net173),
    .A2(_0327_),
    .Y(_0328_),
    .B1(_0186_));
 sg13g2_a221oi_1 _0915_ (.B2(_0328_),
    .C1(_0188_),
    .B1(_0325_),
    .A1(net164),
    .Y(_0329_),
    .A2(_0323_));
 sg13g2_mux4_1 _0916_ (.S0(net178),
    .A0(\cpu0.ram[0][2] ),
    .A1(\cpu0.ram[1][2] ),
    .A2(\cpu0.ram[2][2] ),
    .A3(\cpu0.ram[3][2] ),
    .S1(net171),
    .X(_0330_));
 sg13g2_a21oi_1 _0917_ (.A1(net182),
    .A2(\cpu0.ram[5][2] ),
    .Y(_0331_),
    .B1(net174));
 sg13g2_o21ai_1 _0918_ (.B1(_0331_),
    .Y(_0332_),
    .A1(net182),
    .A2(_0189_));
 sg13g2_nor2b_1 _0919_ (.A(net183),
    .B_N(\cpu0.ram[6][2] ),
    .Y(_0333_));
 sg13g2_a21oi_1 _0920_ (.A1(net183),
    .A2(\cpu0.ram[7][2] ),
    .Y(_0334_),
    .B1(_0333_));
 sg13g2_a21oi_1 _0921_ (.A1(net173),
    .A2(_0334_),
    .Y(_0335_),
    .B1(net164));
 sg13g2_a221oi_1 _0922_ (.B2(_0335_),
    .C1(net168),
    .B1(_0332_),
    .A1(net163),
    .Y(_0336_),
    .A2(_0330_));
 sg13g2_nor3_1 _0923_ (.A(_0251_),
    .B(_0329_),
    .C(_0336_),
    .Y(_0337_));
 sg13g2_or3_1 _0924_ (.A(_0221_),
    .B(_0322_),
    .C(_0337_),
    .X(_0338_));
 sg13g2_o21ai_1 _0925_ (.B1(_0338_),
    .Y(_0339_),
    .A1(\cpu0.pc[2] ),
    .A2(_0222_));
 sg13g2_a21oi_2 _0926_ (.B1(_0311_),
    .Y(_0340_),
    .A2(_0339_),
    .A1(net159));
 sg13g2_mux2_1 _0927_ (.A0(net140),
    .A1(net352),
    .S(_0216_),
    .X(_0006_));
 sg13g2_or2_1 _0928_ (.X(_0341_),
    .B(_0313_),
    .A(\cpu0.b_reg[2] ));
 sg13g2_o21ai_1 _0929_ (.B1(_0341_),
    .Y(_0342_),
    .A1(_0284_),
    .A2(_0285_));
 sg13g2_xor2_1 _0930_ (.B(_0342_),
    .A(\cpu0.b_reg[3] ),
    .X(_0343_));
 sg13g2_nor2_1 _0931_ (.A(\cpu0.a_reg[3] ),
    .B(_0343_),
    .Y(_0344_));
 sg13g2_xnor2_1 _0932_ (.Y(_0345_),
    .A(\cpu0.a_reg[3] ),
    .B(_0343_));
 sg13g2_a21o_1 _0933_ (.A2(_0318_),
    .A1(_0316_),
    .B1(_0345_),
    .X(_0346_));
 sg13g2_nand3_1 _0934_ (.B(_0318_),
    .C(_0345_),
    .A(_0316_),
    .Y(_0347_));
 sg13g2_nand3_1 _0935_ (.B(_0346_),
    .C(_0347_),
    .A(_0261_),
    .Y(_0348_));
 sg13g2_nand2_1 _0936_ (.Y(_0349_),
    .A(\cpu0.a_reg[3] ),
    .B(_0258_));
 sg13g2_a21oi_1 _0937_ (.A1(\cpu0.ir[3] ),
    .A2(_0273_),
    .Y(_0350_),
    .B1(net155));
 sg13g2_nand3_1 _0938_ (.B(_0349_),
    .C(_0350_),
    .A(_0348_),
    .Y(_0351_));
 sg13g2_mux2_1 _0939_ (.A0(\cpu0.ram[12][3] ),
    .A1(\cpu0.ram[13][3] ),
    .S(net188),
    .X(_0352_));
 sg13g2_nor2b_1 _0940_ (.A(\cpu0.ram[15][3] ),
    .B_N(net186),
    .Y(_0353_));
 sg13g2_o21ai_1 _0941_ (.B1(net175),
    .Y(_0354_),
    .A1(net186),
    .A2(\cpu0.ram[14][3] ));
 sg13g2_o21ai_1 _0942_ (.B1(net170),
    .Y(_0355_),
    .A1(_0353_),
    .A2(_0354_));
 sg13g2_a21o_1 _0943_ (.A2(_0352_),
    .A1(net165),
    .B1(_0355_),
    .X(_0356_));
 sg13g2_mux4_1 _0944_ (.S0(net179),
    .A0(\cpu0.ram[8][3] ),
    .A1(\cpu0.ram[9][3] ),
    .A2(\cpu0.ram[10][3] ),
    .A3(\cpu0.ram[11][3] ),
    .S1(net172),
    .X(_0357_));
 sg13g2_o21ai_1 _0945_ (.B1(net167),
    .Y(_0358_),
    .A1(net169),
    .A2(_0357_));
 sg13g2_nand2b_1 _0946_ (.Y(_0359_),
    .B(_0356_),
    .A_N(_0358_));
 sg13g2_a21oi_1 _0947_ (.A1(net177),
    .A2(_0191_),
    .Y(_0360_),
    .B1(net171));
 sg13g2_o21ai_1 _0948_ (.B1(_0360_),
    .Y(_0361_),
    .A1(net178),
    .A2(\cpu0.ram[0][3] ));
 sg13g2_o21ai_1 _0949_ (.B1(net171),
    .Y(_0362_),
    .A1(net177),
    .A2(\cpu0.ram[2][3] ));
 sg13g2_a21oi_1 _0950_ (.A1(net178),
    .A2(_0192_),
    .Y(_0363_),
    .B1(_0362_));
 sg13g2_nor2_1 _0951_ (.A(net169),
    .B(_0363_),
    .Y(_0364_));
 sg13g2_nand2b_1 _0952_ (.Y(_0365_),
    .B(net184),
    .A_N(\cpu0.ram[5][3] ));
 sg13g2_o21ai_1 _0953_ (.B1(_0365_),
    .Y(_0366_),
    .A1(net185),
    .A2(\cpu0.ram[4][3] ));
 sg13g2_o21ai_1 _0954_ (.B1(net173),
    .Y(_0367_),
    .A1(net184),
    .A2(\cpu0.ram[6][3] ));
 sg13g2_a21oi_1 _0955_ (.A1(net184),
    .A2(_0193_),
    .Y(_0368_),
    .B1(_0367_));
 sg13g2_o21ai_1 _0956_ (.B1(net170),
    .Y(_0369_),
    .A1(net174),
    .A2(_0366_));
 sg13g2_a21oi_1 _0957_ (.A1(_0361_),
    .A2(_0364_),
    .Y(_0370_),
    .B1(net168));
 sg13g2_o21ai_1 _0958_ (.B1(_0370_),
    .Y(_0371_),
    .A1(_0368_),
    .A2(_0369_));
 sg13g2_nand3_1 _0959_ (.B(_0359_),
    .C(_0371_),
    .A(net155),
    .Y(_0372_));
 sg13g2_a22oi_1 _0960_ (.Y(_0373_),
    .B1(_0351_),
    .B2(_0372_),
    .A2(_0221_),
    .A1(\cpu0.pc[3] ));
 sg13g2_nor2_1 _0961_ (.A(net4),
    .B(net159),
    .Y(_0374_));
 sg13g2_a21oi_2 _0962_ (.B1(_0374_),
    .Y(_0375_),
    .A2(_0373_),
    .A1(net160));
 sg13g2_mux2_1 _0963_ (.A0(net139),
    .A1(net362),
    .S(_0216_),
    .X(_0007_));
 sg13g2_nor2_1 _0964_ (.A(_0317_),
    .B(_0345_),
    .Y(_0376_));
 sg13g2_nor2_1 _0965_ (.A(_0316_),
    .B(_0344_),
    .Y(_0377_));
 sg13g2_a221oi_1 _0966_ (.B2(_0312_),
    .C1(_0377_),
    .B1(_0376_),
    .A1(\cpu0.a_reg[3] ),
    .Y(_0378_),
    .A2(_0343_));
 sg13g2_nor2_1 _0967_ (.A(\cpu0.b_reg[3] ),
    .B(_0341_),
    .Y(_0379_));
 sg13g2_nor2_1 _0968_ (.A(_0286_),
    .B(_0379_),
    .Y(_0380_));
 sg13g2_xnor2_1 _0969_ (.Y(_0381_),
    .A(_0182_),
    .B(_0380_));
 sg13g2_nor2b_1 _0970_ (.A(_0381_),
    .B_N(\cpu0.a_reg[4] ),
    .Y(_0382_));
 sg13g2_xnor2_1 _0971_ (.Y(_0383_),
    .A(\cpu0.a_reg[4] ),
    .B(_0381_));
 sg13g2_nor2b_1 _0972_ (.A(_0378_),
    .B_N(_0383_),
    .Y(_0384_));
 sg13g2_xnor2_1 _0973_ (.Y(_0385_),
    .A(_0378_),
    .B(_0383_));
 sg13g2_a22oi_1 _0974_ (.Y(_0386_),
    .B1(_0261_),
    .B2(_0385_),
    .A2(_0258_),
    .A1(\cpu0.a_reg[4] ));
 sg13g2_nand2_1 _0975_ (.Y(_0387_),
    .A(_0251_),
    .B(_0386_));
 sg13g2_mux2_1 _0976_ (.A0(\cpu0.ram[12][4] ),
    .A1(\cpu0.ram[13][4] ),
    .S(net188),
    .X(_0388_));
 sg13g2_nor2b_1 _0977_ (.A(\cpu0.ram[15][4] ),
    .B_N(net187),
    .Y(_0389_));
 sg13g2_o21ai_1 _0978_ (.B1(net175),
    .Y(_0390_),
    .A1(net187),
    .A2(\cpu0.ram[14][4] ));
 sg13g2_o21ai_1 _0979_ (.B1(net170),
    .Y(_0391_),
    .A1(_0389_),
    .A2(_0390_));
 sg13g2_a21oi_1 _0980_ (.A1(_0184_),
    .A2(_0388_),
    .Y(_0392_),
    .B1(_0391_));
 sg13g2_mux4_1 _0981_ (.S0(net179),
    .A0(\cpu0.ram[8][4] ),
    .A1(\cpu0.ram[9][4] ),
    .A2(\cpu0.ram[10][4] ),
    .A3(\cpu0.ram[11][4] ),
    .S1(net172),
    .X(_0393_));
 sg13g2_o21ai_1 _0982_ (.B1(net167),
    .Y(_0394_),
    .A1(net169),
    .A2(_0393_));
 sg13g2_nor2_1 _0983_ (.A(_0392_),
    .B(_0394_),
    .Y(_0395_));
 sg13g2_nand2b_1 _0984_ (.Y(_0396_),
    .B(net181),
    .A_N(\cpu0.ram[5][4] ));
 sg13g2_nand2b_1 _0985_ (.Y(_0397_),
    .B(\cpu0.ram[6][4] ),
    .A_N(net181));
 sg13g2_a21oi_1 _0986_ (.A1(net181),
    .A2(\cpu0.ram[7][4] ),
    .Y(_0398_),
    .B1(net165));
 sg13g2_o21ai_1 _0987_ (.B1(_0396_),
    .Y(_0399_),
    .A1(net181),
    .A2(\cpu0.ram[4][4] ));
 sg13g2_a221oi_1 _0988_ (.B2(net165),
    .C1(net163),
    .B1(_0399_),
    .A1(_0397_),
    .Y(_0400_),
    .A2(_0398_));
 sg13g2_mux4_1 _0989_ (.S0(net177),
    .A0(\cpu0.ram[0][4] ),
    .A1(\cpu0.ram[1][4] ),
    .A2(\cpu0.ram[2][4] ),
    .A3(\cpu0.ram[3][4] ),
    .S1(net171),
    .X(_0401_));
 sg13g2_a21oi_1 _0990_ (.A1(net164),
    .A2(_0401_),
    .Y(_0402_),
    .B1(_0400_));
 sg13g2_o21ai_1 _0991_ (.B1(net155),
    .Y(_0403_),
    .A1(net167),
    .A2(_0402_));
 sg13g2_o21ai_1 _0992_ (.B1(_0387_),
    .Y(_0404_),
    .A1(_0395_),
    .A2(_0403_));
 sg13g2_nor2_1 _0993_ (.A(net5),
    .B(net159),
    .Y(_0405_));
 sg13g2_a21oi_2 _0994_ (.B1(_0405_),
    .Y(_0406_),
    .A2(_0404_),
    .A1(net158));
 sg13g2_mux2_1 _0995_ (.A0(net137),
    .A1(net337),
    .S(_0216_),
    .X(_0008_));
 sg13g2_nor2_1 _0996_ (.A(_0382_),
    .B(_0384_),
    .Y(_0407_));
 sg13g2_a21oi_1 _0997_ (.A1(_0182_),
    .A2(_0379_),
    .Y(_0408_),
    .B1(_0286_));
 sg13g2_o21ai_1 _0998_ (.B1(\cpu0.b_reg[5] ),
    .Y(_0409_),
    .A1(_0284_),
    .A2(_0285_));
 sg13g2_xnor2_1 _0999_ (.Y(_0410_),
    .A(\cpu0.b_reg[5] ),
    .B(_0408_));
 sg13g2_and2_1 _1000_ (.A(\cpu0.a_reg[5] ),
    .B(_0410_),
    .X(_0411_));
 sg13g2_xor2_1 _1001_ (.B(_0410_),
    .A(\cpu0.a_reg[5] ),
    .X(_0412_));
 sg13g2_xnor2_1 _1002_ (.Y(_0413_),
    .A(_0407_),
    .B(_0412_));
 sg13g2_a221oi_1 _1003_ (.B2(_0413_),
    .C1(net155),
    .B1(_0261_),
    .A1(\cpu0.a_reg[5] ),
    .Y(_0414_),
    .A2(_0258_));
 sg13g2_mux2_1 _1004_ (.A0(\cpu0.ram[12][5] ),
    .A1(\cpu0.ram[13][5] ),
    .S(net189),
    .X(_0415_));
 sg13g2_nand2_1 _1005_ (.Y(_0416_),
    .A(_0184_),
    .B(_0415_));
 sg13g2_o21ai_1 _1006_ (.B1(net173),
    .Y(_0417_),
    .A1(net184),
    .A2(\cpu0.ram[14][5] ));
 sg13g2_a21oi_1 _1007_ (.A1(net181),
    .A2(_0194_),
    .Y(_0418_),
    .B1(_0417_));
 sg13g2_nor2_1 _1008_ (.A(net163),
    .B(_0418_),
    .Y(_0419_));
 sg13g2_mux4_1 _1009_ (.S0(net179),
    .A0(\cpu0.ram[8][5] ),
    .A1(\cpu0.ram[9][5] ),
    .A2(\cpu0.ram[10][5] ),
    .A3(\cpu0.ram[11][5] ),
    .S1(net172),
    .X(_0420_));
 sg13g2_o21ai_1 _1010_ (.B1(net167),
    .Y(_0421_),
    .A1(net169),
    .A2(_0420_));
 sg13g2_a21oi_1 _1011_ (.A1(_0416_),
    .A2(_0419_),
    .Y(_0422_),
    .B1(_0421_));
 sg13g2_nand2b_1 _1012_ (.Y(_0423_),
    .B(net183),
    .A_N(\cpu0.ram[7][5] ));
 sg13g2_mux2_1 _1013_ (.A0(\cpu0.ram[4][5] ),
    .A1(\cpu0.ram[5][5] ),
    .S(net182),
    .X(_0424_));
 sg13g2_o21ai_1 _1014_ (.B1(_0423_),
    .Y(_0425_),
    .A1(net183),
    .A2(\cpu0.ram[6][5] ));
 sg13g2_a21oi_1 _1015_ (.A1(net173),
    .A2(_0425_),
    .Y(_0426_),
    .B1(net164));
 sg13g2_o21ai_1 _1016_ (.B1(_0426_),
    .Y(_0427_),
    .A1(net174),
    .A2(_0424_));
 sg13g2_mux4_1 _1017_ (.S0(net177),
    .A0(\cpu0.ram[0][5] ),
    .A1(\cpu0.ram[1][5] ),
    .A2(\cpu0.ram[2][5] ),
    .A3(\cpu0.ram[3][5] ),
    .S1(net171),
    .X(_0428_));
 sg13g2_nand2_1 _1018_ (.Y(_0429_),
    .A(net163),
    .B(_0428_));
 sg13g2_a21oi_1 _1019_ (.A1(_0427_),
    .A2(_0429_),
    .Y(_0430_),
    .B1(net168));
 sg13g2_nor3_1 _1020_ (.A(_0251_),
    .B(_0422_),
    .C(_0430_),
    .Y(_0431_));
 sg13g2_or3_1 _1021_ (.A(_0221_),
    .B(_0414_),
    .C(_0431_),
    .X(_0432_));
 sg13g2_nor2_1 _1022_ (.A(net6),
    .B(net157),
    .Y(_0433_));
 sg13g2_a21oi_2 _1023_ (.B1(_0433_),
    .Y(_0434_),
    .A2(_0432_),
    .A1(net157));
 sg13g2_mux2_1 _1024_ (.A0(net133),
    .A1(net444),
    .S(_0216_),
    .X(_0009_));
 sg13g2_nor2_1 _1025_ (.A(net7),
    .B(net157),
    .Y(_0435_));
 sg13g2_nand2_1 _1026_ (.Y(_0436_),
    .A(_0383_),
    .B(_0412_));
 sg13g2_a21oi_1 _1027_ (.A1(_0382_),
    .A2(_0412_),
    .Y(_0437_),
    .B1(_0411_));
 sg13g2_o21ai_1 _1028_ (.B1(_0437_),
    .Y(_0438_),
    .A1(_0378_),
    .A2(_0436_));
 sg13g2_nand2b_1 _1029_ (.Y(_0439_),
    .B(_0409_),
    .A_N(_0408_));
 sg13g2_nor2_1 _1030_ (.A(\cpu0.b_reg[6] ),
    .B(_0439_),
    .Y(_0440_));
 sg13g2_xor2_1 _1031_ (.B(_0439_),
    .A(\cpu0.b_reg[6] ),
    .X(_0441_));
 sg13g2_nor2b_1 _1032_ (.A(_0441_),
    .B_N(\cpu0.a_reg[6] ),
    .Y(_0442_));
 sg13g2_xnor2_1 _1033_ (.Y(_0443_),
    .A(\cpu0.a_reg[6] ),
    .B(_0441_));
 sg13g2_xor2_1 _1034_ (.B(_0443_),
    .A(_0438_),
    .X(_0444_));
 sg13g2_a221oi_1 _1035_ (.B2(_0444_),
    .C1(_0252_),
    .B1(_0261_),
    .A1(\cpu0.a_reg[6] ),
    .Y(_0445_),
    .A2(_0258_));
 sg13g2_o21ai_1 _1036_ (.B1(net165),
    .Y(_0446_),
    .A1(net180),
    .A2(\cpu0.ram[8][6] ));
 sg13g2_a21oi_1 _1037_ (.A1(net180),
    .A2(_0195_),
    .Y(_0447_),
    .B1(_0446_));
 sg13g2_o21ai_1 _1038_ (.B1(net176),
    .Y(_0448_),
    .A1(net179),
    .A2(\cpu0.ram[10][6] ));
 sg13g2_a21oi_1 _1039_ (.A1(net180),
    .A2(_0196_),
    .Y(_0449_),
    .B1(_0448_));
 sg13g2_nor3_1 _1040_ (.A(net170),
    .B(_0447_),
    .C(_0449_),
    .Y(_0450_));
 sg13g2_nand2b_1 _1041_ (.Y(_0451_),
    .B(net186),
    .A_N(\cpu0.ram[13][6] ));
 sg13g2_o21ai_1 _1042_ (.B1(_0451_),
    .Y(_0452_),
    .A1(net187),
    .A2(\cpu0.ram[12][6] ));
 sg13g2_o21ai_1 _1043_ (.B1(net173),
    .Y(_0453_),
    .A1(net184),
    .A2(\cpu0.ram[14][6] ));
 sg13g2_a21oi_1 _1044_ (.A1(net186),
    .A2(_0197_),
    .Y(_0454_),
    .B1(_0453_));
 sg13g2_o21ai_1 _1045_ (.B1(net170),
    .Y(_0455_),
    .A1(net175),
    .A2(_0452_));
 sg13g2_o21ai_1 _1046_ (.B1(_0003_),
    .Y(_0456_),
    .A1(_0454_),
    .A2(_0455_));
 sg13g2_nor2_1 _1047_ (.A(_0450_),
    .B(_0456_),
    .Y(_0457_));
 sg13g2_nand2b_1 _1048_ (.Y(_0458_),
    .B(net177),
    .A_N(\cpu0.ram[3][6] ));
 sg13g2_nand2b_1 _1049_ (.Y(_0459_),
    .B(net183),
    .A_N(\cpu0.ram[7][6] ));
 sg13g2_mux2_1 _1050_ (.A0(\cpu0.ram[0][6] ),
    .A1(\cpu0.ram[1][6] ),
    .S(net177),
    .X(_0460_));
 sg13g2_o21ai_1 _1051_ (.B1(_0458_),
    .Y(_0461_),
    .A1(net177),
    .A2(\cpu0.ram[2][6] ));
 sg13g2_a21oi_1 _1052_ (.A1(net172),
    .A2(_0461_),
    .Y(_0462_),
    .B1(net169));
 sg13g2_o21ai_1 _1053_ (.B1(_0462_),
    .Y(_0463_),
    .A1(net172),
    .A2(_0460_));
 sg13g2_mux2_1 _1054_ (.A0(\cpu0.ram[4][6] ),
    .A1(\cpu0.ram[5][6] ),
    .S(net182),
    .X(_0464_));
 sg13g2_o21ai_1 _1055_ (.B1(_0459_),
    .Y(_0465_),
    .A1(net183),
    .A2(\cpu0.ram[6][6] ));
 sg13g2_a21oi_1 _1056_ (.A1(net173),
    .A2(_0465_),
    .Y(_0466_),
    .B1(net164));
 sg13g2_o21ai_1 _1057_ (.B1(_0466_),
    .Y(_0467_),
    .A1(net174),
    .A2(_0464_));
 sg13g2_a21oi_1 _1058_ (.A1(_0463_),
    .A2(_0467_),
    .Y(_0468_),
    .B1(net168));
 sg13g2_nor3_1 _1059_ (.A(_0251_),
    .B(_0457_),
    .C(_0468_),
    .Y(_0469_));
 sg13g2_or3_1 _1060_ (.A(_0221_),
    .B(_0445_),
    .C(_0469_),
    .X(_0470_));
 sg13g2_a21oi_2 _1061_ (.B1(_0435_),
    .Y(_0471_),
    .A2(_0470_),
    .A1(net157));
 sg13g2_mux2_1 _1062_ (.A0(net135),
    .A1(net324),
    .S(_0216_),
    .X(_0010_));
 sg13g2_a21oi_1 _1063_ (.A1(_0438_),
    .A2(_0443_),
    .Y(_0472_),
    .B1(_0442_));
 sg13g2_nor2_1 _1064_ (.A(_0286_),
    .B(_0440_),
    .Y(_0473_));
 sg13g2_xnor2_1 _1065_ (.Y(_0474_),
    .A(\cpu0.a_reg[7] ),
    .B(\cpu0.b_reg[7] ));
 sg13g2_xnor2_1 _1066_ (.Y(_0475_),
    .A(_0473_),
    .B(_0474_));
 sg13g2_xnor2_1 _1067_ (.Y(_0476_),
    .A(_0472_),
    .B(_0475_));
 sg13g2_a21oi_1 _1068_ (.A1(net290),
    .A2(_0258_),
    .Y(_0477_),
    .B1(_0252_));
 sg13g2_o21ai_1 _1069_ (.B1(_0477_),
    .Y(_0478_),
    .A1(_0262_),
    .A2(_0476_));
 sg13g2_mux2_1 _1070_ (.A0(\cpu0.ram[12][7] ),
    .A1(\cpu0.ram[13][7] ),
    .S(net189),
    .X(_0479_));
 sg13g2_nand2_1 _1071_ (.Y(_0480_),
    .A(_0184_),
    .B(_0479_));
 sg13g2_o21ai_1 _1072_ (.B1(net174),
    .Y(_0481_),
    .A1(net185),
    .A2(\cpu0.ram[14][7] ));
 sg13g2_a21oi_1 _1073_ (.A1(net189),
    .A2(_0198_),
    .Y(_0482_),
    .B1(_0481_));
 sg13g2_nor2_1 _1074_ (.A(net163),
    .B(_0482_),
    .Y(_0483_));
 sg13g2_mux4_1 _1075_ (.S0(net179),
    .A0(\cpu0.ram[8][7] ),
    .A1(\cpu0.ram[9][7] ),
    .A2(\cpu0.ram[10][7] ),
    .A3(\cpu0.ram[11][7] ),
    .S1(net176),
    .X(_0484_));
 sg13g2_o21ai_1 _1076_ (.B1(net167),
    .Y(_0485_),
    .A1(net170),
    .A2(_0484_));
 sg13g2_a21oi_1 _1077_ (.A1(_0480_),
    .A2(_0483_),
    .Y(_0486_),
    .B1(_0485_));
 sg13g2_nand2b_1 _1078_ (.Y(_0487_),
    .B(net182),
    .A_N(\cpu0.ram[5][7] ));
 sg13g2_nand2b_1 _1079_ (.Y(_0488_),
    .B(\cpu0.ram[6][7] ),
    .A_N(net181));
 sg13g2_a21oi_1 _1080_ (.A1(net181),
    .A2(\cpu0.ram[7][7] ),
    .Y(_0489_),
    .B1(net165));
 sg13g2_o21ai_1 _1081_ (.B1(_0487_),
    .Y(_0490_),
    .A1(net181),
    .A2(\cpu0.ram[4][7] ));
 sg13g2_a221oi_1 _1082_ (.B2(net165),
    .C1(net163),
    .B1(_0490_),
    .A1(_0488_),
    .Y(_0491_),
    .A2(_0489_));
 sg13g2_mux4_1 _1083_ (.S0(net177),
    .A0(\cpu0.ram[0][7] ),
    .A1(\cpu0.ram[1][7] ),
    .A2(\cpu0.ram[2][7] ),
    .A3(\cpu0.ram[3][7] ),
    .S1(net171),
    .X(_0492_));
 sg13g2_a21oi_1 _1084_ (.A1(net164),
    .A2(_0492_),
    .Y(_0493_),
    .B1(_0491_));
 sg13g2_o21ai_1 _1085_ (.B1(net155),
    .Y(_0494_),
    .A1(net167),
    .A2(_0493_));
 sg13g2_o21ai_1 _1086_ (.B1(_0222_),
    .Y(_0495_),
    .A1(_0486_),
    .A2(_0494_));
 sg13g2_nand2b_2 _1087_ (.Y(_0496_),
    .B(_0478_),
    .A_N(_0495_));
 sg13g2_nor2_1 _1088_ (.A(net8),
    .B(net158),
    .Y(_0497_));
 sg13g2_a21oi_2 _1089_ (.B1(_0497_),
    .Y(_0498_),
    .A2(_0496_),
    .A1(net157));
 sg13g2_mux2_1 _1090_ (.A0(net131),
    .A1(net320),
    .S(_0216_),
    .X(_0011_));
 sg13g2_a21oi_1 _1091_ (.A1(net456),
    .A2(_0266_),
    .Y(_0499_),
    .B1(_0219_));
 sg13g2_o21ai_1 _1092_ (.B1(net192),
    .Y(_0500_),
    .A1(net457),
    .A2(net152));
 sg13g2_a21oi_1 _1093_ (.A1(_0277_),
    .A2(net152),
    .Y(_0012_),
    .B1(_0500_));
 sg13g2_o21ai_1 _1094_ (.B1(net192),
    .Y(_0501_),
    .A1(net462),
    .A2(net152));
 sg13g2_a21oi_1 _1095_ (.A1(_0309_),
    .A2(net152),
    .Y(_0013_),
    .B1(_0501_));
 sg13g2_o21ai_1 _1096_ (.B1(net192),
    .Y(_0502_),
    .A1(net454),
    .A2(net152));
 sg13g2_a21oi_1 _1097_ (.A1(_0339_),
    .A2(net152),
    .Y(_0014_),
    .B1(_0502_));
 sg13g2_o21ai_1 _1098_ (.B1(net193),
    .Y(_0503_),
    .A1(net452),
    .A2(net153));
 sg13g2_a21oi_1 _1099_ (.A1(_0373_),
    .A2(net152),
    .Y(_0015_),
    .B1(_0503_));
 sg13g2_nand2_1 _1100_ (.Y(_0504_),
    .A(_0213_),
    .B(_0214_));
 sg13g2_nor2_2 _1101_ (.A(_0205_),
    .B(_0207_),
    .Y(_0505_));
 sg13g2_nand2_1 _1102_ (.Y(_0506_),
    .A(_0211_),
    .B(_0505_));
 sg13g2_or2_1 _1103_ (.X(_0507_),
    .B(_0506_),
    .A(_0504_));
 sg13g2_nor2_1 _1104_ (.A(net146),
    .B(net151),
    .Y(_0508_));
 sg13g2_a21oi_1 _1105_ (.A1(_0187_),
    .A2(net151),
    .Y(_0016_),
    .B1(_0508_));
 sg13g2_mux2_1 _1106_ (.A0(net144),
    .A1(net377),
    .S(_0507_),
    .X(_0017_));
 sg13g2_mux2_1 _1107_ (.A0(net141),
    .A1(net367),
    .S(net151),
    .X(_0018_));
 sg13g2_mux2_1 _1108_ (.A0(net139),
    .A1(net429),
    .S(net151),
    .X(_0019_));
 sg13g2_mux2_1 _1109_ (.A0(net137),
    .A1(net422),
    .S(net151),
    .X(_0020_));
 sg13g2_mux2_1 _1110_ (.A0(net133),
    .A1(net335),
    .S(net151),
    .X(_0021_));
 sg13g2_mux2_1 _1111_ (.A0(net135),
    .A1(net391),
    .S(net151),
    .X(_0022_));
 sg13g2_mux2_1 _1112_ (.A0(net131),
    .A1(net376),
    .S(net151),
    .X(_0023_));
 sg13g2_or2_1 _1113_ (.X(_0509_),
    .B(_0504_),
    .A(_0212_));
 sg13g2_mux2_1 _1114_ (.A0(net146),
    .A1(net412),
    .S(_0509_),
    .X(_0024_));
 sg13g2_mux2_1 _1115_ (.A0(net144),
    .A1(net332),
    .S(_0509_),
    .X(_0025_));
 sg13g2_mux2_1 _1116_ (.A0(net141),
    .A1(net398),
    .S(_0509_),
    .X(_0026_));
 sg13g2_mux2_1 _1117_ (.A0(net139),
    .A1(net351),
    .S(_0509_),
    .X(_0027_));
 sg13g2_mux2_1 _1118_ (.A0(net137),
    .A1(net349),
    .S(_0509_),
    .X(_0028_));
 sg13g2_mux2_1 _1119_ (.A0(net133),
    .A1(net311),
    .S(_0509_),
    .X(_0029_));
 sg13g2_mux2_1 _1120_ (.A0(net135),
    .A1(net379),
    .S(_0509_),
    .X(_0030_));
 sg13g2_mux2_1 _1121_ (.A0(net131),
    .A1(net341),
    .S(_0509_),
    .X(_0031_));
 sg13g2_nor3_1 _1122_ (.A(net191),
    .B(_0200_),
    .C(_0254_),
    .Y(_0032_));
 sg13g2_o21ai_1 _1123_ (.B1(_0256_),
    .Y(_0033_),
    .A1(_0201_),
    .A2(_0254_));
 sg13g2_nand2_1 _1124_ (.Y(_0510_),
    .A(_0210_),
    .B(_0505_));
 sg13g2_or2_1 _1125_ (.X(_0511_),
    .B(_0510_),
    .A(_0504_));
 sg13g2_mux2_1 _1126_ (.A0(net146),
    .A1(net316),
    .S(_0511_),
    .X(_0034_));
 sg13g2_mux2_1 _1127_ (.A0(net144),
    .A1(net302),
    .S(_0511_),
    .X(_0035_));
 sg13g2_mux2_1 _1128_ (.A0(net141),
    .A1(net369),
    .S(_0511_),
    .X(_0036_));
 sg13g2_mux2_1 _1129_ (.A0(net139),
    .A1(net396),
    .S(_0511_),
    .X(_0037_));
 sg13g2_mux2_1 _1130_ (.A0(net137),
    .A1(net425),
    .S(_0511_),
    .X(_0038_));
 sg13g2_mux2_1 _1131_ (.A0(net133),
    .A1(net393),
    .S(_0511_),
    .X(_0039_));
 sg13g2_mux2_1 _1132_ (.A0(net135),
    .A1(net353),
    .S(_0511_),
    .X(_0040_));
 sg13g2_mux2_1 _1133_ (.A0(net131),
    .A1(net445),
    .S(_0511_),
    .X(_0041_));
 sg13g2_nor3_1 _1134_ (.A(net191),
    .B(_0217_),
    .C(_0220_),
    .Y(_0042_));
 sg13g2_or2_1 _1135_ (.X(_0512_),
    .B(_0510_),
    .A(_0215_));
 sg13g2_mux2_1 _1136_ (.A0(net145),
    .A1(net368),
    .S(_0512_),
    .X(_0043_));
 sg13g2_mux2_1 _1137_ (.A0(net142),
    .A1(net374),
    .S(_0512_),
    .X(_0044_));
 sg13g2_mux2_1 _1138_ (.A0(net140),
    .A1(net386),
    .S(_0512_),
    .X(_0045_));
 sg13g2_mux2_1 _1139_ (.A0(net139),
    .A1(net327),
    .S(_0512_),
    .X(_0046_));
 sg13g2_mux2_1 _1140_ (.A0(net137),
    .A1(net356),
    .S(_0512_),
    .X(_0047_));
 sg13g2_mux2_1 _1141_ (.A0(net133),
    .A1(net329),
    .S(_0512_),
    .X(_0048_));
 sg13g2_mux2_1 _1142_ (.A0(net135),
    .A1(net423),
    .S(_0512_),
    .X(_0049_));
 sg13g2_mux2_1 _1143_ (.A0(net131),
    .A1(net380),
    .S(_0512_),
    .X(_0050_));
 sg13g2_nor2_2 _1144_ (.A(_0213_),
    .B(_0214_),
    .Y(_0513_));
 sg13g2_nand2_1 _1145_ (.Y(_0514_),
    .A(_0208_),
    .B(_0211_));
 sg13g2_inv_1 _1146_ (.Y(_0515_),
    .A(_0514_));
 sg13g2_nand2_2 _1147_ (.Y(_0516_),
    .A(_0513_),
    .B(_0515_));
 sg13g2_mux2_1 _1148_ (.A0(net145),
    .A1(net426),
    .S(net148),
    .X(_0051_));
 sg13g2_mux2_1 _1149_ (.A0(net142),
    .A1(net359),
    .S(net148),
    .X(_0052_));
 sg13g2_mux2_1 _1150_ (.A0(net140),
    .A1(net411),
    .S(_0516_),
    .X(_0053_));
 sg13g2_nor2_1 _1151_ (.A(net138),
    .B(net148),
    .Y(_0517_));
 sg13g2_a21oi_1 _1152_ (.A1(_0192_),
    .A2(net148),
    .Y(_0054_),
    .B1(_0517_));
 sg13g2_mux2_1 _1153_ (.A0(net136),
    .A1(net331),
    .S(net148),
    .X(_0055_));
 sg13g2_mux2_1 _1154_ (.A0(net132),
    .A1(net357),
    .S(net148),
    .X(_0056_));
 sg13g2_mux2_1 _1155_ (.A0(net134),
    .A1(net303),
    .S(net148),
    .X(_0057_));
 sg13g2_mux2_1 _1156_ (.A0(net130),
    .A1(net363),
    .S(net148),
    .X(_0058_));
 sg13g2_nand3_1 _1157_ (.B(_0505_),
    .C(_0513_),
    .A(_0211_),
    .Y(_0518_));
 sg13g2_mux2_1 _1158_ (.A0(net145),
    .A1(net312),
    .S(_0518_),
    .X(_0059_));
 sg13g2_mux2_1 _1159_ (.A0(net142),
    .A1(net325),
    .S(_0518_),
    .X(_0060_));
 sg13g2_mux2_1 _1160_ (.A0(net140),
    .A1(net343),
    .S(_0518_),
    .X(_0061_));
 sg13g2_mux2_1 _1161_ (.A0(net138),
    .A1(net344),
    .S(_0518_),
    .X(_0062_));
 sg13g2_mux2_1 _1162_ (.A0(net136),
    .A1(net432),
    .S(_0518_),
    .X(_0063_));
 sg13g2_mux2_1 _1163_ (.A0(net132),
    .A1(net392),
    .S(_0518_),
    .X(_0064_));
 sg13g2_mux2_1 _1164_ (.A0(net134),
    .A1(net371),
    .S(_0518_),
    .X(_0065_));
 sg13g2_mux2_1 _1165_ (.A0(net130),
    .A1(net443),
    .S(_0518_),
    .X(_0066_));
 sg13g2_nand3_1 _1166_ (.B(_0210_),
    .C(_0513_),
    .A(_0208_),
    .Y(_0519_));
 sg13g2_mux2_1 _1167_ (.A0(net145),
    .A1(net410),
    .S(net154),
    .X(_0067_));
 sg13g2_mux2_1 _1168_ (.A0(net142),
    .A1(net384),
    .S(net154),
    .X(_0068_));
 sg13g2_mux2_1 _1169_ (.A0(net140),
    .A1(net355),
    .S(_0519_),
    .X(_0069_));
 sg13g2_nor2_1 _1170_ (.A(net138),
    .B(net154),
    .Y(_0520_));
 sg13g2_a21oi_1 _1171_ (.A1(_0191_),
    .A2(net154),
    .Y(_0070_),
    .B1(_0520_));
 sg13g2_mux2_1 _1172_ (.A0(net136),
    .A1(net431),
    .S(net154),
    .X(_0071_));
 sg13g2_mux2_1 _1173_ (.A0(net132),
    .A1(net441),
    .S(net154),
    .X(_0072_));
 sg13g2_mux2_1 _1174_ (.A0(net134),
    .A1(net378),
    .S(net154),
    .X(_0073_));
 sg13g2_mux2_1 _1175_ (.A0(net130),
    .A1(net401),
    .S(net154),
    .X(_0074_));
 sg13g2_or2_1 _1176_ (.X(_0521_),
    .B(_0514_),
    .A(_0504_));
 sg13g2_mux2_1 _1177_ (.A0(net146),
    .A1(net336),
    .S(net150),
    .X(_0075_));
 sg13g2_mux2_1 _1178_ (.A0(net144),
    .A1(net342),
    .S(net150),
    .X(_0076_));
 sg13g2_mux2_1 _1179_ (.A0(net141),
    .A1(net442),
    .S(_0521_),
    .X(_0077_));
 sg13g2_mux2_1 _1180_ (.A0(net139),
    .A1(net345),
    .S(net150),
    .X(_0078_));
 sg13g2_mux2_1 _1181_ (.A0(net137),
    .A1(net322),
    .S(net150),
    .X(_0079_));
 sg13g2_mux2_1 _1182_ (.A0(net133),
    .A1(net358),
    .S(net150),
    .X(_0080_));
 sg13g2_nor2_1 _1183_ (.A(net135),
    .B(net150),
    .Y(_0522_));
 sg13g2_a21oi_1 _1184_ (.A1(_0197_),
    .A2(net150),
    .Y(_0081_),
    .B1(_0522_));
 sg13g2_mux2_1 _1185_ (.A0(net131),
    .A1(net365),
    .S(net150),
    .X(_0082_));
 sg13g2_nor2_1 _1186_ (.A(_0260_),
    .B(_0283_),
    .Y(_0523_));
 sg13g2_or4_1 _1187_ (.A(_0290_),
    .B(_0317_),
    .C(_0345_),
    .D(_0436_),
    .X(_0524_));
 sg13g2_nor4_1 _1188_ (.A(_0264_),
    .B(_0444_),
    .C(_0523_),
    .D(_0524_),
    .Y(_0525_));
 sg13g2_a22oi_1 _1189_ (.Y(_0526_),
    .B1(_0525_),
    .B2(_0476_),
    .A2(_0523_),
    .A1(net451));
 sg13g2_nor2_1 _1190_ (.A(net191),
    .B(_0526_),
    .Y(_0083_));
 sg13g2_and2_1 _1191_ (.A(net193),
    .B(_0247_),
    .X(_0527_));
 sg13g2_nand2_1 _1192_ (.Y(_0528_),
    .A(net347),
    .B(_0527_));
 sg13g2_o21ai_1 _1193_ (.B1(_0528_),
    .Y(_0084_),
    .A1(_0247_),
    .A2(_0277_));
 sg13g2_nand2_1 _1194_ (.Y(_0529_),
    .A(net295),
    .B(_0527_));
 sg13g2_o21ai_1 _1195_ (.B1(_0529_),
    .Y(_0085_),
    .A1(net156),
    .A2(_0309_));
 sg13g2_nand2_1 _1196_ (.Y(_0530_),
    .A(net283),
    .B(_0527_));
 sg13g2_o21ai_1 _1197_ (.B1(_0530_),
    .Y(_0086_),
    .A1(net156),
    .A2(_0339_));
 sg13g2_nand2_1 _1198_ (.Y(_0531_),
    .A(net297),
    .B(_0527_));
 sg13g2_o21ai_1 _1199_ (.B1(_0531_),
    .Y(_0087_),
    .A1(net156),
    .A2(_0373_));
 sg13g2_nand2_1 _1200_ (.Y(_0532_),
    .A(net272),
    .B(_0527_));
 sg13g2_o21ai_1 _1201_ (.B1(_0532_),
    .Y(_0088_),
    .A1(net156),
    .A2(_0404_));
 sg13g2_nand2_1 _1202_ (.Y(_0533_),
    .A(net372),
    .B(_0527_));
 sg13g2_o21ai_1 _1203_ (.B1(_0533_),
    .Y(_0089_),
    .A1(net156),
    .A2(_0432_));
 sg13g2_nand2_1 _1204_ (.Y(_0534_),
    .A(net304),
    .B(_0527_));
 sg13g2_o21ai_1 _1205_ (.B1(_0534_),
    .Y(_0090_),
    .A1(net156),
    .A2(_0470_));
 sg13g2_nand2_1 _1206_ (.Y(_0535_),
    .A(net278),
    .B(_0527_));
 sg13g2_o21ai_1 _1207_ (.B1(_0535_),
    .Y(_0091_),
    .A1(net156),
    .A2(_0496_));
 sg13g2_a21oi_2 _1208_ (.B1(_0261_),
    .Y(_0536_),
    .A2(_0240_),
    .A1(_0203_));
 sg13g2_nor2b_2 _1209_ (.A(_0271_),
    .B_N(_0536_),
    .Y(_0537_));
 sg13g2_and2_1 _1210_ (.A(net193),
    .B(_0537_),
    .X(_0538_));
 sg13g2_nand2_1 _1211_ (.Y(_0539_),
    .A(net292),
    .B(_0538_));
 sg13g2_o21ai_1 _1212_ (.B1(_0539_),
    .Y(_0092_),
    .A1(_0277_),
    .A2(_0537_));
 sg13g2_nand2_1 _1213_ (.Y(_0540_),
    .A(net301),
    .B(_0538_));
 sg13g2_o21ai_1 _1214_ (.B1(_0540_),
    .Y(_0093_),
    .A1(_0309_),
    .A2(_0537_));
 sg13g2_nand2_1 _1215_ (.Y(_0541_),
    .A(net300),
    .B(_0538_));
 sg13g2_o21ai_1 _1216_ (.B1(_0541_),
    .Y(_0094_),
    .A1(_0339_),
    .A2(_0537_));
 sg13g2_nand2_1 _1217_ (.Y(_0542_),
    .A(net450),
    .B(_0538_));
 sg13g2_o21ai_1 _1218_ (.B1(_0542_),
    .Y(_0095_),
    .A1(_0373_),
    .A2(_0537_));
 sg13g2_nand2_1 _1219_ (.Y(_0543_),
    .A(net298),
    .B(_0538_));
 sg13g2_o21ai_1 _1220_ (.B1(_0543_),
    .Y(_0096_),
    .A1(_0404_),
    .A2(_0536_));
 sg13g2_nand2_1 _1221_ (.Y(_0544_),
    .A(net404),
    .B(_0538_));
 sg13g2_o21ai_1 _1222_ (.B1(_0544_),
    .Y(_0097_),
    .A1(_0432_),
    .A2(_0536_));
 sg13g2_nand2_1 _1223_ (.Y(_0545_),
    .A(net333),
    .B(_0538_));
 sg13g2_o21ai_1 _1224_ (.B1(_0545_),
    .Y(_0098_),
    .A1(_0470_),
    .A2(_0536_));
 sg13g2_nand2_1 _1225_ (.Y(_0546_),
    .A(net290),
    .B(_0538_));
 sg13g2_o21ai_1 _1226_ (.B1(_0546_),
    .Y(_0099_),
    .A1(_0496_),
    .A2(_0536_));
 sg13g2_a21oi_2 _1227_ (.B1(_0183_),
    .Y(_0547_),
    .A2(_0248_),
    .A1(_0218_));
 sg13g2_nand2_1 _1228_ (.Y(_0548_),
    .A(net270),
    .B(_0547_));
 sg13g2_o21ai_1 _1229_ (.B1(_0548_),
    .Y(_0100_),
    .A1(net162),
    .A2(_0277_));
 sg13g2_nand2_1 _1230_ (.Y(_0549_),
    .A(net274),
    .B(_0547_));
 sg13g2_o21ai_1 _1231_ (.B1(_0549_),
    .Y(_0101_),
    .A1(net162),
    .A2(_0309_));
 sg13g2_nand2_1 _1232_ (.Y(_0550_),
    .A(net271),
    .B(_0547_));
 sg13g2_o21ai_1 _1233_ (.B1(_0550_),
    .Y(_0102_),
    .A1(net162),
    .A2(_0339_));
 sg13g2_nand2_1 _1234_ (.Y(_0551_),
    .A(net276),
    .B(_0547_));
 sg13g2_o21ai_1 _1235_ (.B1(_0551_),
    .Y(_0103_),
    .A1(net162),
    .A2(_0373_));
 sg13g2_nand2_1 _1236_ (.Y(_0552_),
    .A(net449),
    .B(_0547_));
 sg13g2_o21ai_1 _1237_ (.B1(_0552_),
    .Y(_0104_),
    .A1(net162),
    .A2(_0404_));
 sg13g2_nand2_1 _1238_ (.Y(_0553_),
    .A(net413),
    .B(_0547_));
 sg13g2_o21ai_1 _1239_ (.B1(_0553_),
    .Y(_0105_),
    .A1(_0249_),
    .A2(_0432_));
 sg13g2_nand2_1 _1240_ (.Y(_0554_),
    .A(net286),
    .B(_0547_));
 sg13g2_o21ai_1 _1241_ (.B1(_0554_),
    .Y(_0106_),
    .A1(_0249_),
    .A2(_0470_));
 sg13g2_nand2_1 _1242_ (.Y(_0555_),
    .A(net446),
    .B(_0547_));
 sg13g2_o21ai_1 _1243_ (.B1(_0555_),
    .Y(_0107_),
    .A1(net162),
    .A2(_0496_));
 sg13g2_nand3_1 _1244_ (.B(_0218_),
    .C(_0248_),
    .A(net461),
    .Y(_0556_));
 sg13g2_xor2_1 _1245_ (.B(_0249_),
    .A(net461),
    .X(_0557_));
 sg13g2_mux2_1 _1246_ (.A0(_0277_),
    .A1(_0557_),
    .S(_0270_),
    .X(_0558_));
 sg13g2_nor2_1 _1247_ (.A(net191),
    .B(_0558_),
    .Y(_0112_));
 sg13g2_nor2_1 _1248_ (.A(_0180_),
    .B(_0556_),
    .Y(_0559_));
 sg13g2_and2_1 _1249_ (.A(_0180_),
    .B(_0556_),
    .X(_0560_));
 sg13g2_mux2_1 _1250_ (.A0(_0309_),
    .A1(_0560_),
    .S(_0270_),
    .X(_0561_));
 sg13g2_nor3_1 _1251_ (.A(net191),
    .B(_0559_),
    .C(_0561_),
    .Y(_0113_));
 sg13g2_nand2_1 _1252_ (.Y(_0562_),
    .A(net465),
    .B(_0559_));
 sg13g2_and2_1 _1253_ (.A(_0270_),
    .B(_0562_),
    .X(_0563_));
 sg13g2_o21ai_1 _1254_ (.B1(_0563_),
    .Y(_0564_),
    .A1(net465),
    .A2(_0559_));
 sg13g2_o21ai_1 _1255_ (.B1(_0564_),
    .Y(_0565_),
    .A1(_0270_),
    .A2(_0339_));
 sg13g2_and2_1 _1256_ (.A(net192),
    .B(_0565_),
    .X(_0114_));
 sg13g2_nor2_1 _1257_ (.A(net458),
    .B(_0562_),
    .Y(_0566_));
 sg13g2_a21oi_1 _1258_ (.A1(net458),
    .A2(_0563_),
    .Y(_0567_),
    .B1(_0566_));
 sg13g2_o21ai_1 _1259_ (.B1(_0567_),
    .Y(_0568_),
    .A1(_0270_),
    .A2(_0373_));
 sg13g2_and2_1 _1260_ (.A(net192),
    .B(_0568_),
    .X(_0115_));
 sg13g2_and2_1 _1261_ (.A(net193),
    .B(net161),
    .X(_0569_));
 sg13g2_nand2_1 _1262_ (.Y(_0570_),
    .A(net288),
    .B(_0569_));
 sg13g2_o21ai_1 _1263_ (.B1(_0570_),
    .Y(_0116_),
    .A1(_0257_),
    .A2(_0277_));
 sg13g2_nand2_1 _1264_ (.Y(_0571_),
    .A(net293),
    .B(_0569_));
 sg13g2_o21ai_1 _1265_ (.B1(_0571_),
    .Y(_0117_),
    .A1(_0257_),
    .A2(_0309_));
 sg13g2_nand2_1 _1266_ (.Y(_0572_),
    .A(net313),
    .B(_0569_));
 sg13g2_o21ai_1 _1267_ (.B1(_0572_),
    .Y(_0118_),
    .A1(net161),
    .A2(_0339_));
 sg13g2_nand2_1 _1268_ (.Y(_0573_),
    .A(net399),
    .B(_0569_));
 sg13g2_o21ai_1 _1269_ (.B1(_0573_),
    .Y(_0119_),
    .A1(net161),
    .A2(_0373_));
 sg13g2_nand2_1 _1270_ (.Y(_0574_),
    .A(net436),
    .B(_0569_));
 sg13g2_o21ai_1 _1271_ (.B1(_0574_),
    .Y(_0120_),
    .A1(net161),
    .A2(_0404_));
 sg13g2_nand2_1 _1272_ (.Y(_0575_),
    .A(net306),
    .B(_0569_));
 sg13g2_o21ai_1 _1273_ (.B1(_0575_),
    .Y(_0121_),
    .A1(net161),
    .A2(_0432_));
 sg13g2_nand2_1 _1274_ (.Y(_0576_),
    .A(net309),
    .B(_0569_));
 sg13g2_o21ai_1 _1275_ (.B1(_0576_),
    .Y(_0122_),
    .A1(net161),
    .A2(_0470_));
 sg13g2_nand2_1 _1276_ (.Y(_0577_),
    .A(net408),
    .B(_0569_));
 sg13g2_o21ai_1 _1277_ (.B1(_0577_),
    .Y(_0123_),
    .A1(net161),
    .A2(_0496_));
 sg13g2_or2_1 _1278_ (.X(_0578_),
    .B(_0506_),
    .A(_0215_));
 sg13g2_mux2_1 _1279_ (.A0(net146),
    .A1(net360),
    .S(_0578_),
    .X(_0124_));
 sg13g2_mux2_1 _1280_ (.A0(net142),
    .A1(net319),
    .S(_0578_),
    .X(_0125_));
 sg13g2_mux2_1 _1281_ (.A0(net141),
    .A1(net375),
    .S(_0578_),
    .X(_0126_));
 sg13g2_mux2_1 _1282_ (.A0(net139),
    .A1(net435),
    .S(_0578_),
    .X(_0127_));
 sg13g2_mux2_1 _1283_ (.A0(net137),
    .A1(net361),
    .S(_0578_),
    .X(_0128_));
 sg13g2_mux2_1 _1284_ (.A0(net133),
    .A1(net388),
    .S(_0578_),
    .X(_0129_));
 sg13g2_mux2_1 _1285_ (.A0(net135),
    .A1(net406),
    .S(_0578_),
    .X(_0130_));
 sg13g2_mux2_1 _1286_ (.A0(net131),
    .A1(net382),
    .S(_0578_),
    .X(_0131_));
 sg13g2_or2_1 _1287_ (.X(_0579_),
    .B(_0514_),
    .A(_0215_));
 sg13g2_mux2_1 _1288_ (.A0(_0279_),
    .A1(net434),
    .S(net149),
    .X(_0132_));
 sg13g2_mux2_1 _1289_ (.A0(net142),
    .A1(net433),
    .S(net149),
    .X(_0133_));
 sg13g2_mux2_1 _1290_ (.A0(_0340_),
    .A1(net407),
    .S(net149),
    .X(_0134_));
 sg13g2_nor2_1 _1291_ (.A(net139),
    .B(net149),
    .Y(_0580_));
 sg13g2_a21oi_1 _1292_ (.A1(_0193_),
    .A2(net149),
    .Y(_0135_),
    .B1(_0580_));
 sg13g2_mux2_1 _1293_ (.A0(net137),
    .A1(net447),
    .S(net149),
    .X(_0136_));
 sg13g2_mux2_1 _1294_ (.A0(net133),
    .A1(net420),
    .S(net149),
    .X(_0137_));
 sg13g2_mux2_1 _1295_ (.A0(net135),
    .A1(net317),
    .S(_0579_),
    .X(_0138_));
 sg13g2_mux2_1 _1296_ (.A0(net131),
    .A1(net318),
    .S(net149),
    .X(_0139_));
 sg13g2_nor2b_2 _1297_ (.A(_0213_),
    .B_N(_0214_),
    .Y(_0581_));
 sg13g2_nand3_1 _1298_ (.B(_0505_),
    .C(_0581_),
    .A(_0211_),
    .Y(_0582_));
 sg13g2_mux2_1 _1299_ (.A0(net145),
    .A1(net323),
    .S(_0582_),
    .X(_0140_));
 sg13g2_mux2_1 _1300_ (.A0(net143),
    .A1(net430),
    .S(_0582_),
    .X(_0141_));
 sg13g2_mux2_1 _1301_ (.A0(net140),
    .A1(net438),
    .S(_0582_),
    .X(_0142_));
 sg13g2_mux2_1 _1302_ (.A0(net138),
    .A1(net427),
    .S(_0582_),
    .X(_0143_));
 sg13g2_mux2_1 _1303_ (.A0(net136),
    .A1(net448),
    .S(_0582_),
    .X(_0144_));
 sg13g2_mux2_1 _1304_ (.A0(net132),
    .A1(net419),
    .S(_0582_),
    .X(_0145_));
 sg13g2_mux2_1 _1305_ (.A0(net134),
    .A1(net415),
    .S(_0582_),
    .X(_0146_));
 sg13g2_mux2_1 _1306_ (.A0(net130),
    .A1(net424),
    .S(_0582_),
    .X(_0147_));
 sg13g2_nand2_1 _1307_ (.Y(_0583_),
    .A(_0515_),
    .B(_0581_));
 sg13g2_mux2_1 _1308_ (.A0(net145),
    .A1(net370),
    .S(net147),
    .X(_0148_));
 sg13g2_mux2_1 _1309_ (.A0(net143),
    .A1(net403),
    .S(net147),
    .X(_0149_));
 sg13g2_mux2_1 _1310_ (.A0(net140),
    .A1(net321),
    .S(net147),
    .X(_0150_));
 sg13g2_mux2_1 _1311_ (.A0(net138),
    .A1(net387),
    .S(net147),
    .X(_0151_));
 sg13g2_mux2_1 _1312_ (.A0(net136),
    .A1(net328),
    .S(net147),
    .X(_0152_));
 sg13g2_mux2_1 _1313_ (.A0(net132),
    .A1(net340),
    .S(net147),
    .X(_0153_));
 sg13g2_nor2_1 _1314_ (.A(net134),
    .B(net147),
    .Y(_0584_));
 sg13g2_a21oi_1 _1315_ (.A1(_0196_),
    .A2(_0583_),
    .Y(_0154_),
    .B1(_0584_));
 sg13g2_mux2_1 _1316_ (.A0(net130),
    .A1(net366),
    .S(net147),
    .X(_0155_));
 sg13g2_nand3_1 _1317_ (.B(_0505_),
    .C(_0513_),
    .A(_0210_),
    .Y(_0585_));
 sg13g2_mux2_1 _1318_ (.A0(net145),
    .A1(net390),
    .S(_0585_),
    .X(_0156_));
 sg13g2_mux2_1 _1319_ (.A0(net142),
    .A1(net308),
    .S(_0585_),
    .X(_0157_));
 sg13g2_mux2_1 _1320_ (.A0(net140),
    .A1(net385),
    .S(_0585_),
    .X(_0158_));
 sg13g2_mux2_1 _1321_ (.A0(net138),
    .A1(net381),
    .S(_0585_),
    .X(_0159_));
 sg13g2_mux2_1 _1322_ (.A0(net136),
    .A1(net315),
    .S(_0585_),
    .X(_0160_));
 sg13g2_mux2_1 _1323_ (.A0(net132),
    .A1(net421),
    .S(_0585_),
    .X(_0161_));
 sg13g2_mux2_1 _1324_ (.A0(net134),
    .A1(net394),
    .S(_0585_),
    .X(_0162_));
 sg13g2_mux2_1 _1325_ (.A0(net130),
    .A1(net428),
    .S(_0585_),
    .X(_0163_));
 sg13g2_nand3_1 _1326_ (.B(_0505_),
    .C(_0581_),
    .A(_0210_),
    .Y(_0586_));
 sg13g2_mux2_1 _1327_ (.A0(net145),
    .A1(net397),
    .S(_0586_),
    .X(_0164_));
 sg13g2_mux2_1 _1328_ (.A0(net143),
    .A1(net389),
    .S(_0586_),
    .X(_0165_));
 sg13g2_mux2_1 _1329_ (.A0(net141),
    .A1(net395),
    .S(_0586_),
    .X(_0166_));
 sg13g2_mux2_1 _1330_ (.A0(net138),
    .A1(net402),
    .S(_0586_),
    .X(_0167_));
 sg13g2_mux2_1 _1331_ (.A0(net136),
    .A1(net418),
    .S(_0586_),
    .X(_0168_));
 sg13g2_mux2_1 _1332_ (.A0(net132),
    .A1(net440),
    .S(_0586_),
    .X(_0169_));
 sg13g2_mux2_1 _1333_ (.A0(net134),
    .A1(net350),
    .S(_0586_),
    .X(_0170_));
 sg13g2_mux2_1 _1334_ (.A0(net130),
    .A1(net326),
    .S(_0586_),
    .X(_0171_));
 sg13g2_nand3_1 _1335_ (.B(_0210_),
    .C(_0581_),
    .A(_0208_),
    .Y(_0587_));
 sg13g2_mux2_1 _1336_ (.A0(net146),
    .A1(net338),
    .S(_0587_),
    .X(_0172_));
 sg13g2_mux2_1 _1337_ (.A0(net143),
    .A1(net416),
    .S(_0587_),
    .X(_0173_));
 sg13g2_mux2_1 _1338_ (.A0(net141),
    .A1(net346),
    .S(_0587_),
    .X(_0174_));
 sg13g2_mux2_1 _1339_ (.A0(net138),
    .A1(net339),
    .S(_0587_),
    .X(_0175_));
 sg13g2_mux2_1 _1340_ (.A0(net136),
    .A1(net439),
    .S(_0587_),
    .X(_0176_));
 sg13g2_mux2_1 _1341_ (.A0(net132),
    .A1(net330),
    .S(_0587_),
    .X(_0177_));
 sg13g2_mux2_1 _1342_ (.A0(net134),
    .A1(net354),
    .S(_0587_),
    .X(_0178_));
 sg13g2_mux2_1 _1343_ (.A0(net130),
    .A1(net417),
    .S(_0587_),
    .X(_0179_));
 sg13g2_a21oi_1 _1344_ (.A1(_0277_),
    .A2(net153),
    .Y(_0108_),
    .B1(_0500_));
 sg13g2_a21oi_1 _1345_ (.A1(_0309_),
    .A2(net152),
    .Y(_0109_),
    .B1(_0501_));
 sg13g2_a21oi_1 _1346_ (.A1(_0339_),
    .A2(net153),
    .Y(_0110_),
    .B1(_0502_));
 sg13g2_a21oi_1 _1347_ (.A1(_0373_),
    .A2(net153),
    .Y(_0111_),
    .B1(_0503_));
 sg13g2_dfrbpq_1 _1348_ (.RESET_B(net40),
    .D(_0004_),
    .Q(\cpu0.ram[5][0] ),
    .CLK(clknet_5_16__leaf_clk));
 sg13g2_dfrbpq_1 _1349_ (.RESET_B(net263),
    .D(_0005_),
    .Q(\cpu0.ram[5][1] ),
    .CLK(clknet_5_5__leaf_clk));
 sg13g2_dfrbpq_1 _1350_ (.RESET_B(net262),
    .D(_0006_),
    .Q(\cpu0.ram[5][2] ),
    .CLK(clknet_5_16__leaf_clk));
 sg13g2_dfrbpq_1 _1351_ (.RESET_B(net261),
    .D(_0007_),
    .Q(\cpu0.ram[5][3] ),
    .CLK(clknet_5_17__leaf_clk));
 sg13g2_dfrbpq_1 _1352_ (.RESET_B(net260),
    .D(_0008_),
    .Q(\cpu0.ram[5][4] ),
    .CLK(clknet_5_16__leaf_clk));
 sg13g2_dfrbpq_1 _1353_ (.RESET_B(net259),
    .D(_0009_),
    .Q(\cpu0.ram[5][5] ),
    .CLK(clknet_5_20__leaf_clk));
 sg13g2_dfrbpq_1 _1354_ (.RESET_B(net258),
    .D(_0010_),
    .Q(\cpu0.ram[5][6] ),
    .CLK(clknet_5_20__leaf_clk));
 sg13g2_dfrbpq_1 _1355_ (.RESET_B(net257),
    .D(_0011_),
    .Q(\cpu0.ram[5][7] ),
    .CLK(clknet_5_17__leaf_clk));
 sg13g2_dfrbpq_1 _1356_ (.RESET_B(net256),
    .D(_0012_),
    .Q(_0000_),
    .CLK(clknet_5_25__leaf_clk));
 sg13g2_dfrbpq_1 _1357_ (.RESET_B(net255),
    .D(_0013_),
    .Q(_0001_),
    .CLK(clknet_5_30__leaf_clk));
 sg13g2_dfrbpq_1 _1358_ (.RESET_B(net254),
    .D(net455),
    .Q(_0002_),
    .CLK(clknet_5_31__leaf_clk));
 sg13g2_dfrbpq_2 _1359_ (.RESET_B(net253),
    .D(net453),
    .Q(_0003_),
    .CLK(clknet_5_25__leaf_clk));
 sg13g2_dfrbpq_1 _1360_ (.RESET_B(net252),
    .D(_0016_),
    .Q(\cpu0.ram[14][0] ),
    .CLK(clknet_5_22__leaf_clk));
 sg13g2_dfrbpq_1 _1361_ (.RESET_B(net251),
    .D(_0017_),
    .Q(\cpu0.ram[14][1] ),
    .CLK(clknet_5_22__leaf_clk));
 sg13g2_dfrbpq_1 _1362_ (.RESET_B(net250),
    .D(_0018_),
    .Q(\cpu0.ram[14][2] ),
    .CLK(clknet_5_22__leaf_clk));
 sg13g2_dfrbpq_1 _1363_ (.RESET_B(net249),
    .D(_0019_),
    .Q(\cpu0.ram[14][3] ),
    .CLK(clknet_5_23__leaf_clk));
 sg13g2_dfrbpq_1 _1364_ (.RESET_B(net248),
    .D(_0020_),
    .Q(\cpu0.ram[14][4] ),
    .CLK(clknet_5_28__leaf_clk));
 sg13g2_dfrbpq_1 _1365_ (.RESET_B(net247),
    .D(_0021_),
    .Q(\cpu0.ram[14][5] ),
    .CLK(clknet_5_22__leaf_clk));
 sg13g2_dfrbpq_1 _1366_ (.RESET_B(net246),
    .D(_0022_),
    .Q(\cpu0.ram[14][6] ),
    .CLK(clknet_5_23__leaf_clk));
 sg13g2_dfrbpq_1 _1367_ (.RESET_B(net245),
    .D(_0023_),
    .Q(\cpu0.ram[14][7] ),
    .CLK(clknet_5_19__leaf_clk));
 sg13g2_dfrbpq_1 _1368_ (.RESET_B(net244),
    .D(_0024_),
    .Q(\cpu0.ram[13][0] ),
    .CLK(clknet_5_29__leaf_clk));
 sg13g2_dfrbpq_1 _1369_ (.RESET_B(net243),
    .D(_0025_),
    .Q(\cpu0.ram[13][1] ),
    .CLK(clknet_5_28__leaf_clk));
 sg13g2_dfrbpq_1 _1370_ (.RESET_B(net242),
    .D(_0026_),
    .Q(\cpu0.ram[13][2] ),
    .CLK(clknet_5_24__leaf_clk));
 sg13g2_dfrbpq_1 _1371_ (.RESET_B(net241),
    .D(_0027_),
    .Q(\cpu0.ram[13][3] ),
    .CLK(clknet_5_30__leaf_clk));
 sg13g2_dfrbpq_1 _1372_ (.RESET_B(net240),
    .D(_0028_),
    .Q(\cpu0.ram[13][4] ),
    .CLK(clknet_5_25__leaf_clk));
 sg13g2_dfrbpq_1 _1373_ (.RESET_B(net239),
    .D(_0029_),
    .Q(\cpu0.ram[13][5] ),
    .CLK(clknet_5_19__leaf_clk));
 sg13g2_dfrbpq_1 _1374_ (.RESET_B(net238),
    .D(_0030_),
    .Q(\cpu0.ram[13][6] ),
    .CLK(clknet_5_29__leaf_clk));
 sg13g2_dfrbpq_1 _1375_ (.RESET_B(net237),
    .D(_0031_),
    .Q(\cpu0.ram[13][7] ),
    .CLK(clknet_5_24__leaf_clk));
 sg13g2_dfrbpq_2 _1376_ (.RESET_B(net236),
    .D(_0032_),
    .Q(\cpu0.step[1] ),
    .CLK(clknet_5_30__leaf_clk));
 sg13g2_dfrbpq_2 _1377_ (.RESET_B(net235),
    .D(net460),
    .Q(\cpu0.step[2] ),
    .CLK(clknet_5_31__leaf_clk));
 sg13g2_dfrbpq_1 _1378_ (.RESET_B(net234),
    .D(_0034_),
    .Q(\cpu0.ram[12][0] ),
    .CLK(clknet_5_28__leaf_clk));
 sg13g2_dfrbpq_1 _1379_ (.RESET_B(net233),
    .D(_0035_),
    .Q(\cpu0.ram[12][1] ),
    .CLK(clknet_5_28__leaf_clk));
 sg13g2_dfrbpq_1 _1380_ (.RESET_B(net232),
    .D(_0036_),
    .Q(\cpu0.ram[12][2] ),
    .CLK(clknet_5_18__leaf_clk));
 sg13g2_dfrbpq_1 _1381_ (.RESET_B(net231),
    .D(_0037_),
    .Q(\cpu0.ram[12][3] ),
    .CLK(clknet_5_29__leaf_clk));
 sg13g2_dfrbpq_1 _1382_ (.RESET_B(net230),
    .D(_0038_),
    .Q(\cpu0.ram[12][4] ),
    .CLK(clknet_5_24__leaf_clk));
 sg13g2_dfrbpq_1 _1383_ (.RESET_B(net229),
    .D(_0039_),
    .Q(\cpu0.ram[12][5] ),
    .CLK(clknet_5_19__leaf_clk));
 sg13g2_dfrbpq_1 _1384_ (.RESET_B(net228),
    .D(_0040_),
    .Q(\cpu0.ram[12][6] ),
    .CLK(clknet_5_28__leaf_clk));
 sg13g2_dfrbpq_1 _1385_ (.RESET_B(net227),
    .D(_0041_),
    .Q(\cpu0.ram[12][7] ),
    .CLK(clknet_5_24__leaf_clk));
 sg13g2_dfrbpq_2 _1386_ (.RESET_B(net226),
    .D(_0042_),
    .Q(\cpu0.step[0] ),
    .CLK(clknet_5_30__leaf_clk));
 sg13g2_dfrbpq_1 _1387_ (.RESET_B(net225),
    .D(_0043_),
    .Q(\cpu0.ram[4][0] ),
    .CLK(clknet_5_5__leaf_clk));
 sg13g2_dfrbpq_1 _1388_ (.RESET_B(net224),
    .D(_0044_),
    .Q(\cpu0.ram[4][1] ),
    .CLK(clknet_5_5__leaf_clk));
 sg13g2_dfrbpq_1 _1389_ (.RESET_B(net223),
    .D(_0045_),
    .Q(\cpu0.ram[4][2] ),
    .CLK(clknet_5_5__leaf_clk));
 sg13g2_dfrbpq_1 _1390_ (.RESET_B(net222),
    .D(_0046_),
    .Q(\cpu0.ram[4][3] ),
    .CLK(clknet_5_17__leaf_clk));
 sg13g2_dfrbpq_1 _1391_ (.RESET_B(net221),
    .D(_0047_),
    .Q(\cpu0.ram[4][4] ),
    .CLK(clknet_5_18__leaf_clk));
 sg13g2_dfrbpq_1 _1392_ (.RESET_B(net220),
    .D(_0048_),
    .Q(\cpu0.ram[4][5] ),
    .CLK(clknet_5_20__leaf_clk));
 sg13g2_dfrbpq_1 _1393_ (.RESET_B(net219),
    .D(_0049_),
    .Q(\cpu0.ram[4][6] ),
    .CLK(clknet_5_20__leaf_clk));
 sg13g2_dfrbpq_1 _1394_ (.RESET_B(net218),
    .D(_0050_),
    .Q(\cpu0.ram[4][7] ),
    .CLK(clknet_5_17__leaf_clk));
 sg13g2_dfrbpq_1 _1395_ (.RESET_B(net217),
    .D(_0051_),
    .Q(\cpu0.ram[3][0] ),
    .CLK(clknet_5_4__leaf_clk));
 sg13g2_dfrbpq_1 _1396_ (.RESET_B(net216),
    .D(_0052_),
    .Q(\cpu0.ram[3][1] ),
    .CLK(clknet_5_4__leaf_clk));
 sg13g2_dfrbpq_1 _1397_ (.RESET_B(net215),
    .D(_0053_),
    .Q(\cpu0.ram[3][2] ),
    .CLK(clknet_5_7__leaf_clk));
 sg13g2_dfrbpq_1 _1398_ (.RESET_B(net214),
    .D(_0054_),
    .Q(\cpu0.ram[3][3] ),
    .CLK(clknet_5_7__leaf_clk));
 sg13g2_dfrbpq_1 _1399_ (.RESET_B(net213),
    .D(_0055_),
    .Q(\cpu0.ram[3][4] ),
    .CLK(clknet_5_1__leaf_clk));
 sg13g2_dfrbpq_1 _1400_ (.RESET_B(net212),
    .D(_0056_),
    .Q(\cpu0.ram[3][5] ),
    .CLK(clknet_5_1__leaf_clk));
 sg13g2_dfrbpq_1 _1401_ (.RESET_B(net211),
    .D(_0057_),
    .Q(\cpu0.ram[3][6] ),
    .CLK(clknet_5_3__leaf_clk));
 sg13g2_dfrbpq_1 _1402_ (.RESET_B(net210),
    .D(_0058_),
    .Q(\cpu0.ram[3][7] ),
    .CLK(clknet_5_1__leaf_clk));
 sg13g2_dfrbpq_1 _1403_ (.RESET_B(net209),
    .D(_0059_),
    .Q(\cpu0.ram[2][0] ),
    .CLK(clknet_5_4__leaf_clk));
 sg13g2_dfrbpq_1 _1404_ (.RESET_B(net208),
    .D(_0060_),
    .Q(\cpu0.ram[2][1] ),
    .CLK(clknet_5_5__leaf_clk));
 sg13g2_dfrbpq_1 _1405_ (.RESET_B(net207),
    .D(_0061_),
    .Q(\cpu0.ram[2][2] ),
    .CLK(clknet_5_7__leaf_clk));
 sg13g2_dfrbpq_1 _1406_ (.RESET_B(net206),
    .D(_0062_),
    .Q(\cpu0.ram[2][3] ),
    .CLK(clknet_5_6__leaf_clk));
 sg13g2_dfrbpq_1 _1407_ (.RESET_B(net205),
    .D(_0063_),
    .Q(\cpu0.ram[2][4] ),
    .CLK(clknet_5_2__leaf_clk));
 sg13g2_dfrbpq_1 _1408_ (.RESET_B(net204),
    .D(_0064_),
    .Q(\cpu0.ram[2][5] ),
    .CLK(clknet_5_0__leaf_clk));
 sg13g2_dfrbpq_1 _1409_ (.RESET_B(net203),
    .D(_0065_),
    .Q(\cpu0.ram[2][6] ),
    .CLK(clknet_5_6__leaf_clk));
 sg13g2_dfrbpq_1 _1410_ (.RESET_B(net202),
    .D(_0066_),
    .Q(\cpu0.ram[2][7] ),
    .CLK(clknet_5_0__leaf_clk));
 sg13g2_dfrbpq_1 _1411_ (.RESET_B(net201),
    .D(_0067_),
    .Q(\cpu0.ram[1][0] ),
    .CLK(clknet_5_4__leaf_clk));
 sg13g2_dfrbpq_1 _1412_ (.RESET_B(net200),
    .D(_0068_),
    .Q(\cpu0.ram[1][1] ),
    .CLK(clknet_5_4__leaf_clk));
 sg13g2_dfrbpq_1 _1413_ (.RESET_B(net199),
    .D(_0069_),
    .Q(\cpu0.ram[1][2] ),
    .CLK(clknet_5_7__leaf_clk));
 sg13g2_dfrbpq_1 _1414_ (.RESET_B(net198),
    .D(_0070_),
    .Q(\cpu0.ram[1][3] ),
    .CLK(clknet_5_6__leaf_clk));
 sg13g2_dfrbpq_1 _1415_ (.RESET_B(net197),
    .D(_0071_),
    .Q(\cpu0.ram[1][4] ),
    .CLK(clknet_5_2__leaf_clk));
 sg13g2_dfrbpq_1 _1416_ (.RESET_B(net196),
    .D(_0072_),
    .Q(\cpu0.ram[1][5] ),
    .CLK(clknet_5_0__leaf_clk));
 sg13g2_dfrbpq_1 _1417_ (.RESET_B(net195),
    .D(_0073_),
    .Q(\cpu0.ram[1][6] ),
    .CLK(clknet_5_3__leaf_clk));
 sg13g2_dfrbpq_1 _1418_ (.RESET_B(net194),
    .D(_0074_),
    .Q(\cpu0.ram[1][7] ),
    .CLK(clknet_5_1__leaf_clk));
 sg13g2_dfrbpq_1 _1419_ (.RESET_B(net129),
    .D(_0075_),
    .Q(\cpu0.ram[15][0] ),
    .CLK(clknet_5_29__leaf_clk));
 sg13g2_dfrbpq_1 _1420_ (.RESET_B(net128),
    .D(_0076_),
    .Q(\cpu0.ram[15][1] ),
    .CLK(clknet_5_22__leaf_clk));
 sg13g2_dfrbpq_1 _1421_ (.RESET_B(net127),
    .D(_0077_),
    .Q(\cpu0.ram[15][2] ),
    .CLK(clknet_5_19__leaf_clk));
 sg13g2_dfrbpq_1 _1422_ (.RESET_B(net126),
    .D(_0078_),
    .Q(\cpu0.ram[15][3] ),
    .CLK(clknet_5_29__leaf_clk));
 sg13g2_dfrbpq_1 _1423_ (.RESET_B(net125),
    .D(_0079_),
    .Q(\cpu0.ram[15][4] ),
    .CLK(clknet_5_28__leaf_clk));
 sg13g2_dfrbpq_1 _1424_ (.RESET_B(net124),
    .D(_0080_),
    .Q(\cpu0.ram[15][5] ),
    .CLK(clknet_5_18__leaf_clk));
 sg13g2_dfrbpq_1 _1425_ (.RESET_B(net123),
    .D(_0081_),
    .Q(\cpu0.ram[15][6] ),
    .CLK(clknet_5_22__leaf_clk));
 sg13g2_dfrbpq_1 _1426_ (.RESET_B(net122),
    .D(_0082_),
    .Q(\cpu0.ram[15][7] ),
    .CLK(clknet_5_18__leaf_clk));
 sg13g2_dfrbpq_1 _1427_ (.RESET_B(net121),
    .D(_0083_),
    .Q(\cpu0.zero_flag ),
    .CLK(clknet_5_27__leaf_clk));
 sg13g2_dfrbpq_2 _1428_ (.RESET_B(net119),
    .D(net348),
    .Q(\cpu0.b_reg[0] ),
    .CLK(clknet_5_26__leaf_clk));
 sg13g2_dfrbpq_1 _1429_ (.RESET_B(net117),
    .D(net296),
    .Q(\cpu0.b_reg[1] ),
    .CLK(clknet_5_15__leaf_clk));
 sg13g2_dfrbpq_2 _1430_ (.RESET_B(net115),
    .D(net284),
    .Q(\cpu0.b_reg[2] ),
    .CLK(clknet_5_11__leaf_clk));
 sg13g2_dfrbpq_2 _1431_ (.RESET_B(net113),
    .D(_0087_),
    .Q(\cpu0.b_reg[3] ),
    .CLK(clknet_5_11__leaf_clk));
 sg13g2_dfrbpq_1 _1432_ (.RESET_B(net111),
    .D(net273),
    .Q(\cpu0.b_reg[4] ),
    .CLK(clknet_5_11__leaf_clk));
 sg13g2_dfrbpq_1 _1433_ (.RESET_B(net109),
    .D(net373),
    .Q(\cpu0.b_reg[5] ),
    .CLK(clknet_5_14__leaf_clk));
 sg13g2_dfrbpq_1 _1434_ (.RESET_B(net107),
    .D(net305),
    .Q(\cpu0.b_reg[6] ),
    .CLK(clknet_5_14__leaf_clk));
 sg13g2_dfrbpq_1 _1435_ (.RESET_B(net105),
    .D(net279),
    .Q(\cpu0.b_reg[7] ),
    .CLK(clknet_5_10__leaf_clk));
 sg13g2_dfrbpq_2 _1436_ (.RESET_B(net103),
    .D(_0092_),
    .Q(\cpu0.a_reg[0] ),
    .CLK(clknet_5_15__leaf_clk));
 sg13g2_dfrbpq_2 _1437_ (.RESET_B(net101),
    .D(_0093_),
    .Q(\cpu0.a_reg[1] ),
    .CLK(clknet_5_14__leaf_clk));
 sg13g2_dfrbpq_2 _1438_ (.RESET_B(net99),
    .D(_0094_),
    .Q(\cpu0.a_reg[2] ),
    .CLK(clknet_5_15__leaf_clk));
 sg13g2_dfrbpq_2 _1439_ (.RESET_B(net97),
    .D(_0095_),
    .Q(\cpu0.a_reg[3] ),
    .CLK(clknet_5_14__leaf_clk));
 sg13g2_dfrbpq_2 _1440_ (.RESET_B(net95),
    .D(net299),
    .Q(\cpu0.a_reg[4] ),
    .CLK(clknet_5_14__leaf_clk));
 sg13g2_dfrbpq_2 _1441_ (.RESET_B(net93),
    .D(net405),
    .Q(\cpu0.a_reg[5] ),
    .CLK(clknet_5_14__leaf_clk));
 sg13g2_dfrbpq_2 _1442_ (.RESET_B(net91),
    .D(net334),
    .Q(\cpu0.a_reg[6] ),
    .CLK(clknet_5_11__leaf_clk));
 sg13g2_dfrbpq_2 _1443_ (.RESET_B(net89),
    .D(net291),
    .Q(\cpu0.a_reg[7] ),
    .CLK(clknet_5_11__leaf_clk));
 sg13g2_dfrbpq_1 _1444_ (.RESET_B(net87),
    .D(_0100_),
    .Q(\cpu0.ir[0] ),
    .CLK(clknet_5_26__leaf_clk));
 sg13g2_dfrbpq_1 _1445_ (.RESET_B(net85),
    .D(_0101_),
    .Q(\cpu0.ir[1] ),
    .CLK(clknet_5_26__leaf_clk));
 sg13g2_dfrbpq_1 _1446_ (.RESET_B(net83),
    .D(_0102_),
    .Q(\cpu0.ir[2] ),
    .CLK(clknet_5_27__leaf_clk));
 sg13g2_dfrbpq_1 _1447_ (.RESET_B(net81),
    .D(_0103_),
    .Q(\cpu0.ir[3] ),
    .CLK(clknet_5_26__leaf_clk));
 sg13g2_dfrbpq_2 _1448_ (.RESET_B(net79),
    .D(_0104_),
    .Q(\cpu0.ir[4] ),
    .CLK(clknet_5_26__leaf_clk));
 sg13g2_dfrbpq_2 _1449_ (.RESET_B(net77),
    .D(net414),
    .Q(\cpu0.ir[5] ),
    .CLK(clknet_5_27__leaf_clk));
 sg13g2_dfrbpq_2 _1450_ (.RESET_B(net75),
    .D(net287),
    .Q(\cpu0.ir[6] ),
    .CLK(clknet_5_27__leaf_clk));
 sg13g2_dfrbpq_2 _1451_ (.RESET_B(net73),
    .D(_0107_),
    .Q(\cpu0.ir[7] ),
    .CLK(clknet_5_26__leaf_clk));
 sg13g2_dfrbpq_1 _1452_ (.RESET_B(net71),
    .D(_0108_),
    .Q(\cpu0.mar[0] ),
    .CLK(clknet_5_25__leaf_clk));
 sg13g2_dfrbpq_2 _1453_ (.RESET_B(net69),
    .D(_0109_),
    .Q(\cpu0.mar[1] ),
    .CLK(clknet_5_30__leaf_clk));
 sg13g2_dfrbpq_1 _1454_ (.RESET_B(net67),
    .D(_0110_),
    .Q(\cpu0.mar[2] ),
    .CLK(clknet_5_27__leaf_clk));
 sg13g2_dfrbpq_1 _1455_ (.RESET_B(net65),
    .D(_0111_),
    .Q(\cpu0.mar[3] ),
    .CLK(clknet_5_25__leaf_clk));
 sg13g2_dfrbpq_2 _1456_ (.RESET_B(net63),
    .D(_0112_),
    .Q(\cpu0.pc[0] ),
    .CLK(clknet_5_31__leaf_clk));
 sg13g2_dfrbpq_1 _1457_ (.RESET_B(net61),
    .D(_0113_),
    .Q(\cpu0.pc[1] ),
    .CLK(clknet_5_31__leaf_clk));
 sg13g2_dfrbpq_1 _1458_ (.RESET_B(net59),
    .D(_0114_),
    .Q(\cpu0.pc[2] ),
    .CLK(clknet_5_30__leaf_clk));
 sg13g2_dfrbpq_2 _1459_ (.RESET_B(net57),
    .D(_0115_),
    .Q(\cpu0.pc[3] ),
    .CLK(clknet_5_31__leaf_clk));
 sg13g2_dfrbpq_1 _1460_ (.RESET_B(net55),
    .D(net289),
    .Q(uo_out[0]),
    .CLK(clknet_5_15__leaf_clk));
 sg13g2_dfrbpq_1 _1461_ (.RESET_B(net53),
    .D(net294),
    .Q(uo_out[1]),
    .CLK(clknet_5_15__leaf_clk));
 sg13g2_dfrbpq_2 _1462_ (.RESET_B(net51),
    .D(net314),
    .Q(uo_out[2]),
    .CLK(clknet_5_10__leaf_clk));
 sg13g2_dfrbpq_2 _1463_ (.RESET_B(net49),
    .D(net400),
    .Q(uo_out[3]),
    .CLK(clknet_5_10__leaf_clk));
 sg13g2_dfrbpq_2 _1464_ (.RESET_B(net47),
    .D(net437),
    .Q(uo_out[4]),
    .CLK(clknet_5_10__leaf_clk));
 sg13g2_dfrbpq_2 _1465_ (.RESET_B(net45),
    .D(net307),
    .Q(uo_out[5]),
    .CLK(clknet_5_10__leaf_clk));
 sg13g2_dfrbpq_2 _1466_ (.RESET_B(net43),
    .D(net310),
    .Q(uo_out[6]),
    .CLK(clknet_5_10__leaf_clk));
 sg13g2_dfrbpq_2 _1467_ (.RESET_B(net41),
    .D(net409),
    .Q(uo_out[7]),
    .CLK(clknet_5_8__leaf_clk));
 sg13g2_dfrbpq_1 _1468_ (.RESET_B(net39),
    .D(_0124_),
    .Q(\cpu0.ram[6][0] ),
    .CLK(clknet_5_21__leaf_clk));
 sg13g2_dfrbpq_1 _1469_ (.RESET_B(net38),
    .D(_0125_),
    .Q(\cpu0.ram[6][1] ),
    .CLK(clknet_5_16__leaf_clk));
 sg13g2_dfrbpq_1 _1470_ (.RESET_B(net37),
    .D(_0126_),
    .Q(\cpu0.ram[6][2] ),
    .CLK(clknet_5_21__leaf_clk));
 sg13g2_dfrbpq_1 _1471_ (.RESET_B(net36),
    .D(_0127_),
    .Q(\cpu0.ram[6][3] ),
    .CLK(clknet_5_23__leaf_clk));
 sg13g2_dfrbpq_1 _1472_ (.RESET_B(net35),
    .D(_0128_),
    .Q(\cpu0.ram[6][4] ),
    .CLK(clknet_5_18__leaf_clk));
 sg13g2_dfrbpq_1 _1473_ (.RESET_B(net34),
    .D(_0129_),
    .Q(\cpu0.ram[6][5] ),
    .CLK(clknet_5_20__leaf_clk));
 sg13g2_dfrbpq_1 _1474_ (.RESET_B(net33),
    .D(_0130_),
    .Q(\cpu0.ram[6][6] ),
    .CLK(clknet_5_21__leaf_clk));
 sg13g2_dfrbpq_1 _1475_ (.RESET_B(net32),
    .D(_0131_),
    .Q(\cpu0.ram[6][7] ),
    .CLK(clknet_5_16__leaf_clk));
 sg13g2_dfrbpq_1 _1476_ (.RESET_B(net31),
    .D(_0132_),
    .Q(\cpu0.ram[7][0] ),
    .CLK(clknet_5_21__leaf_clk));
 sg13g2_dfrbpq_1 _1477_ (.RESET_B(net30),
    .D(_0133_),
    .Q(\cpu0.ram[7][1] ),
    .CLK(clknet_5_16__leaf_clk));
 sg13g2_dfrbpq_1 _1478_ (.RESET_B(net269),
    .D(_0134_),
    .Q(\cpu0.ram[7][2] ),
    .CLK(clknet_5_23__leaf_clk));
 sg13g2_dfrbpq_1 _1479_ (.RESET_B(net268),
    .D(_0135_),
    .Q(\cpu0.ram[7][3] ),
    .CLK(clknet_5_23__leaf_clk));
 sg13g2_dfrbpq_1 _1480_ (.RESET_B(net267),
    .D(_0136_),
    .Q(\cpu0.ram[7][4] ),
    .CLK(clknet_5_19__leaf_clk));
 sg13g2_dfrbpq_1 _1481_ (.RESET_B(net266),
    .D(_0137_),
    .Q(\cpu0.ram[7][5] ),
    .CLK(clknet_5_21__leaf_clk));
 sg13g2_dfrbpq_1 _1482_ (.RESET_B(net265),
    .D(_0138_),
    .Q(\cpu0.ram[7][6] ),
    .CLK(clknet_5_20__leaf_clk));
 sg13g2_dfrbpq_1 _1483_ (.RESET_B(net264),
    .D(_0139_),
    .Q(\cpu0.ram[7][7] ),
    .CLK(clknet_5_17__leaf_clk));
 sg13g2_dfrbpq_1 _1484_ (.RESET_B(net120),
    .D(_0140_),
    .Q(\cpu0.ram[10][0] ),
    .CLK(clknet_5_13__leaf_clk));
 sg13g2_dfrbpq_1 _1485_ (.RESET_B(net118),
    .D(_0141_),
    .Q(\cpu0.ram[10][1] ),
    .CLK(clknet_5_12__leaf_clk));
 sg13g2_dfrbpq_1 _1486_ (.RESET_B(net116),
    .D(_0142_),
    .Q(\cpu0.ram[10][2] ),
    .CLK(clknet_5_6__leaf_clk));
 sg13g2_dfrbpq_1 _1487_ (.RESET_B(net114),
    .D(_0143_),
    .Q(\cpu0.ram[10][3] ),
    .CLK(clknet_5_12__leaf_clk));
 sg13g2_dfrbpq_1 _1488_ (.RESET_B(net112),
    .D(_0144_),
    .Q(\cpu0.ram[10][4] ),
    .CLK(clknet_5_8__leaf_clk));
 sg13g2_dfrbpq_1 _1489_ (.RESET_B(net110),
    .D(_0145_),
    .Q(\cpu0.ram[10][5] ),
    .CLK(clknet_5_2__leaf_clk));
 sg13g2_dfrbpq_1 _1490_ (.RESET_B(net108),
    .D(_0146_),
    .Q(\cpu0.ram[10][6] ),
    .CLK(clknet_5_13__leaf_clk));
 sg13g2_dfrbpq_1 _1491_ (.RESET_B(net106),
    .D(_0147_),
    .Q(\cpu0.ram[10][7] ),
    .CLK(clknet_5_9__leaf_clk));
 sg13g2_dfrbpq_1 _1492_ (.RESET_B(net104),
    .D(_0148_),
    .Q(\cpu0.ram[11][0] ),
    .CLK(clknet_5_24__leaf_clk));
 sg13g2_dfrbpq_1 _1493_ (.RESET_B(net102),
    .D(_0149_),
    .Q(\cpu0.ram[11][1] ),
    .CLK(clknet_5_12__leaf_clk));
 sg13g2_dfrbpq_1 _1494_ (.RESET_B(net100),
    .D(_0150_),
    .Q(\cpu0.ram[11][2] ),
    .CLK(clknet_5_6__leaf_clk));
 sg13g2_dfrbpq_1 _1495_ (.RESET_B(net98),
    .D(_0151_),
    .Q(\cpu0.ram[11][3] ),
    .CLK(clknet_5_12__leaf_clk));
 sg13g2_dfrbpq_1 _1496_ (.RESET_B(net96),
    .D(_0152_),
    .Q(\cpu0.ram[11][4] ),
    .CLK(clknet_5_8__leaf_clk));
 sg13g2_dfrbpq_1 _1497_ (.RESET_B(net94),
    .D(_0153_),
    .Q(\cpu0.ram[11][5] ),
    .CLK(clknet_5_2__leaf_clk));
 sg13g2_dfrbpq_1 _1498_ (.RESET_B(net92),
    .D(_0154_),
    .Q(\cpu0.ram[11][6] ),
    .CLK(clknet_5_18__leaf_clk));
 sg13g2_dfrbpq_1 _1499_ (.RESET_B(net90),
    .D(_0155_),
    .Q(\cpu0.ram[11][7] ),
    .CLK(clknet_5_9__leaf_clk));
 sg13g2_dfrbpq_1 _1500_ (.RESET_B(net88),
    .D(_0156_),
    .Q(\cpu0.ram[0][0] ),
    .CLK(clknet_5_1__leaf_clk));
 sg13g2_dfrbpq_1 _1501_ (.RESET_B(net86),
    .D(_0157_),
    .Q(\cpu0.ram[0][1] ),
    .CLK(clknet_5_4__leaf_clk));
 sg13g2_dfrbpq_1 _1502_ (.RESET_B(net84),
    .D(_0158_),
    .Q(\cpu0.ram[0][2] ),
    .CLK(clknet_5_7__leaf_clk));
 sg13g2_dfrbpq_1 _1503_ (.RESET_B(net82),
    .D(_0159_),
    .Q(\cpu0.ram[0][3] ),
    .CLK(clknet_5_6__leaf_clk));
 sg13g2_dfrbpq_1 _1504_ (.RESET_B(net80),
    .D(_0160_),
    .Q(\cpu0.ram[0][4] ),
    .CLK(clknet_5_0__leaf_clk));
 sg13g2_dfrbpq_1 _1505_ (.RESET_B(net78),
    .D(_0161_),
    .Q(\cpu0.ram[0][5] ),
    .CLK(clknet_5_0__leaf_clk));
 sg13g2_dfrbpq_1 _1506_ (.RESET_B(net76),
    .D(_0162_),
    .Q(\cpu0.ram[0][6] ),
    .CLK(clknet_5_3__leaf_clk));
 sg13g2_dfrbpq_1 _1507_ (.RESET_B(net74),
    .D(_0163_),
    .Q(\cpu0.ram[0][7] ),
    .CLK(clknet_5_0__leaf_clk));
 sg13g2_dfrbpq_1 _1508_ (.RESET_B(net72),
    .D(_0164_),
    .Q(\cpu0.ram[8][0] ),
    .CLK(clknet_5_13__leaf_clk));
 sg13g2_dfrbpq_1 _1509_ (.RESET_B(net70),
    .D(_0165_),
    .Q(\cpu0.ram[8][1] ),
    .CLK(clknet_5_9__leaf_clk));
 sg13g2_dfrbpq_1 _1510_ (.RESET_B(net68),
    .D(_0166_),
    .Q(\cpu0.ram[8][2] ),
    .CLK(clknet_5_3__leaf_clk));
 sg13g2_dfrbpq_1 _1511_ (.RESET_B(net66),
    .D(_0167_),
    .Q(\cpu0.ram[8][3] ),
    .CLK(clknet_5_12__leaf_clk));
 sg13g2_dfrbpq_1 _1512_ (.RESET_B(net64),
    .D(_0168_),
    .Q(\cpu0.ram[8][4] ),
    .CLK(clknet_5_8__leaf_clk));
 sg13g2_dfrbpq_1 _1513_ (.RESET_B(net62),
    .D(_0169_),
    .Q(\cpu0.ram[8][5] ),
    .CLK(clknet_5_2__leaf_clk));
 sg13g2_dfrbpq_1 _1514_ (.RESET_B(net60),
    .D(_0170_),
    .Q(\cpu0.ram[8][6] ),
    .CLK(clknet_5_13__leaf_clk));
 sg13g2_dfrbpq_1 _1515_ (.RESET_B(net58),
    .D(_0171_),
    .Q(\cpu0.ram[8][7] ),
    .CLK(clknet_5_9__leaf_clk));
 sg13g2_dfrbpq_1 _1516_ (.RESET_B(net56),
    .D(_0172_),
    .Q(\cpu0.ram[9][0] ),
    .CLK(clknet_5_24__leaf_clk));
 sg13g2_dfrbpq_1 _1517_ (.RESET_B(net54),
    .D(_0173_),
    .Q(\cpu0.ram[9][1] ),
    .CLK(clknet_5_9__leaf_clk));
 sg13g2_dfrbpq_1 _1518_ (.RESET_B(net52),
    .D(_0174_),
    .Q(\cpu0.ram[9][2] ),
    .CLK(clknet_5_3__leaf_clk));
 sg13g2_dfrbpq_1 _1519_ (.RESET_B(net50),
    .D(_0175_),
    .Q(\cpu0.ram[9][3] ),
    .CLK(clknet_5_12__leaf_clk));
 sg13g2_dfrbpq_1 _1520_ (.RESET_B(net48),
    .D(_0176_),
    .Q(\cpu0.ram[9][4] ),
    .CLK(clknet_5_8__leaf_clk));
 sg13g2_dfrbpq_1 _1521_ (.RESET_B(net46),
    .D(_0177_),
    .Q(\cpu0.ram[9][5] ),
    .CLK(clknet_5_2__leaf_clk));
 sg13g2_dfrbpq_1 _1522_ (.RESET_B(net44),
    .D(_0178_),
    .Q(\cpu0.ram[9][6] ),
    .CLK(clknet_5_13__leaf_clk));
 sg13g2_dfrbpq_1 _1523_ (.RESET_B(net42),
    .D(_0179_),
    .Q(\cpu0.ram[9][7] ),
    .CLK(clknet_5_8__leaf_clk));
 sg13g2_tiehi _1476__31 (.L_HI(net31));
 sg13g2_tiehi _1475__32 (.L_HI(net32));
 sg13g2_tiehi _1474__33 (.L_HI(net33));
 sg13g2_tiehi _1473__34 (.L_HI(net34));
 sg13g2_tiehi _1472__35 (.L_HI(net35));
 sg13g2_tiehi _1471__36 (.L_HI(net36));
 sg13g2_tiehi _1470__37 (.L_HI(net37));
 sg13g2_tiehi _1469__38 (.L_HI(net38));
 sg13g2_tiehi _1468__39 (.L_HI(net39));
 sg13g2_tiehi _1348__40 (.L_HI(net40));
 sg13g2_tiehi _1467__41 (.L_HI(net41));
 sg13g2_tiehi _1523__42 (.L_HI(net42));
 sg13g2_tiehi _1466__43 (.L_HI(net43));
 sg13g2_tiehi _1522__44 (.L_HI(net44));
 sg13g2_tiehi _1465__45 (.L_HI(net45));
 sg13g2_tiehi _1521__46 (.L_HI(net46));
 sg13g2_tiehi _1464__47 (.L_HI(net47));
 sg13g2_tiehi _1520__48 (.L_HI(net48));
 sg13g2_tiehi _1463__49 (.L_HI(net49));
 sg13g2_tiehi _1519__50 (.L_HI(net50));
 sg13g2_tiehi _1462__51 (.L_HI(net51));
 sg13g2_tiehi _1518__52 (.L_HI(net52));
 sg13g2_tiehi _1461__53 (.L_HI(net53));
 sg13g2_tiehi _1517__54 (.L_HI(net54));
 sg13g2_tiehi _1460__55 (.L_HI(net55));
 sg13g2_tiehi _1516__56 (.L_HI(net56));
 sg13g2_tiehi _1459__57 (.L_HI(net57));
 sg13g2_tiehi _1515__58 (.L_HI(net58));
 sg13g2_tiehi _1458__59 (.L_HI(net59));
 sg13g2_tiehi _1514__60 (.L_HI(net60));
 sg13g2_tiehi _1457__61 (.L_HI(net61));
 sg13g2_tiehi _1513__62 (.L_HI(net62));
 sg13g2_tiehi _1456__63 (.L_HI(net63));
 sg13g2_tiehi _1512__64 (.L_HI(net64));
 sg13g2_tiehi _1455__65 (.L_HI(net65));
 sg13g2_tiehi _1511__66 (.L_HI(net66));
 sg13g2_tiehi _1454__67 (.L_HI(net67));
 sg13g2_tiehi _1510__68 (.L_HI(net68));
 sg13g2_tiehi _1453__69 (.L_HI(net69));
 sg13g2_tiehi _1509__70 (.L_HI(net70));
 sg13g2_tiehi _1452__71 (.L_HI(net71));
 sg13g2_tiehi _1508__72 (.L_HI(net72));
 sg13g2_tiehi _1451__73 (.L_HI(net73));
 sg13g2_tiehi _1507__74 (.L_HI(net74));
 sg13g2_tiehi _1450__75 (.L_HI(net75));
 sg13g2_tiehi _1506__76 (.L_HI(net76));
 sg13g2_tiehi _1449__77 (.L_HI(net77));
 sg13g2_tiehi _1505__78 (.L_HI(net78));
 sg13g2_tiehi _1448__79 (.L_HI(net79));
 sg13g2_tiehi _1504__80 (.L_HI(net80));
 sg13g2_tiehi _1447__81 (.L_HI(net81));
 sg13g2_tiehi _1503__82 (.L_HI(net82));
 sg13g2_tiehi _1446__83 (.L_HI(net83));
 sg13g2_tiehi _1502__84 (.L_HI(net84));
 sg13g2_tiehi _1445__85 (.L_HI(net85));
 sg13g2_tiehi _1501__86 (.L_HI(net86));
 sg13g2_tiehi _1444__87 (.L_HI(net87));
 sg13g2_tiehi _1500__88 (.L_HI(net88));
 sg13g2_tiehi _1443__89 (.L_HI(net89));
 sg13g2_tiehi _1499__90 (.L_HI(net90));
 sg13g2_tiehi _1442__91 (.L_HI(net91));
 sg13g2_tiehi _1498__92 (.L_HI(net92));
 sg13g2_tiehi _1441__93 (.L_HI(net93));
 sg13g2_tiehi _1497__94 (.L_HI(net94));
 sg13g2_tiehi _1440__95 (.L_HI(net95));
 sg13g2_tiehi _1496__96 (.L_HI(net96));
 sg13g2_tiehi _1439__97 (.L_HI(net97));
 sg13g2_tiehi _1495__98 (.L_HI(net98));
 sg13g2_tiehi _1438__99 (.L_HI(net99));
 sg13g2_tiehi _1494__100 (.L_HI(net100));
 sg13g2_tiehi _1437__101 (.L_HI(net101));
 sg13g2_tiehi _1493__102 (.L_HI(net102));
 sg13g2_tiehi _1436__103 (.L_HI(net103));
 sg13g2_tiehi _1492__104 (.L_HI(net104));
 sg13g2_tiehi _1435__105 (.L_HI(net105));
 sg13g2_tiehi _1491__106 (.L_HI(net106));
 sg13g2_tiehi _1434__107 (.L_HI(net107));
 sg13g2_tiehi _1490__108 (.L_HI(net108));
 sg13g2_tiehi _1433__109 (.L_HI(net109));
 sg13g2_tiehi _1489__110 (.L_HI(net110));
 sg13g2_tiehi _1432__111 (.L_HI(net111));
 sg13g2_tiehi _1488__112 (.L_HI(net112));
 sg13g2_tiehi _1431__113 (.L_HI(net113));
 sg13g2_tiehi _1487__114 (.L_HI(net114));
 sg13g2_tiehi _1430__115 (.L_HI(net115));
 sg13g2_tiehi _1486__116 (.L_HI(net116));
 sg13g2_tiehi _1429__117 (.L_HI(net117));
 sg13g2_tiehi _1485__118 (.L_HI(net118));
 sg13g2_tiehi _1428__119 (.L_HI(net119));
 sg13g2_tiehi _1484__120 (.L_HI(net120));
 sg13g2_tiehi _1427__121 (.L_HI(net121));
 sg13g2_tiehi _1426__122 (.L_HI(net122));
 sg13g2_tiehi _1425__123 (.L_HI(net123));
 sg13g2_tiehi _1424__124 (.L_HI(net124));
 sg13g2_tiehi _1423__125 (.L_HI(net125));
 sg13g2_tiehi _1422__126 (.L_HI(net126));
 sg13g2_tiehi _1421__127 (.L_HI(net127));
 sg13g2_tiehi _1420__128 (.L_HI(net128));
 sg13g2_tiehi _1419__129 (.L_HI(net129));
 sg13g2_tiehi _1418__130 (.L_HI(net194));
 sg13g2_tiehi _1417__131 (.L_HI(net195));
 sg13g2_tiehi _1416__132 (.L_HI(net196));
 sg13g2_tiehi _1415__133 (.L_HI(net197));
 sg13g2_tiehi _1414__134 (.L_HI(net198));
 sg13g2_tiehi _1413__135 (.L_HI(net199));
 sg13g2_tiehi _1412__136 (.L_HI(net200));
 sg13g2_tiehi _1411__137 (.L_HI(net201));
 sg13g2_tiehi _1410__138 (.L_HI(net202));
 sg13g2_tiehi _1409__139 (.L_HI(net203));
 sg13g2_tiehi _1408__140 (.L_HI(net204));
 sg13g2_tiehi _1407__141 (.L_HI(net205));
 sg13g2_tiehi _1406__142 (.L_HI(net206));
 sg13g2_tiehi _1405__143 (.L_HI(net207));
 sg13g2_tiehi _1404__144 (.L_HI(net208));
 sg13g2_tiehi _1403__145 (.L_HI(net209));
 sg13g2_tiehi _1402__146 (.L_HI(net210));
 sg13g2_tiehi _1401__147 (.L_HI(net211));
 sg13g2_tiehi _1400__148 (.L_HI(net212));
 sg13g2_tiehi _1399__149 (.L_HI(net213));
 sg13g2_tiehi _1398__150 (.L_HI(net214));
 sg13g2_tiehi _1397__151 (.L_HI(net215));
 sg13g2_tiehi _1396__152 (.L_HI(net216));
 sg13g2_tiehi _1395__153 (.L_HI(net217));
 sg13g2_tiehi _1394__154 (.L_HI(net218));
 sg13g2_tiehi _1393__155 (.L_HI(net219));
 sg13g2_tiehi _1392__156 (.L_HI(net220));
 sg13g2_tiehi _1391__157 (.L_HI(net221));
 sg13g2_tiehi _1390__158 (.L_HI(net222));
 sg13g2_tiehi _1389__159 (.L_HI(net223));
 sg13g2_tiehi _1388__160 (.L_HI(net224));
 sg13g2_tiehi _1387__161 (.L_HI(net225));
 sg13g2_tiehi _1386__162 (.L_HI(net226));
 sg13g2_tiehi _1385__163 (.L_HI(net227));
 sg13g2_tiehi _1384__164 (.L_HI(net228));
 sg13g2_tiehi _1383__165 (.L_HI(net229));
 sg13g2_tiehi _1382__166 (.L_HI(net230));
 sg13g2_tiehi _1381__167 (.L_HI(net231));
 sg13g2_tiehi _1380__168 (.L_HI(net232));
 sg13g2_tiehi _1379__169 (.L_HI(net233));
 sg13g2_tiehi _1378__170 (.L_HI(net234));
 sg13g2_tiehi _1377__171 (.L_HI(net235));
 sg13g2_tiehi _1376__172 (.L_HI(net236));
 sg13g2_tiehi _1375__173 (.L_HI(net237));
 sg13g2_tiehi _1374__174 (.L_HI(net238));
 sg13g2_tiehi _1373__175 (.L_HI(net239));
 sg13g2_tiehi _1372__176 (.L_HI(net240));
 sg13g2_tiehi _1371__177 (.L_HI(net241));
 sg13g2_tiehi _1370__178 (.L_HI(net242));
 sg13g2_tiehi _1369__179 (.L_HI(net243));
 sg13g2_tiehi _1368__180 (.L_HI(net244));
 sg13g2_tiehi _1367__181 (.L_HI(net245));
 sg13g2_tiehi _1366__182 (.L_HI(net246));
 sg13g2_tiehi _1365__183 (.L_HI(net247));
 sg13g2_tiehi _1364__184 (.L_HI(net248));
 sg13g2_tiehi _1363__185 (.L_HI(net249));
 sg13g2_tiehi _1362__186 (.L_HI(net250));
 sg13g2_tiehi _1361__187 (.L_HI(net251));
 sg13g2_tiehi _1360__188 (.L_HI(net252));
 sg13g2_tiehi _1359__189 (.L_HI(net253));
 sg13g2_tiehi _1358__190 (.L_HI(net254));
 sg13g2_tiehi _1357__191 (.L_HI(net255));
 sg13g2_tiehi _1356__192 (.L_HI(net256));
 sg13g2_tiehi _1355__193 (.L_HI(net257));
 sg13g2_tiehi _1354__194 (.L_HI(net258));
 sg13g2_tiehi _1353__195 (.L_HI(net259));
 sg13g2_tiehi _1352__196 (.L_HI(net260));
 sg13g2_tiehi _1351__197 (.L_HI(net261));
 sg13g2_tiehi _1350__198 (.L_HI(net262));
 sg13g2_tiehi _1349__199 (.L_HI(net263));
 sg13g2_tiehi _1483__200 (.L_HI(net264));
 sg13g2_tiehi _1482__201 (.L_HI(net265));
 sg13g2_tiehi _1481__202 (.L_HI(net266));
 sg13g2_tiehi _1480__203 (.L_HI(net267));
 sg13g2_tiehi _1479__204 (.L_HI(net268));
 sg13g2_tiehi _1478__205 (.L_HI(net269));
 sg13g2_buf_8 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_tielo tt_um_dranoel06_SAP1_15 (.L_LO(net15));
 sg13g2_tielo tt_um_dranoel06_SAP1_16 (.L_LO(net16));
 sg13g2_tielo tt_um_dranoel06_SAP1_17 (.L_LO(net17));
 sg13g2_tielo tt_um_dranoel06_SAP1_18 (.L_LO(net18));
 sg13g2_tielo tt_um_dranoel06_SAP1_19 (.L_LO(net19));
 sg13g2_tielo tt_um_dranoel06_SAP1_20 (.L_LO(net20));
 sg13g2_tielo tt_um_dranoel06_SAP1_21 (.L_LO(net21));
 sg13g2_tielo tt_um_dranoel06_SAP1_22 (.L_LO(net22));
 sg13g2_tielo tt_um_dranoel06_SAP1_23 (.L_LO(net23));
 sg13g2_tielo tt_um_dranoel06_SAP1_24 (.L_LO(net24));
 sg13g2_tielo tt_um_dranoel06_SAP1_25 (.L_LO(net25));
 sg13g2_tielo tt_um_dranoel06_SAP1_26 (.L_LO(net26));
 sg13g2_tielo tt_um_dranoel06_SAP1_27 (.L_LO(net27));
 sg13g2_tielo tt_um_dranoel06_SAP1_28 (.L_LO(net28));
 sg13g2_tielo tt_um_dranoel06_SAP1_29 (.L_LO(net29));
 sg13g2_tiehi _1477__30 (.L_HI(net30));
 sg13g2_buf_8 fanout130 (.A(_0498_),
    .X(net130));
 sg13g2_buf_8 fanout131 (.A(_0498_),
    .X(net131));
 sg13g2_buf_8 fanout132 (.A(_0434_),
    .X(net132));
 sg13g2_buf_8 fanout133 (.A(_0434_),
    .X(net133));
 sg13g2_buf_8 fanout134 (.A(_0471_),
    .X(net134));
 sg13g2_buf_8 fanout135 (.A(_0471_),
    .X(net135));
 sg13g2_buf_8 fanout136 (.A(_0406_),
    .X(net136));
 sg13g2_buf_8 fanout137 (.A(_0406_),
    .X(net137));
 sg13g2_buf_8 fanout138 (.A(_0375_),
    .X(net138));
 sg13g2_buf_8 fanout139 (.A(_0375_),
    .X(net139));
 sg13g2_buf_8 fanout140 (.A(net141),
    .X(net140));
 sg13g2_buf_8 fanout141 (.A(_0340_),
    .X(net141));
 sg13g2_buf_8 fanout142 (.A(net144),
    .X(net142));
 sg13g2_buf_1 fanout143 (.A(net144),
    .X(net143));
 sg13g2_buf_8 fanout144 (.A(_0310_),
    .X(net144));
 sg13g2_buf_8 fanout145 (.A(net146),
    .X(net145));
 sg13g2_buf_8 fanout146 (.A(_0279_),
    .X(net146));
 sg13g2_buf_8 fanout147 (.A(_0583_),
    .X(net147));
 sg13g2_buf_8 fanout148 (.A(_0516_),
    .X(net148));
 sg13g2_buf_8 fanout149 (.A(_0579_),
    .X(net149));
 sg13g2_buf_8 fanout150 (.A(_0521_),
    .X(net150));
 sg13g2_buf_8 fanout151 (.A(_0507_),
    .X(net151));
 sg13g2_buf_8 fanout152 (.A(_0499_),
    .X(net152));
 sg13g2_buf_1 fanout153 (.A(_0499_),
    .X(net153));
 sg13g2_buf_8 fanout154 (.A(_0519_),
    .X(net154));
 sg13g2_buf_8 fanout155 (.A(_0252_),
    .X(net155));
 sg13g2_buf_8 fanout156 (.A(_0247_),
    .X(net156));
 sg13g2_buf_8 fanout157 (.A(net160),
    .X(net157));
 sg13g2_buf_1 fanout158 (.A(net160),
    .X(net158));
 sg13g2_buf_8 fanout159 (.A(net160),
    .X(net159));
 sg13g2_buf_2 fanout160 (.A(_0206_),
    .X(net160));
 sg13g2_buf_8 fanout161 (.A(_0257_),
    .X(net161));
 sg13g2_buf_8 fanout162 (.A(_0249_),
    .X(net162));
 sg13g2_buf_8 fanout163 (.A(net164),
    .X(net163));
 sg13g2_buf_8 fanout164 (.A(_0186_),
    .X(net164));
 sg13g2_buf_8 fanout165 (.A(_0184_),
    .X(net165));
 sg13g2_buf_8 fanout166 (.A(net456),
    .X(net166));
 sg13g2_buf_8 fanout167 (.A(net168),
    .X(net167));
 sg13g2_buf_8 fanout168 (.A(_0003_),
    .X(net168));
 sg13g2_buf_8 fanout169 (.A(net170),
    .X(net169));
 sg13g2_buf_8 fanout170 (.A(_0002_),
    .X(net170));
 sg13g2_buf_8 fanout171 (.A(net172),
    .X(net171));
 sg13g2_buf_8 fanout172 (.A(net176),
    .X(net172));
 sg13g2_buf_8 fanout173 (.A(net174),
    .X(net173));
 sg13g2_buf_8 fanout174 (.A(net175),
    .X(net174));
 sg13g2_buf_8 fanout175 (.A(net176),
    .X(net175));
 sg13g2_buf_8 fanout176 (.A(_0001_),
    .X(net176));
 sg13g2_buf_8 fanout177 (.A(net178),
    .X(net177));
 sg13g2_buf_8 fanout178 (.A(net190),
    .X(net178));
 sg13g2_buf_8 fanout179 (.A(net190),
    .X(net179));
 sg13g2_buf_1 fanout180 (.A(net190),
    .X(net180));
 sg13g2_buf_8 fanout181 (.A(net185),
    .X(net181));
 sg13g2_buf_8 fanout182 (.A(net185),
    .X(net182));
 sg13g2_buf_8 fanout183 (.A(net185),
    .X(net183));
 sg13g2_buf_8 fanout184 (.A(net185),
    .X(net184));
 sg13g2_buf_8 fanout185 (.A(net190),
    .X(net185));
 sg13g2_buf_8 fanout186 (.A(net187),
    .X(net186));
 sg13g2_buf_1 fanout187 (.A(net188),
    .X(net187));
 sg13g2_buf_1 fanout188 (.A(net189),
    .X(net188));
 sg13g2_buf_8 fanout189 (.A(net190),
    .X(net189));
 sg13g2_buf_8 fanout190 (.A(_0000_),
    .X(net190));
 sg13g2_buf_8 fanout191 (.A(_0183_),
    .X(net191));
 sg13g2_buf_8 fanout192 (.A(net193),
    .X(net192));
 sg13g2_buf_8 fanout193 (.A(rst_n),
    .X(net193));
 sg13g2_buf_1 input1 (.A(ui_in[0]),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[1]),
    .X(net2));
 sg13g2_buf_1 input3 (.A(ui_in[2]),
    .X(net3));
 sg13g2_buf_1 input4 (.A(ui_in[3]),
    .X(net4));
 sg13g2_buf_1 input5 (.A(ui_in[4]),
    .X(net5));
 sg13g2_buf_1 input6 (.A(ui_in[5]),
    .X(net6));
 sg13g2_buf_1 input7 (.A(ui_in[6]),
    .X(net7));
 sg13g2_buf_1 input8 (.A(ui_in[7]),
    .X(net8));
 sg13g2_buf_1 input9 (.A(uio_in[0]),
    .X(net9));
 sg13g2_buf_1 input10 (.A(uio_in[1]),
    .X(net10));
 sg13g2_buf_1 input11 (.A(uio_in[2]),
    .X(net11));
 sg13g2_buf_1 input12 (.A(uio_in[3]),
    .X(net12));
 sg13g2_buf_1 input13 (.A(uio_in[7]),
    .X(net13));
 sg13g2_tielo tt_um_dranoel06_SAP1_14 (.L_LO(net14));
 sg13g2_buf_8 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sg13g2_buf_8 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sg13g2_buf_8 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sg13g2_buf_8 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sg13g2_buf_8 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sg13g2_buf_8 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sg13g2_buf_8 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sg13g2_buf_8 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sg13g2_buf_8 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sg13g2_buf_8 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sg13g2_buf_8 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sg13g2_buf_8 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sg13g2_buf_8 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sg13g2_buf_8 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sg13g2_buf_8 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sg13g2_buf_8 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sg13g2_buf_8 clkbuf_5_0__f_clk (.A(clknet_4_0_0_clk),
    .X(clknet_5_0__leaf_clk));
 sg13g2_buf_8 clkbuf_5_1__f_clk (.A(clknet_4_0_0_clk),
    .X(clknet_5_1__leaf_clk));
 sg13g2_buf_8 clkbuf_5_2__f_clk (.A(clknet_4_1_0_clk),
    .X(clknet_5_2__leaf_clk));
 sg13g2_buf_8 clkbuf_5_3__f_clk (.A(clknet_4_1_0_clk),
    .X(clknet_5_3__leaf_clk));
 sg13g2_buf_8 clkbuf_5_4__f_clk (.A(clknet_4_2_0_clk),
    .X(clknet_5_4__leaf_clk));
 sg13g2_buf_8 clkbuf_5_5__f_clk (.A(clknet_4_2_0_clk),
    .X(clknet_5_5__leaf_clk));
 sg13g2_buf_8 clkbuf_5_6__f_clk (.A(clknet_4_3_0_clk),
    .X(clknet_5_6__leaf_clk));
 sg13g2_buf_8 clkbuf_5_7__f_clk (.A(clknet_4_3_0_clk),
    .X(clknet_5_7__leaf_clk));
 sg13g2_buf_8 clkbuf_5_8__f_clk (.A(clknet_4_4_0_clk),
    .X(clknet_5_8__leaf_clk));
 sg13g2_buf_8 clkbuf_5_9__f_clk (.A(clknet_4_4_0_clk),
    .X(clknet_5_9__leaf_clk));
 sg13g2_buf_8 clkbuf_5_10__f_clk (.A(clknet_4_5_0_clk),
    .X(clknet_5_10__leaf_clk));
 sg13g2_buf_8 clkbuf_5_11__f_clk (.A(clknet_4_5_0_clk),
    .X(clknet_5_11__leaf_clk));
 sg13g2_buf_8 clkbuf_5_12__f_clk (.A(clknet_4_6_0_clk),
    .X(clknet_5_12__leaf_clk));
 sg13g2_buf_8 clkbuf_5_13__f_clk (.A(clknet_4_6_0_clk),
    .X(clknet_5_13__leaf_clk));
 sg13g2_buf_8 clkbuf_5_14__f_clk (.A(clknet_4_7_0_clk),
    .X(clknet_5_14__leaf_clk));
 sg13g2_buf_8 clkbuf_5_15__f_clk (.A(clknet_4_7_0_clk),
    .X(clknet_5_15__leaf_clk));
 sg13g2_buf_8 clkbuf_5_16__f_clk (.A(clknet_4_8_0_clk),
    .X(clknet_5_16__leaf_clk));
 sg13g2_buf_8 clkbuf_5_17__f_clk (.A(clknet_4_8_0_clk),
    .X(clknet_5_17__leaf_clk));
 sg13g2_buf_8 clkbuf_5_18__f_clk (.A(clknet_4_9_0_clk),
    .X(clknet_5_18__leaf_clk));
 sg13g2_buf_8 clkbuf_5_19__f_clk (.A(clknet_4_9_0_clk),
    .X(clknet_5_19__leaf_clk));
 sg13g2_buf_8 clkbuf_5_20__f_clk (.A(clknet_4_10_0_clk),
    .X(clknet_5_20__leaf_clk));
 sg13g2_buf_8 clkbuf_5_21__f_clk (.A(clknet_4_10_0_clk),
    .X(clknet_5_21__leaf_clk));
 sg13g2_buf_8 clkbuf_5_22__f_clk (.A(clknet_4_11_0_clk),
    .X(clknet_5_22__leaf_clk));
 sg13g2_buf_8 clkbuf_5_23__f_clk (.A(clknet_4_11_0_clk),
    .X(clknet_5_23__leaf_clk));
 sg13g2_buf_8 clkbuf_5_24__f_clk (.A(clknet_4_12_0_clk),
    .X(clknet_5_24__leaf_clk));
 sg13g2_buf_8 clkbuf_5_25__f_clk (.A(clknet_4_12_0_clk),
    .X(clknet_5_25__leaf_clk));
 sg13g2_buf_8 clkbuf_5_26__f_clk (.A(clknet_4_13_0_clk),
    .X(clknet_5_26__leaf_clk));
 sg13g2_buf_8 clkbuf_5_27__f_clk (.A(clknet_4_13_0_clk),
    .X(clknet_5_27__leaf_clk));
 sg13g2_buf_8 clkbuf_5_28__f_clk (.A(clknet_4_14_0_clk),
    .X(clknet_5_28__leaf_clk));
 sg13g2_buf_8 clkbuf_5_29__f_clk (.A(clknet_4_14_0_clk),
    .X(clknet_5_29__leaf_clk));
 sg13g2_buf_8 clkbuf_5_30__f_clk (.A(clknet_4_15_0_clk),
    .X(clknet_5_30__leaf_clk));
 sg13g2_buf_8 clkbuf_5_31__f_clk (.A(clknet_4_15_0_clk),
    .X(clknet_5_31__leaf_clk));
 sg13g2_inv_1 clkload0 (.A(clknet_5_1__leaf_clk));
 sg13g2_inv_1 clkload1 (.A(clknet_5_3__leaf_clk));
 sg13g2_inv_1 clkload2 (.A(clknet_5_5__leaf_clk));
 sg13g2_inv_1 clkload3 (.A(clknet_5_7__leaf_clk));
 sg13g2_inv_1 clkload4 (.A(clknet_5_9__leaf_clk));
 sg13g2_inv_1 clkload5 (.A(clknet_5_11__leaf_clk));
 sg13g2_inv_1 clkload6 (.A(clknet_5_13__leaf_clk));
 sg13g2_inv_1 clkload7 (.A(clknet_5_15__leaf_clk));
 sg13g2_inv_1 clkload8 (.A(clknet_5_17__leaf_clk));
 sg13g2_inv_1 clkload9 (.A(clknet_5_19__leaf_clk));
 sg13g2_inv_1 clkload10 (.A(clknet_5_21__leaf_clk));
 sg13g2_inv_1 clkload11 (.A(clknet_5_23__leaf_clk));
 sg13g2_inv_1 clkload12 (.A(clknet_5_25__leaf_clk));
 sg13g2_inv_1 clkload13 (.A(clknet_5_27__leaf_clk));
 sg13g2_inv_1 clkload14 (.A(clknet_5_29__leaf_clk));
 sg13g2_inv_1 clkload15 (.A(clknet_5_31__leaf_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(\cpu0.ir[0] ),
    .X(net270));
 sg13g2_dlygate4sd3_1 hold2 (.A(\cpu0.ir[2] ),
    .X(net271));
 sg13g2_dlygate4sd3_1 hold3 (.A(\cpu0.b_reg[4] ),
    .X(net272));
 sg13g2_dlygate4sd3_1 hold4 (.A(_0088_),
    .X(net273));
 sg13g2_dlygate4sd3_1 hold5 (.A(\cpu0.ir[1] ),
    .X(net274));
 sg13g2_dlygate4sd3_1 hold6 (.A(\cpu0.ram[3][3] ),
    .X(net275));
 sg13g2_dlygate4sd3_1 hold7 (.A(\cpu0.ir[3] ),
    .X(net276));
 sg13g2_dlygate4sd3_1 hold8 (.A(\cpu0.ram[15][6] ),
    .X(net277));
 sg13g2_dlygate4sd3_1 hold9 (.A(\cpu0.b_reg[7] ),
    .X(net278));
 sg13g2_dlygate4sd3_1 hold10 (.A(_0091_),
    .X(net279));
 sg13g2_dlygate4sd3_1 hold11 (.A(\cpu0.ram[7][3] ),
    .X(net280));
 sg13g2_dlygate4sd3_1 hold12 (.A(\cpu0.ram[14][0] ),
    .X(net281));
 sg13g2_dlygate4sd3_1 hold13 (.A(\cpu0.ram[11][6] ),
    .X(net282));
 sg13g2_dlygate4sd3_1 hold14 (.A(\cpu0.b_reg[2] ),
    .X(net283));
 sg13g2_dlygate4sd3_1 hold15 (.A(_0086_),
    .X(net284));
 sg13g2_dlygate4sd3_1 hold16 (.A(\cpu0.ram[1][3] ),
    .X(net285));
 sg13g2_dlygate4sd3_1 hold17 (.A(\cpu0.ir[6] ),
    .X(net286));
 sg13g2_dlygate4sd3_1 hold18 (.A(_0106_),
    .X(net287));
 sg13g2_dlygate4sd3_1 hold19 (.A(uo_out[0]),
    .X(net288));
 sg13g2_dlygate4sd3_1 hold20 (.A(_0116_),
    .X(net289));
 sg13g2_dlygate4sd3_1 hold21 (.A(\cpu0.a_reg[7] ),
    .X(net290));
 sg13g2_dlygate4sd3_1 hold22 (.A(_0099_),
    .X(net291));
 sg13g2_dlygate4sd3_1 hold23 (.A(\cpu0.a_reg[0] ),
    .X(net292));
 sg13g2_dlygate4sd3_1 hold24 (.A(uo_out[1]),
    .X(net293));
 sg13g2_dlygate4sd3_1 hold25 (.A(_0117_),
    .X(net294));
 sg13g2_dlygate4sd3_1 hold26 (.A(\cpu0.b_reg[1] ),
    .X(net295));
 sg13g2_dlygate4sd3_1 hold27 (.A(_0085_),
    .X(net296));
 sg13g2_dlygate4sd3_1 hold28 (.A(\cpu0.b_reg[3] ),
    .X(net297));
 sg13g2_dlygate4sd3_1 hold29 (.A(\cpu0.a_reg[4] ),
    .X(net298));
 sg13g2_dlygate4sd3_1 hold30 (.A(_0096_),
    .X(net299));
 sg13g2_dlygate4sd3_1 hold31 (.A(\cpu0.a_reg[2] ),
    .X(net300));
 sg13g2_dlygate4sd3_1 hold32 (.A(\cpu0.a_reg[1] ),
    .X(net301));
 sg13g2_dlygate4sd3_1 hold33 (.A(\cpu0.ram[12][1] ),
    .X(net302));
 sg13g2_dlygate4sd3_1 hold34 (.A(\cpu0.ram[3][6] ),
    .X(net303));
 sg13g2_dlygate4sd3_1 hold35 (.A(\cpu0.b_reg[6] ),
    .X(net304));
 sg13g2_dlygate4sd3_1 hold36 (.A(_0090_),
    .X(net305));
 sg13g2_dlygate4sd3_1 hold37 (.A(uo_out[5]),
    .X(net306));
 sg13g2_dlygate4sd3_1 hold38 (.A(_0121_),
    .X(net307));
 sg13g2_dlygate4sd3_1 hold39 (.A(\cpu0.ram[0][1] ),
    .X(net308));
 sg13g2_dlygate4sd3_1 hold40 (.A(uo_out[6]),
    .X(net309));
 sg13g2_dlygate4sd3_1 hold41 (.A(_0122_),
    .X(net310));
 sg13g2_dlygate4sd3_1 hold42 (.A(\cpu0.ram[13][5] ),
    .X(net311));
 sg13g2_dlygate4sd3_1 hold43 (.A(\cpu0.ram[2][0] ),
    .X(net312));
 sg13g2_dlygate4sd3_1 hold44 (.A(uo_out[2]),
    .X(net313));
 sg13g2_dlygate4sd3_1 hold45 (.A(_0118_),
    .X(net314));
 sg13g2_dlygate4sd3_1 hold46 (.A(\cpu0.ram[0][4] ),
    .X(net315));
 sg13g2_dlygate4sd3_1 hold47 (.A(\cpu0.ram[12][0] ),
    .X(net316));
 sg13g2_dlygate4sd3_1 hold48 (.A(\cpu0.ram[7][6] ),
    .X(net317));
 sg13g2_dlygate4sd3_1 hold49 (.A(\cpu0.ram[7][7] ),
    .X(net318));
 sg13g2_dlygate4sd3_1 hold50 (.A(\cpu0.ram[6][1] ),
    .X(net319));
 sg13g2_dlygate4sd3_1 hold51 (.A(\cpu0.ram[5][7] ),
    .X(net320));
 sg13g2_dlygate4sd3_1 hold52 (.A(\cpu0.ram[11][2] ),
    .X(net321));
 sg13g2_dlygate4sd3_1 hold53 (.A(\cpu0.ram[15][4] ),
    .X(net322));
 sg13g2_dlygate4sd3_1 hold54 (.A(\cpu0.ram[10][0] ),
    .X(net323));
 sg13g2_dlygate4sd3_1 hold55 (.A(\cpu0.ram[5][6] ),
    .X(net324));
 sg13g2_dlygate4sd3_1 hold56 (.A(\cpu0.ram[2][1] ),
    .X(net325));
 sg13g2_dlygate4sd3_1 hold57 (.A(\cpu0.ram[8][7] ),
    .X(net326));
 sg13g2_dlygate4sd3_1 hold58 (.A(\cpu0.ram[4][3] ),
    .X(net327));
 sg13g2_dlygate4sd3_1 hold59 (.A(\cpu0.ram[11][4] ),
    .X(net328));
 sg13g2_dlygate4sd3_1 hold60 (.A(\cpu0.ram[4][5] ),
    .X(net329));
 sg13g2_dlygate4sd3_1 hold61 (.A(\cpu0.ram[9][5] ),
    .X(net330));
 sg13g2_dlygate4sd3_1 hold62 (.A(\cpu0.ram[3][4] ),
    .X(net331));
 sg13g2_dlygate4sd3_1 hold63 (.A(\cpu0.ram[13][1] ),
    .X(net332));
 sg13g2_dlygate4sd3_1 hold64 (.A(\cpu0.a_reg[6] ),
    .X(net333));
 sg13g2_dlygate4sd3_1 hold65 (.A(_0098_),
    .X(net334));
 sg13g2_dlygate4sd3_1 hold66 (.A(\cpu0.ram[14][5] ),
    .X(net335));
 sg13g2_dlygate4sd3_1 hold67 (.A(\cpu0.ram[15][0] ),
    .X(net336));
 sg13g2_dlygate4sd3_1 hold68 (.A(\cpu0.ram[5][4] ),
    .X(net337));
 sg13g2_dlygate4sd3_1 hold69 (.A(\cpu0.ram[9][0] ),
    .X(net338));
 sg13g2_dlygate4sd3_1 hold70 (.A(\cpu0.ram[9][3] ),
    .X(net339));
 sg13g2_dlygate4sd3_1 hold71 (.A(\cpu0.ram[11][5] ),
    .X(net340));
 sg13g2_dlygate4sd3_1 hold72 (.A(\cpu0.ram[13][7] ),
    .X(net341));
 sg13g2_dlygate4sd3_1 hold73 (.A(\cpu0.ram[15][1] ),
    .X(net342));
 sg13g2_dlygate4sd3_1 hold74 (.A(\cpu0.ram[2][2] ),
    .X(net343));
 sg13g2_dlygate4sd3_1 hold75 (.A(\cpu0.ram[2][3] ),
    .X(net344));
 sg13g2_dlygate4sd3_1 hold76 (.A(\cpu0.ram[15][3] ),
    .X(net345));
 sg13g2_dlygate4sd3_1 hold77 (.A(\cpu0.ram[9][2] ),
    .X(net346));
 sg13g2_dlygate4sd3_1 hold78 (.A(\cpu0.b_reg[0] ),
    .X(net347));
 sg13g2_dlygate4sd3_1 hold79 (.A(_0084_),
    .X(net348));
 sg13g2_dlygate4sd3_1 hold80 (.A(\cpu0.ram[13][4] ),
    .X(net349));
 sg13g2_dlygate4sd3_1 hold81 (.A(\cpu0.ram[8][6] ),
    .X(net350));
 sg13g2_dlygate4sd3_1 hold82 (.A(\cpu0.ram[13][3] ),
    .X(net351));
 sg13g2_dlygate4sd3_1 hold83 (.A(\cpu0.ram[5][2] ),
    .X(net352));
 sg13g2_dlygate4sd3_1 hold84 (.A(\cpu0.ram[12][6] ),
    .X(net353));
 sg13g2_dlygate4sd3_1 hold85 (.A(\cpu0.ram[9][6] ),
    .X(net354));
 sg13g2_dlygate4sd3_1 hold86 (.A(\cpu0.ram[1][2] ),
    .X(net355));
 sg13g2_dlygate4sd3_1 hold87 (.A(\cpu0.ram[4][4] ),
    .X(net356));
 sg13g2_dlygate4sd3_1 hold88 (.A(\cpu0.ram[3][5] ),
    .X(net357));
 sg13g2_dlygate4sd3_1 hold89 (.A(\cpu0.ram[15][5] ),
    .X(net358));
 sg13g2_dlygate4sd3_1 hold90 (.A(\cpu0.ram[3][1] ),
    .X(net359));
 sg13g2_dlygate4sd3_1 hold91 (.A(\cpu0.ram[6][0] ),
    .X(net360));
 sg13g2_dlygate4sd3_1 hold92 (.A(\cpu0.ram[6][4] ),
    .X(net361));
 sg13g2_dlygate4sd3_1 hold93 (.A(\cpu0.ram[5][3] ),
    .X(net362));
 sg13g2_dlygate4sd3_1 hold94 (.A(\cpu0.ram[3][7] ),
    .X(net363));
 sg13g2_dlygate4sd3_1 hold95 (.A(\cpu0.ram[5][0] ),
    .X(net364));
 sg13g2_dlygate4sd3_1 hold96 (.A(\cpu0.ram[15][7] ),
    .X(net365));
 sg13g2_dlygate4sd3_1 hold97 (.A(\cpu0.ram[11][7] ),
    .X(net366));
 sg13g2_dlygate4sd3_1 hold98 (.A(\cpu0.ram[14][2] ),
    .X(net367));
 sg13g2_dlygate4sd3_1 hold99 (.A(\cpu0.ram[4][0] ),
    .X(net368));
 sg13g2_dlygate4sd3_1 hold100 (.A(\cpu0.ram[12][2] ),
    .X(net369));
 sg13g2_dlygate4sd3_1 hold101 (.A(\cpu0.ram[11][0] ),
    .X(net370));
 sg13g2_dlygate4sd3_1 hold102 (.A(\cpu0.ram[2][6] ),
    .X(net371));
 sg13g2_dlygate4sd3_1 hold103 (.A(\cpu0.b_reg[5] ),
    .X(net372));
 sg13g2_dlygate4sd3_1 hold104 (.A(_0089_),
    .X(net373));
 sg13g2_dlygate4sd3_1 hold105 (.A(\cpu0.ram[4][1] ),
    .X(net374));
 sg13g2_dlygate4sd3_1 hold106 (.A(\cpu0.ram[6][2] ),
    .X(net375));
 sg13g2_dlygate4sd3_1 hold107 (.A(\cpu0.ram[14][7] ),
    .X(net376));
 sg13g2_dlygate4sd3_1 hold108 (.A(\cpu0.ram[14][1] ),
    .X(net377));
 sg13g2_dlygate4sd3_1 hold109 (.A(\cpu0.ram[1][6] ),
    .X(net378));
 sg13g2_dlygate4sd3_1 hold110 (.A(\cpu0.ram[13][6] ),
    .X(net379));
 sg13g2_dlygate4sd3_1 hold111 (.A(\cpu0.ram[4][7] ),
    .X(net380));
 sg13g2_dlygate4sd3_1 hold112 (.A(\cpu0.ram[0][3] ),
    .X(net381));
 sg13g2_dlygate4sd3_1 hold113 (.A(\cpu0.ram[6][7] ),
    .X(net382));
 sg13g2_dlygate4sd3_1 hold114 (.A(\cpu0.ram[5][1] ),
    .X(net383));
 sg13g2_dlygate4sd3_1 hold115 (.A(\cpu0.ram[1][1] ),
    .X(net384));
 sg13g2_dlygate4sd3_1 hold116 (.A(\cpu0.ram[0][2] ),
    .X(net385));
 sg13g2_dlygate4sd3_1 hold117 (.A(\cpu0.ram[4][2] ),
    .X(net386));
 sg13g2_dlygate4sd3_1 hold118 (.A(\cpu0.ram[11][3] ),
    .X(net387));
 sg13g2_dlygate4sd3_1 hold119 (.A(\cpu0.ram[6][5] ),
    .X(net388));
 sg13g2_dlygate4sd3_1 hold120 (.A(\cpu0.ram[8][1] ),
    .X(net389));
 sg13g2_dlygate4sd3_1 hold121 (.A(\cpu0.ram[0][0] ),
    .X(net390));
 sg13g2_dlygate4sd3_1 hold122 (.A(\cpu0.ram[14][6] ),
    .X(net391));
 sg13g2_dlygate4sd3_1 hold123 (.A(\cpu0.ram[2][5] ),
    .X(net392));
 sg13g2_dlygate4sd3_1 hold124 (.A(\cpu0.ram[12][5] ),
    .X(net393));
 sg13g2_dlygate4sd3_1 hold125 (.A(\cpu0.ram[0][6] ),
    .X(net394));
 sg13g2_dlygate4sd3_1 hold126 (.A(\cpu0.ram[8][2] ),
    .X(net395));
 sg13g2_dlygate4sd3_1 hold127 (.A(\cpu0.ram[12][3] ),
    .X(net396));
 sg13g2_dlygate4sd3_1 hold128 (.A(\cpu0.ram[8][0] ),
    .X(net397));
 sg13g2_dlygate4sd3_1 hold129 (.A(\cpu0.ram[13][2] ),
    .X(net398));
 sg13g2_dlygate4sd3_1 hold130 (.A(uo_out[3]),
    .X(net399));
 sg13g2_dlygate4sd3_1 hold131 (.A(_0119_),
    .X(net400));
 sg13g2_dlygate4sd3_1 hold132 (.A(\cpu0.ram[1][7] ),
    .X(net401));
 sg13g2_dlygate4sd3_1 hold133 (.A(\cpu0.ram[8][3] ),
    .X(net402));
 sg13g2_dlygate4sd3_1 hold134 (.A(\cpu0.ram[11][1] ),
    .X(net403));
 sg13g2_dlygate4sd3_1 hold135 (.A(\cpu0.a_reg[5] ),
    .X(net404));
 sg13g2_dlygate4sd3_1 hold136 (.A(_0097_),
    .X(net405));
 sg13g2_dlygate4sd3_1 hold137 (.A(\cpu0.ram[6][6] ),
    .X(net406));
 sg13g2_dlygate4sd3_1 hold138 (.A(\cpu0.ram[7][2] ),
    .X(net407));
 sg13g2_dlygate4sd3_1 hold139 (.A(uo_out[7]),
    .X(net408));
 sg13g2_dlygate4sd3_1 hold140 (.A(_0123_),
    .X(net409));
 sg13g2_dlygate4sd3_1 hold141 (.A(\cpu0.ram[1][0] ),
    .X(net410));
 sg13g2_dlygate4sd3_1 hold142 (.A(\cpu0.ram[3][2] ),
    .X(net411));
 sg13g2_dlygate4sd3_1 hold143 (.A(\cpu0.ram[13][0] ),
    .X(net412));
 sg13g2_dlygate4sd3_1 hold144 (.A(\cpu0.ir[5] ),
    .X(net413));
 sg13g2_dlygate4sd3_1 hold145 (.A(_0105_),
    .X(net414));
 sg13g2_dlygate4sd3_1 hold146 (.A(\cpu0.ram[10][6] ),
    .X(net415));
 sg13g2_dlygate4sd3_1 hold147 (.A(\cpu0.ram[9][1] ),
    .X(net416));
 sg13g2_dlygate4sd3_1 hold148 (.A(\cpu0.ram[9][7] ),
    .X(net417));
 sg13g2_dlygate4sd3_1 hold149 (.A(\cpu0.ram[8][4] ),
    .X(net418));
 sg13g2_dlygate4sd3_1 hold150 (.A(\cpu0.ram[10][5] ),
    .X(net419));
 sg13g2_dlygate4sd3_1 hold151 (.A(\cpu0.ram[7][5] ),
    .X(net420));
 sg13g2_dlygate4sd3_1 hold152 (.A(\cpu0.ram[0][5] ),
    .X(net421));
 sg13g2_dlygate4sd3_1 hold153 (.A(\cpu0.ram[14][4] ),
    .X(net422));
 sg13g2_dlygate4sd3_1 hold154 (.A(\cpu0.ram[4][6] ),
    .X(net423));
 sg13g2_dlygate4sd3_1 hold155 (.A(\cpu0.ram[10][7] ),
    .X(net424));
 sg13g2_dlygate4sd3_1 hold156 (.A(\cpu0.ram[12][4] ),
    .X(net425));
 sg13g2_dlygate4sd3_1 hold157 (.A(\cpu0.ram[3][0] ),
    .X(net426));
 sg13g2_dlygate4sd3_1 hold158 (.A(\cpu0.ram[10][3] ),
    .X(net427));
 sg13g2_dlygate4sd3_1 hold159 (.A(\cpu0.ram[0][7] ),
    .X(net428));
 sg13g2_dlygate4sd3_1 hold160 (.A(\cpu0.ram[14][3] ),
    .X(net429));
 sg13g2_dlygate4sd3_1 hold161 (.A(\cpu0.ram[10][1] ),
    .X(net430));
 sg13g2_dlygate4sd3_1 hold162 (.A(\cpu0.ram[1][4] ),
    .X(net431));
 sg13g2_dlygate4sd3_1 hold163 (.A(\cpu0.ram[2][4] ),
    .X(net432));
 sg13g2_dlygate4sd3_1 hold164 (.A(\cpu0.ram[7][1] ),
    .X(net433));
 sg13g2_dlygate4sd3_1 hold165 (.A(\cpu0.ram[7][0] ),
    .X(net434));
 sg13g2_dlygate4sd3_1 hold166 (.A(\cpu0.ram[6][3] ),
    .X(net435));
 sg13g2_dlygate4sd3_1 hold167 (.A(uo_out[4]),
    .X(net436));
 sg13g2_dlygate4sd3_1 hold168 (.A(_0120_),
    .X(net437));
 sg13g2_dlygate4sd3_1 hold169 (.A(\cpu0.ram[10][2] ),
    .X(net438));
 sg13g2_dlygate4sd3_1 hold170 (.A(\cpu0.ram[9][4] ),
    .X(net439));
 sg13g2_dlygate4sd3_1 hold171 (.A(\cpu0.ram[8][5] ),
    .X(net440));
 sg13g2_dlygate4sd3_1 hold172 (.A(\cpu0.ram[1][5] ),
    .X(net441));
 sg13g2_dlygate4sd3_1 hold173 (.A(\cpu0.ram[15][2] ),
    .X(net442));
 sg13g2_dlygate4sd3_1 hold174 (.A(\cpu0.ram[2][7] ),
    .X(net443));
 sg13g2_dlygate4sd3_1 hold175 (.A(\cpu0.ram[5][5] ),
    .X(net444));
 sg13g2_dlygate4sd3_1 hold176 (.A(\cpu0.ram[12][7] ),
    .X(net445));
 sg13g2_dlygate4sd3_1 hold177 (.A(\cpu0.ir[7] ),
    .X(net446));
 sg13g2_dlygate4sd3_1 hold178 (.A(\cpu0.ram[7][4] ),
    .X(net447));
 sg13g2_dlygate4sd3_1 hold179 (.A(\cpu0.ram[10][4] ),
    .X(net448));
 sg13g2_dlygate4sd3_1 hold180 (.A(\cpu0.ir[4] ),
    .X(net449));
 sg13g2_dlygate4sd3_1 hold181 (.A(\cpu0.a_reg[3] ),
    .X(net450));
 sg13g2_dlygate4sd3_1 hold182 (.A(\cpu0.zero_flag ),
    .X(net451));
 sg13g2_dlygate4sd3_1 hold183 (.A(\cpu0.mar[3] ),
    .X(net452));
 sg13g2_dlygate4sd3_1 hold184 (.A(_0015_),
    .X(net453));
 sg13g2_dlygate4sd3_1 hold185 (.A(\cpu0.mar[2] ),
    .X(net454));
 sg13g2_dlygate4sd3_1 hold186 (.A(_0014_),
    .X(net455));
 sg13g2_dlygate4sd3_1 hold187 (.A(\cpu0.step[1] ),
    .X(net456));
 sg13g2_dlygate4sd3_1 hold188 (.A(\cpu0.mar[0] ),
    .X(net457));
 sg13g2_dlygate4sd3_1 hold189 (.A(\cpu0.pc[3] ),
    .X(net458));
 sg13g2_dlygate4sd3_1 hold190 (.A(\cpu0.step[2] ),
    .X(net459));
 sg13g2_dlygate4sd3_1 hold191 (.A(_0033_),
    .X(net460));
 sg13g2_dlygate4sd3_1 hold192 (.A(\cpu0.pc[0] ),
    .X(net461));
 sg13g2_dlygate4sd3_1 hold193 (.A(\cpu0.mar[1] ),
    .X(net462));
 sg13g2_dlygate4sd3_1 hold194 (.A(\cpu0.pc[1] ),
    .X(net463));
 sg13g2_dlygate4sd3_1 hold195 (.A(\cpu0.step[0] ),
    .X(net464));
 sg13g2_dlygate4sd3_1 hold196 (.A(\cpu0.pc[2] ),
    .X(net465));
 sg13g2_dlygate4sd3_1 hold197 (.A(\cpu0.step[0] ),
    .X(net466));
 sg13g2_dlygate4sd3_1 hold198 (.A(\cpu0.step[2] ),
    .X(net467));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_4 FILLER_0_112 ();
 sg13g2_fill_1 FILLER_0_116 ();
 sg13g2_decap_8 FILLER_0_144 ();
 sg13g2_decap_8 FILLER_0_151 ();
 sg13g2_decap_4 FILLER_0_158 ();
 sg13g2_fill_1 FILLER_0_162 ();
 sg13g2_decap_8 FILLER_0_199 ();
 sg13g2_decap_8 FILLER_0_206 ();
 sg13g2_decap_4 FILLER_0_213 ();
 sg13g2_fill_2 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_246 ();
 sg13g2_decap_8 FILLER_0_253 ();
 sg13g2_fill_2 FILLER_0_260 ();
 sg13g2_decap_8 FILLER_0_270 ();
 sg13g2_decap_8 FILLER_0_277 ();
 sg13g2_decap_8 FILLER_0_284 ();
 sg13g2_decap_8 FILLER_0_291 ();
 sg13g2_decap_4 FILLER_0_298 ();
 sg13g2_fill_2 FILLER_0_302 ();
 sg13g2_decap_8 FILLER_0_331 ();
 sg13g2_decap_8 FILLER_0_338 ();
 sg13g2_fill_2 FILLER_0_345 ();
 sg13g2_decap_8 FILLER_0_374 ();
 sg13g2_decap_8 FILLER_0_381 ();
 sg13g2_decap_8 FILLER_0_388 ();
 sg13g2_decap_8 FILLER_0_395 ();
 sg13g2_decap_8 FILLER_0_402 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_fill_1 FILLER_1_105 ();
 sg13g2_fill_2 FILLER_1_115 ();
 sg13g2_decap_8 FILLER_1_153 ();
 sg13g2_decap_4 FILLER_1_160 ();
 sg13g2_fill_1 FILLER_1_164 ();
 sg13g2_decap_8 FILLER_1_201 ();
 sg13g2_decap_8 FILLER_1_208 ();
 sg13g2_fill_1 FILLER_1_215 ();
 sg13g2_decap_8 FILLER_1_243 ();
 sg13g2_decap_8 FILLER_1_250 ();
 sg13g2_fill_1 FILLER_1_257 ();
 sg13g2_decap_8 FILLER_1_285 ();
 sg13g2_fill_1 FILLER_1_292 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_4 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_374 ();
 sg13g2_decap_8 FILLER_1_381 ();
 sg13g2_decap_8 FILLER_1_388 ();
 sg13g2_decap_8 FILLER_1_395 ();
 sg13g2_decap_8 FILLER_1_402 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_4 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_43 ();
 sg13g2_decap_8 FILLER_2_50 ();
 sg13g2_decap_8 FILLER_2_57 ();
 sg13g2_decap_8 FILLER_2_64 ();
 sg13g2_decap_8 FILLER_2_71 ();
 sg13g2_decap_8 FILLER_2_78 ();
 sg13g2_decap_8 FILLER_2_85 ();
 sg13g2_fill_1 FILLER_2_92 ();
 sg13g2_fill_2 FILLER_2_103 ();
 sg13g2_fill_1 FILLER_2_105 ();
 sg13g2_fill_2 FILLER_2_116 ();
 sg13g2_fill_1 FILLER_2_212 ();
 sg13g2_fill_1 FILLER_2_284 ();
 sg13g2_fill_2 FILLER_2_359 ();
 sg13g2_fill_2 FILLER_2_370 ();
 sg13g2_decap_8 FILLER_2_381 ();
 sg13g2_decap_8 FILLER_2_388 ();
 sg13g2_decap_8 FILLER_2_395 ();
 sg13g2_decap_8 FILLER_2_402 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_fill_2 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_43 ();
 sg13g2_decap_8 FILLER_3_50 ();
 sg13g2_decap_8 FILLER_3_57 ();
 sg13g2_decap_8 FILLER_3_64 ();
 sg13g2_decap_8 FILLER_3_71 ();
 sg13g2_decap_8 FILLER_3_78 ();
 sg13g2_fill_2 FILLER_3_85 ();
 sg13g2_fill_2 FILLER_3_140 ();
 sg13g2_fill_2 FILLER_3_169 ();
 sg13g2_fill_1 FILLER_3_171 ();
 sg13g2_fill_2 FILLER_3_196 ();
 sg13g2_fill_1 FILLER_3_198 ();
 sg13g2_decap_8 FILLER_3_208 ();
 sg13g2_decap_4 FILLER_3_215 ();
 sg13g2_decap_4 FILLER_3_246 ();
 sg13g2_fill_2 FILLER_3_293 ();
 sg13g2_fill_2 FILLER_3_322 ();
 sg13g2_fill_1 FILLER_3_324 ();
 sg13g2_fill_1 FILLER_3_338 ();
 sg13g2_fill_2 FILLER_3_354 ();
 sg13g2_fill_1 FILLER_3_356 ();
 sg13g2_fill_1 FILLER_3_376 ();
 sg13g2_decap_4 FILLER_3_404 ();
 sg13g2_fill_1 FILLER_3_408 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_fill_2 FILLER_4_7 ();
 sg13g2_fill_1 FILLER_4_9 ();
 sg13g2_decap_8 FILLER_4_55 ();
 sg13g2_decap_8 FILLER_4_62 ();
 sg13g2_decap_4 FILLER_4_69 ();
 sg13g2_fill_2 FILLER_4_131 ();
 sg13g2_fill_1 FILLER_4_133 ();
 sg13g2_decap_4 FILLER_4_181 ();
 sg13g2_fill_2 FILLER_4_206 ();
 sg13g2_fill_1 FILLER_4_226 ();
 sg13g2_fill_1 FILLER_4_346 ();
 sg13g2_decap_8 FILLER_4_402 ();
 sg13g2_decap_4 FILLER_5_0 ();
 sg13g2_fill_1 FILLER_5_4 ();
 sg13g2_fill_2 FILLER_5_72 ();
 sg13g2_decap_8 FILLER_5_123 ();
 sg13g2_decap_8 FILLER_5_130 ();
 sg13g2_decap_4 FILLER_5_137 ();
 sg13g2_decap_8 FILLER_5_175 ();
 sg13g2_fill_1 FILLER_5_182 ();
 sg13g2_decap_8 FILLER_5_196 ();
 sg13g2_decap_4 FILLER_5_203 ();
 sg13g2_fill_2 FILLER_5_207 ();
 sg13g2_decap_4 FILLER_5_236 ();
 sg13g2_decap_8 FILLER_5_276 ();
 sg13g2_fill_2 FILLER_5_303 ();
 sg13g2_fill_1 FILLER_5_356 ();
 sg13g2_fill_2 FILLER_5_362 ();
 sg13g2_decap_4 FILLER_5_404 ();
 sg13g2_fill_1 FILLER_5_408 ();
 sg13g2_fill_1 FILLER_6_39 ();
 sg13g2_decap_4 FILLER_6_61 ();
 sg13g2_decap_8 FILLER_6_68 ();
 sg13g2_decap_8 FILLER_6_75 ();
 sg13g2_fill_2 FILLER_6_82 ();
 sg13g2_fill_1 FILLER_6_84 ();
 sg13g2_fill_2 FILLER_6_104 ();
 sg13g2_fill_1 FILLER_6_106 ();
 sg13g2_decap_8 FILLER_6_128 ();
 sg13g2_fill_2 FILLER_6_135 ();
 sg13g2_fill_1 FILLER_6_137 ();
 sg13g2_fill_2 FILLER_6_151 ();
 sg13g2_decap_8 FILLER_6_171 ();
 sg13g2_fill_1 FILLER_6_178 ();
 sg13g2_decap_4 FILLER_6_206 ();
 sg13g2_fill_2 FILLER_6_248 ();
 sg13g2_decap_8 FILLER_6_274 ();
 sg13g2_decap_8 FILLER_6_281 ();
 sg13g2_fill_2 FILLER_6_288 ();
 sg13g2_decap_4 FILLER_6_305 ();
 sg13g2_fill_2 FILLER_6_322 ();
 sg13g2_decap_4 FILLER_6_338 ();
 sg13g2_fill_1 FILLER_6_356 ();
 sg13g2_fill_1 FILLER_6_382 ();
 sg13g2_decap_8 FILLER_6_387 ();
 sg13g2_decap_8 FILLER_6_394 ();
 sg13g2_decap_8 FILLER_6_401 ();
 sg13g2_fill_1 FILLER_6_408 ();
 sg13g2_decap_4 FILLER_7_0 ();
 sg13g2_fill_2 FILLER_7_4 ();
 sg13g2_fill_1 FILLER_7_52 ();
 sg13g2_fill_2 FILLER_7_66 ();
 sg13g2_decap_8 FILLER_7_81 ();
 sg13g2_fill_2 FILLER_7_88 ();
 sg13g2_decap_8 FILLER_7_94 ();
 sg13g2_fill_2 FILLER_7_105 ();
 sg13g2_fill_1 FILLER_7_116 ();
 sg13g2_decap_4 FILLER_7_130 ();
 sg13g2_fill_1 FILLER_7_134 ();
 sg13g2_fill_1 FILLER_7_172 ();
 sg13g2_decap_4 FILLER_7_210 ();
 sg13g2_decap_4 FILLER_7_224 ();
 sg13g2_fill_1 FILLER_7_228 ();
 sg13g2_decap_8 FILLER_7_234 ();
 sg13g2_decap_8 FILLER_7_241 ();
 sg13g2_fill_2 FILLER_7_248 ();
 sg13g2_decap_8 FILLER_7_258 ();
 sg13g2_fill_1 FILLER_7_265 ();
 sg13g2_decap_8 FILLER_7_279 ();
 sg13g2_decap_8 FILLER_7_330 ();
 sg13g2_fill_2 FILLER_7_337 ();
 sg13g2_fill_1 FILLER_7_339 ();
 sg13g2_decap_4 FILLER_7_381 ();
 sg13g2_fill_2 FILLER_7_385 ();
 sg13g2_fill_2 FILLER_7_396 ();
 sg13g2_fill_1 FILLER_7_398 ();
 sg13g2_decap_8 FILLER_7_402 ();
 sg13g2_fill_2 FILLER_8_0 ();
 sg13g2_fill_1 FILLER_8_2 ();
 sg13g2_decap_8 FILLER_8_43 ();
 sg13g2_fill_1 FILLER_8_50 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_fill_1 FILLER_8_104 ();
 sg13g2_fill_2 FILLER_8_129 ();
 sg13g2_fill_1 FILLER_8_131 ();
 sg13g2_fill_2 FILLER_8_145 ();
 sg13g2_fill_1 FILLER_8_147 ();
 sg13g2_fill_2 FILLER_8_193 ();
 sg13g2_fill_2 FILLER_8_204 ();
 sg13g2_decap_8 FILLER_8_209 ();
 sg13g2_fill_1 FILLER_8_216 ();
 sg13g2_decap_8 FILLER_8_225 ();
 sg13g2_fill_1 FILLER_8_242 ();
 sg13g2_decap_8 FILLER_8_275 ();
 sg13g2_decap_8 FILLER_8_282 ();
 sg13g2_decap_4 FILLER_8_289 ();
 sg13g2_fill_1 FILLER_8_293 ();
 sg13g2_fill_2 FILLER_8_330 ();
 sg13g2_fill_2 FILLER_8_407 ();
 sg13g2_decap_4 FILLER_9_0 ();
 sg13g2_decap_4 FILLER_9_45 ();
 sg13g2_decap_8 FILLER_9_130 ();
 sg13g2_fill_1 FILLER_9_137 ();
 sg13g2_fill_1 FILLER_9_183 ();
 sg13g2_decap_4 FILLER_9_188 ();
 sg13g2_fill_1 FILLER_9_192 ();
 sg13g2_fill_2 FILLER_9_229 ();
 sg13g2_fill_1 FILLER_9_231 ();
 sg13g2_decap_4 FILLER_9_281 ();
 sg13g2_fill_2 FILLER_9_336 ();
 sg13g2_fill_2 FILLER_9_361 ();
 sg13g2_fill_1 FILLER_9_399 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_4 FILLER_10_62 ();
 sg13g2_fill_2 FILLER_10_66 ();
 sg13g2_fill_2 FILLER_10_96 ();
 sg13g2_fill_2 FILLER_10_164 ();
 sg13g2_decap_8 FILLER_10_190 ();
 sg13g2_decap_8 FILLER_10_197 ();
 sg13g2_fill_1 FILLER_10_204 ();
 sg13g2_decap_4 FILLER_10_236 ();
 sg13g2_fill_2 FILLER_10_250 ();
 sg13g2_fill_1 FILLER_10_288 ();
 sg13g2_fill_1 FILLER_10_309 ();
 sg13g2_fill_1 FILLER_10_341 ();
 sg13g2_fill_2 FILLER_10_374 ();
 sg13g2_fill_1 FILLER_10_376 ();
 sg13g2_fill_2 FILLER_10_407 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_fill_2 FILLER_11_7 ();
 sg13g2_fill_1 FILLER_11_9 ();
 sg13g2_decap_8 FILLER_11_43 ();
 sg13g2_decap_8 FILLER_11_63 ();
 sg13g2_decap_8 FILLER_11_70 ();
 sg13g2_fill_1 FILLER_11_77 ();
 sg13g2_fill_1 FILLER_11_96 ();
 sg13g2_fill_2 FILLER_11_151 ();
 sg13g2_decap_8 FILLER_11_197 ();
 sg13g2_fill_2 FILLER_11_204 ();
 sg13g2_fill_1 FILLER_11_206 ();
 sg13g2_fill_2 FILLER_11_248 ();
 sg13g2_fill_1 FILLER_11_265 ();
 sg13g2_fill_1 FILLER_11_306 ();
 sg13g2_fill_1 FILLER_11_325 ();
 sg13g2_fill_1 FILLER_11_377 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_4 FILLER_12_7 ();
 sg13g2_decap_4 FILLER_12_72 ();
 sg13g2_fill_1 FILLER_12_103 ();
 sg13g2_fill_1 FILLER_12_122 ();
 sg13g2_fill_2 FILLER_12_128 ();
 sg13g2_decap_8 FILLER_12_133 ();
 sg13g2_decap_8 FILLER_12_140 ();
 sg13g2_decap_4 FILLER_12_147 ();
 sg13g2_fill_2 FILLER_12_151 ();
 sg13g2_decap_8 FILLER_12_190 ();
 sg13g2_decap_4 FILLER_12_197 ();
 sg13g2_fill_2 FILLER_12_214 ();
 sg13g2_fill_1 FILLER_12_216 ();
 sg13g2_fill_2 FILLER_12_310 ();
 sg13g2_fill_2 FILLER_12_354 ();
 sg13g2_fill_1 FILLER_12_356 ();
 sg13g2_fill_1 FILLER_12_376 ();
 sg13g2_decap_4 FILLER_12_404 ();
 sg13g2_fill_1 FILLER_12_408 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_fill_2 FILLER_13_7 ();
 sg13g2_fill_2 FILLER_13_80 ();
 sg13g2_fill_1 FILLER_13_82 ();
 sg13g2_fill_2 FILLER_13_120 ();
 sg13g2_fill_1 FILLER_13_122 ();
 sg13g2_decap_8 FILLER_13_133 ();
 sg13g2_fill_1 FILLER_13_140 ();
 sg13g2_decap_8 FILLER_13_190 ();
 sg13g2_decap_8 FILLER_13_197 ();
 sg13g2_decap_8 FILLER_13_204 ();
 sg13g2_fill_1 FILLER_13_211 ();
 sg13g2_decap_4 FILLER_13_217 ();
 sg13g2_fill_2 FILLER_13_267 ();
 sg13g2_fill_2 FILLER_13_309 ();
 sg13g2_fill_1 FILLER_13_311 ();
 sg13g2_fill_2 FILLER_13_351 ();
 sg13g2_fill_1 FILLER_13_353 ();
 sg13g2_decap_4 FILLER_13_363 ();
 sg13g2_decap_4 FILLER_13_404 ();
 sg13g2_fill_1 FILLER_13_408 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_fill_2 FILLER_14_7 ();
 sg13g2_decap_4 FILLER_14_54 ();
 sg13g2_fill_2 FILLER_14_67 ();
 sg13g2_fill_1 FILLER_14_69 ();
 sg13g2_fill_2 FILLER_14_120 ();
 sg13g2_fill_1 FILLER_14_122 ();
 sg13g2_fill_2 FILLER_14_150 ();
 sg13g2_fill_1 FILLER_14_152 ();
 sg13g2_decap_8 FILLER_14_185 ();
 sg13g2_decap_8 FILLER_14_192 ();
 sg13g2_decap_8 FILLER_14_199 ();
 sg13g2_fill_2 FILLER_14_206 ();
 sg13g2_fill_1 FILLER_14_208 ();
 sg13g2_fill_2 FILLER_14_218 ();
 sg13g2_fill_1 FILLER_14_220 ();
 sg13g2_fill_2 FILLER_14_234 ();
 sg13g2_fill_1 FILLER_14_236 ();
 sg13g2_fill_2 FILLER_14_312 ();
 sg13g2_fill_1 FILLER_14_314 ();
 sg13g2_fill_1 FILLER_14_342 ();
 sg13g2_decap_8 FILLER_14_400 ();
 sg13g2_fill_2 FILLER_14_407 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_66 ();
 sg13g2_fill_2 FILLER_15_73 ();
 sg13g2_fill_1 FILLER_15_115 ();
 sg13g2_decap_8 FILLER_15_143 ();
 sg13g2_decap_8 FILLER_15_150 ();
 sg13g2_decap_8 FILLER_15_157 ();
 sg13g2_fill_2 FILLER_15_164 ();
 sg13g2_decap_8 FILLER_15_171 ();
 sg13g2_decap_4 FILLER_15_178 ();
 sg13g2_fill_2 FILLER_15_192 ();
 sg13g2_decap_8 FILLER_15_229 ();
 sg13g2_decap_8 FILLER_15_236 ();
 sg13g2_decap_4 FILLER_15_243 ();
 sg13g2_fill_1 FILLER_15_247 ();
 sg13g2_decap_8 FILLER_15_275 ();
 sg13g2_fill_1 FILLER_15_282 ();
 sg13g2_decap_8 FILLER_15_287 ();
 sg13g2_decap_8 FILLER_15_294 ();
 sg13g2_fill_1 FILLER_15_301 ();
 sg13g2_decap_4 FILLER_15_338 ();
 sg13g2_fill_1 FILLER_15_355 ();
 sg13g2_decap_8 FILLER_15_396 ();
 sg13g2_decap_4 FILLER_15_403 ();
 sg13g2_fill_2 FILLER_15_407 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_fill_2 FILLER_16_41 ();
 sg13g2_fill_2 FILLER_16_53 ();
 sg13g2_fill_1 FILLER_16_55 ();
 sg13g2_fill_1 FILLER_16_65 ();
 sg13g2_fill_2 FILLER_16_102 ();
 sg13g2_fill_1 FILLER_16_104 ();
 sg13g2_fill_1 FILLER_16_114 ();
 sg13g2_decap_8 FILLER_16_142 ();
 sg13g2_decap_4 FILLER_16_149 ();
 sg13g2_fill_2 FILLER_16_153 ();
 sg13g2_fill_1 FILLER_16_188 ();
 sg13g2_fill_2 FILLER_16_234 ();
 sg13g2_fill_1 FILLER_16_236 ();
 sg13g2_fill_2 FILLER_16_294 ();
 sg13g2_fill_1 FILLER_16_296 ();
 sg13g2_decap_4 FILLER_16_325 ();
 sg13g2_decap_8 FILLER_16_333 ();
 sg13g2_decap_8 FILLER_16_340 ();
 sg13g2_decap_4 FILLER_16_347 ();
 sg13g2_fill_1 FILLER_16_356 ();
 sg13g2_decap_8 FILLER_16_400 ();
 sg13g2_fill_2 FILLER_16_407 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_4 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_65 ();
 sg13g2_decap_4 FILLER_17_72 ();
 sg13g2_fill_2 FILLER_17_103 ();
 sg13g2_decap_8 FILLER_17_142 ();
 sg13g2_decap_8 FILLER_17_186 ();
 sg13g2_decap_8 FILLER_17_193 ();
 sg13g2_fill_2 FILLER_17_200 ();
 sg13g2_fill_1 FILLER_17_202 ();
 sg13g2_decap_4 FILLER_17_207 ();
 sg13g2_fill_1 FILLER_17_211 ();
 sg13g2_fill_2 FILLER_17_222 ();
 sg13g2_fill_2 FILLER_17_242 ();
 sg13g2_decap_8 FILLER_17_290 ();
 sg13g2_fill_2 FILLER_17_297 ();
 sg13g2_decap_8 FILLER_17_335 ();
 sg13g2_decap_8 FILLER_17_342 ();
 sg13g2_fill_2 FILLER_17_349 ();
 sg13g2_fill_1 FILLER_17_351 ();
 sg13g2_fill_1 FILLER_17_376 ();
 sg13g2_decap_4 FILLER_17_404 ();
 sg13g2_fill_1 FILLER_17_408 ();
 sg13g2_decap_4 FILLER_18_0 ();
 sg13g2_fill_2 FILLER_18_4 ();
 sg13g2_fill_2 FILLER_18_103 ();
 sg13g2_fill_2 FILLER_18_130 ();
 sg13g2_decap_8 FILLER_18_141 ();
 sg13g2_fill_2 FILLER_18_148 ();
 sg13g2_fill_1 FILLER_18_150 ();
 sg13g2_decap_8 FILLER_18_191 ();
 sg13g2_fill_2 FILLER_18_247 ();
 sg13g2_fill_1 FILLER_18_249 ();
 sg13g2_decap_8 FILLER_18_283 ();
 sg13g2_decap_4 FILLER_18_290 ();
 sg13g2_decap_8 FILLER_18_325 ();
 sg13g2_decap_8 FILLER_18_332 ();
 sg13g2_decap_4 FILLER_18_339 ();
 sg13g2_fill_2 FILLER_18_343 ();
 sg13g2_decap_8 FILLER_18_401 ();
 sg13g2_fill_1 FILLER_18_408 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_4 FILLER_19_7 ();
 sg13g2_fill_2 FILLER_19_11 ();
 sg13g2_decap_8 FILLER_19_65 ();
 sg13g2_decap_4 FILLER_19_72 ();
 sg13g2_decap_8 FILLER_19_84 ();
 sg13g2_decap_8 FILLER_19_110 ();
 sg13g2_fill_1 FILLER_19_117 ();
 sg13g2_decap_8 FILLER_19_137 ();
 sg13g2_decap_8 FILLER_19_144 ();
 sg13g2_fill_1 FILLER_19_165 ();
 sg13g2_fill_1 FILLER_19_180 ();
 sg13g2_decap_8 FILLER_19_188 ();
 sg13g2_decap_8 FILLER_19_195 ();
 sg13g2_decap_4 FILLER_19_202 ();
 sg13g2_fill_1 FILLER_19_206 ();
 sg13g2_fill_2 FILLER_19_238 ();
 sg13g2_decap_8 FILLER_19_250 ();
 sg13g2_fill_2 FILLER_19_257 ();
 sg13g2_fill_1 FILLER_19_259 ();
 sg13g2_decap_8 FILLER_19_281 ();
 sg13g2_decap_4 FILLER_19_288 ();
 sg13g2_fill_1 FILLER_19_292 ();
 sg13g2_fill_1 FILLER_19_307 ();
 sg13g2_decap_4 FILLER_19_327 ();
 sg13g2_fill_1 FILLER_19_331 ();
 sg13g2_decap_4 FILLER_19_371 ();
 sg13g2_fill_2 FILLER_19_375 ();
 sg13g2_decap_4 FILLER_19_404 ();
 sg13g2_fill_1 FILLER_19_408 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_decap_4 FILLER_20_57 ();
 sg13g2_decap_4 FILLER_20_74 ();
 sg13g2_decap_4 FILLER_20_115 ();
 sg13g2_fill_2 FILLER_20_119 ();
 sg13g2_decap_8 FILLER_20_125 ();
 sg13g2_decap_8 FILLER_20_132 ();
 sg13g2_decap_8 FILLER_20_139 ();
 sg13g2_fill_1 FILLER_20_146 ();
 sg13g2_decap_4 FILLER_20_174 ();
 sg13g2_fill_2 FILLER_20_188 ();
 sg13g2_decap_8 FILLER_20_195 ();
 sg13g2_fill_2 FILLER_20_202 ();
 sg13g2_fill_2 FILLER_20_227 ();
 sg13g2_fill_1 FILLER_20_229 ();
 sg13g2_fill_2 FILLER_20_233 ();
 sg13g2_fill_1 FILLER_20_235 ();
 sg13g2_decap_8 FILLER_20_272 ();
 sg13g2_decap_8 FILLER_20_279 ();
 sg13g2_decap_8 FILLER_20_286 ();
 sg13g2_decap_8 FILLER_20_293 ();
 sg13g2_decap_4 FILLER_20_342 ();
 sg13g2_fill_2 FILLER_20_346 ();
 sg13g2_decap_4 FILLER_20_353 ();
 sg13g2_decap_8 FILLER_20_394 ();
 sg13g2_decap_8 FILLER_20_401 ();
 sg13g2_fill_1 FILLER_20_408 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_fill_2 FILLER_21_7 ();
 sg13g2_fill_1 FILLER_21_9 ();
 sg13g2_fill_2 FILLER_21_78 ();
 sg13g2_decap_8 FILLER_21_134 ();
 sg13g2_fill_1 FILLER_21_141 ();
 sg13g2_fill_2 FILLER_21_204 ();
 sg13g2_fill_1 FILLER_21_206 ();
 sg13g2_decap_4 FILLER_21_226 ();
 sg13g2_fill_2 FILLER_21_230 ();
 sg13g2_decap_4 FILLER_21_273 ();
 sg13g2_fill_1 FILLER_21_277 ();
 sg13g2_fill_2 FILLER_21_305 ();
 sg13g2_fill_2 FILLER_21_334 ();
 sg13g2_fill_1 FILLER_21_336 ();
 sg13g2_fill_2 FILLER_21_341 ();
 sg13g2_fill_1 FILLER_21_365 ();
 sg13g2_fill_2 FILLER_21_381 ();
 sg13g2_decap_4 FILLER_21_403 ();
 sg13g2_fill_2 FILLER_21_407 ();
 sg13g2_fill_2 FILLER_22_0 ();
 sg13g2_fill_1 FILLER_22_2 ();
 sg13g2_fill_2 FILLER_22_44 ();
 sg13g2_fill_2 FILLER_22_73 ();
 sg13g2_fill_1 FILLER_22_75 ();
 sg13g2_decap_4 FILLER_22_137 ();
 sg13g2_decap_4 FILLER_22_161 ();
 sg13g2_fill_1 FILLER_22_174 ();
 sg13g2_decap_4 FILLER_22_212 ();
 sg13g2_fill_2 FILLER_22_231 ();
 sg13g2_decap_8 FILLER_22_273 ();
 sg13g2_fill_1 FILLER_22_280 ();
 sg13g2_fill_1 FILLER_22_323 ();
 sg13g2_fill_2 FILLER_22_338 ();
 sg13g2_fill_2 FILLER_22_350 ();
 sg13g2_fill_1 FILLER_22_352 ();
 sg13g2_fill_2 FILLER_22_363 ();
 sg13g2_fill_1 FILLER_22_365 ();
 sg13g2_fill_1 FILLER_22_376 ();
 sg13g2_fill_1 FILLER_22_386 ();
 sg13g2_fill_1 FILLER_22_408 ();
 sg13g2_decap_4 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_40 ();
 sg13g2_decap_8 FILLER_23_61 ();
 sg13g2_decap_8 FILLER_23_68 ();
 sg13g2_decap_4 FILLER_23_75 ();
 sg13g2_fill_2 FILLER_23_79 ();
 sg13g2_decap_4 FILLER_23_103 ();
 sg13g2_decap_8 FILLER_23_126 ();
 sg13g2_decap_8 FILLER_23_133 ();
 sg13g2_decap_8 FILLER_23_140 ();
 sg13g2_fill_1 FILLER_23_151 ();
 sg13g2_fill_2 FILLER_23_187 ();
 sg13g2_fill_1 FILLER_23_189 ();
 sg13g2_decap_8 FILLER_23_205 ();
 sg13g2_fill_1 FILLER_23_217 ();
 sg13g2_decap_8 FILLER_23_227 ();
 sg13g2_fill_1 FILLER_23_239 ();
 sg13g2_fill_2 FILLER_23_253 ();
 sg13g2_fill_1 FILLER_23_255 ();
 sg13g2_fill_1 FILLER_23_308 ();
 sg13g2_decap_4 FILLER_23_403 ();
 sg13g2_fill_2 FILLER_23_407 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_fill_2 FILLER_24_14 ();
 sg13g2_fill_1 FILLER_24_16 ();
 sg13g2_fill_1 FILLER_24_37 ();
 sg13g2_fill_2 FILLER_24_47 ();
 sg13g2_decap_8 FILLER_24_58 ();
 sg13g2_decap_8 FILLER_24_65 ();
 sg13g2_decap_8 FILLER_24_72 ();
 sg13g2_fill_1 FILLER_24_79 ();
 sg13g2_decap_8 FILLER_24_126 ();
 sg13g2_fill_2 FILLER_24_193 ();
 sg13g2_decap_8 FILLER_24_202 ();
 sg13g2_decap_4 FILLER_24_209 ();
 sg13g2_fill_1 FILLER_24_213 ();
 sg13g2_decap_8 FILLER_24_235 ();
 sg13g2_fill_2 FILLER_24_242 ();
 sg13g2_decap_8 FILLER_24_262 ();
 sg13g2_decap_4 FILLER_24_269 ();
 sg13g2_decap_4 FILLER_24_314 ();
 sg13g2_decap_8 FILLER_24_322 ();
 sg13g2_fill_2 FILLER_24_338 ();
 sg13g2_fill_1 FILLER_24_340 ();
 sg13g2_decap_4 FILLER_24_345 ();
 sg13g2_fill_1 FILLER_24_349 ();
 sg13g2_decap_4 FILLER_24_370 ();
 sg13g2_fill_1 FILLER_24_374 ();
 sg13g2_decap_8 FILLER_24_402 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_decap_4 FILLER_25_125 ();
 sg13g2_decap_8 FILLER_25_187 ();
 sg13g2_decap_8 FILLER_25_194 ();
 sg13g2_fill_2 FILLER_25_201 ();
 sg13g2_fill_1 FILLER_25_203 ();
 sg13g2_fill_1 FILLER_25_225 ();
 sg13g2_decap_8 FILLER_25_245 ();
 sg13g2_decap_8 FILLER_25_265 ();
 sg13g2_decap_4 FILLER_25_272 ();
 sg13g2_fill_2 FILLER_25_276 ();
 sg13g2_fill_1 FILLER_25_291 ();
 sg13g2_decap_8 FILLER_25_309 ();
 sg13g2_decap_8 FILLER_25_316 ();
 sg13g2_fill_2 FILLER_25_323 ();
 sg13g2_fill_1 FILLER_25_325 ();
 sg13g2_decap_8 FILLER_25_334 ();
 sg13g2_decap_4 FILLER_25_341 ();
 sg13g2_fill_1 FILLER_25_345 ();
 sg13g2_decap_4 FILLER_25_404 ();
 sg13g2_fill_1 FILLER_25_408 ();
 sg13g2_decap_4 FILLER_26_0 ();
 sg13g2_fill_2 FILLER_26_104 ();
 sg13g2_fill_1 FILLER_26_106 ();
 sg13g2_fill_2 FILLER_26_147 ();
 sg13g2_fill_2 FILLER_26_158 ();
 sg13g2_fill_1 FILLER_26_160 ();
 sg13g2_fill_2 FILLER_26_175 ();
 sg13g2_fill_1 FILLER_26_177 ();
 sg13g2_decap_8 FILLER_26_191 ();
 sg13g2_decap_8 FILLER_26_198 ();
 sg13g2_fill_1 FILLER_26_205 ();
 sg13g2_fill_2 FILLER_26_249 ();
 sg13g2_decap_8 FILLER_26_255 ();
 sg13g2_fill_1 FILLER_26_262 ();
 sg13g2_fill_2 FILLER_26_349 ();
 sg13g2_fill_1 FILLER_26_386 ();
 sg13g2_fill_1 FILLER_26_408 ();
 sg13g2_fill_2 FILLER_27_0 ();
 sg13g2_fill_1 FILLER_27_2 ();
 sg13g2_decap_4 FILLER_27_60 ();
 sg13g2_fill_2 FILLER_27_64 ();
 sg13g2_decap_8 FILLER_27_123 ();
 sg13g2_decap_8 FILLER_27_162 ();
 sg13g2_decap_8 FILLER_27_169 ();
 sg13g2_decap_8 FILLER_27_189 ();
 sg13g2_decap_8 FILLER_27_196 ();
 sg13g2_decap_8 FILLER_27_203 ();
 sg13g2_fill_1 FILLER_27_241 ();
 sg13g2_decap_4 FILLER_27_260 ();
 sg13g2_fill_1 FILLER_27_264 ();
 sg13g2_fill_2 FILLER_27_282 ();
 sg13g2_fill_2 FILLER_27_319 ();
 sg13g2_fill_2 FILLER_27_376 ();
 sg13g2_fill_2 FILLER_27_387 ();
 sg13g2_fill_2 FILLER_27_406 ();
 sg13g2_fill_1 FILLER_27_408 ();
 sg13g2_decap_4 FILLER_28_0 ();
 sg13g2_decap_4 FILLER_28_52 ();
 sg13g2_fill_2 FILLER_28_56 ();
 sg13g2_fill_1 FILLER_28_71 ();
 sg13g2_fill_2 FILLER_28_81 ();
 sg13g2_fill_1 FILLER_28_83 ();
 sg13g2_decap_8 FILLER_28_103 ();
 sg13g2_decap_8 FILLER_28_110 ();
 sg13g2_decap_8 FILLER_28_117 ();
 sg13g2_decap_4 FILLER_28_124 ();
 sg13g2_fill_1 FILLER_28_128 ();
 sg13g2_fill_1 FILLER_28_142 ();
 sg13g2_fill_2 FILLER_28_176 ();
 sg13g2_fill_1 FILLER_28_178 ();
 sg13g2_decap_8 FILLER_28_207 ();
 sg13g2_decap_4 FILLER_28_214 ();
 sg13g2_decap_4 FILLER_28_238 ();
 sg13g2_fill_1 FILLER_28_242 ();
 sg13g2_decap_8 FILLER_28_251 ();
 sg13g2_decap_8 FILLER_28_258 ();
 sg13g2_decap_8 FILLER_28_265 ();
 sg13g2_decap_8 FILLER_28_272 ();
 sg13g2_decap_8 FILLER_28_279 ();
 sg13g2_decap_4 FILLER_28_286 ();
 sg13g2_fill_2 FILLER_28_290 ();
 sg13g2_fill_2 FILLER_28_296 ();
 sg13g2_fill_1 FILLER_28_298 ();
 sg13g2_fill_2 FILLER_28_309 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_decap_8 FILLER_29_14 ();
 sg13g2_decap_4 FILLER_29_21 ();
 sg13g2_fill_1 FILLER_29_25 ();
 sg13g2_decap_4 FILLER_29_62 ();
 sg13g2_fill_2 FILLER_29_84 ();
 sg13g2_fill_2 FILLER_29_95 ();
 sg13g2_fill_1 FILLER_29_97 ();
 sg13g2_decap_8 FILLER_29_116 ();
 sg13g2_fill_2 FILLER_29_123 ();
 sg13g2_fill_1 FILLER_29_125 ();
 sg13g2_fill_1 FILLER_29_158 ();
 sg13g2_decap_4 FILLER_29_163 ();
 sg13g2_decap_4 FILLER_29_176 ();
 sg13g2_fill_1 FILLER_29_180 ();
 sg13g2_decap_8 FILLER_29_190 ();
 sg13g2_decap_8 FILLER_29_206 ();
 sg13g2_decap_4 FILLER_29_232 ();
 sg13g2_decap_8 FILLER_29_241 ();
 sg13g2_fill_2 FILLER_29_248 ();
 sg13g2_fill_1 FILLER_29_250 ();
 sg13g2_decap_8 FILLER_29_256 ();
 sg13g2_decap_8 FILLER_29_263 ();
 sg13g2_decap_4 FILLER_29_270 ();
 sg13g2_decap_8 FILLER_29_291 ();
 sg13g2_fill_1 FILLER_29_298 ();
 sg13g2_decap_4 FILLER_29_303 ();
 sg13g2_fill_2 FILLER_29_307 ();
 sg13g2_decap_4 FILLER_29_337 ();
 sg13g2_fill_1 FILLER_29_341 ();
 sg13g2_fill_1 FILLER_29_370 ();
 sg13g2_decap_8 FILLER_29_402 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_fill_2 FILLER_30_14 ();
 sg13g2_fill_1 FILLER_30_20 ();
 sg13g2_fill_1 FILLER_30_58 ();
 sg13g2_fill_2 FILLER_30_132 ();
 sg13g2_fill_1 FILLER_30_150 ();
 sg13g2_fill_1 FILLER_30_179 ();
 sg13g2_fill_2 FILLER_30_190 ();
 sg13g2_decap_4 FILLER_30_198 ();
 sg13g2_fill_2 FILLER_30_202 ();
 sg13g2_fill_1 FILLER_30_212 ();
 sg13g2_fill_1 FILLER_30_218 ();
 sg13g2_fill_2 FILLER_30_238 ();
 sg13g2_fill_1 FILLER_30_240 ();
 sg13g2_fill_1 FILLER_30_253 ();
 sg13g2_fill_2 FILLER_30_287 ();
 sg13g2_decap_8 FILLER_30_298 ();
 sg13g2_decap_8 FILLER_30_305 ();
 sg13g2_decap_8 FILLER_30_312 ();
 sg13g2_fill_1 FILLER_30_319 ();
 sg13g2_fill_1 FILLER_30_347 ();
 sg13g2_fill_2 FILLER_30_352 ();
 sg13g2_fill_1 FILLER_30_354 ();
 sg13g2_fill_1 FILLER_30_360 ();
 sg13g2_fill_1 FILLER_30_366 ();
 sg13g2_decap_8 FILLER_30_394 ();
 sg13g2_decap_8 FILLER_30_401 ();
 sg13g2_fill_1 FILLER_30_408 ();
 sg13g2_fill_2 FILLER_31_0 ();
 sg13g2_fill_1 FILLER_31_2 ();
 sg13g2_fill_1 FILLER_31_57 ();
 sg13g2_fill_1 FILLER_31_138 ();
 sg13g2_fill_2 FILLER_31_187 ();
 sg13g2_fill_1 FILLER_31_189 ();
 sg13g2_fill_1 FILLER_31_203 ();
 sg13g2_decap_4 FILLER_31_228 ();
 sg13g2_fill_1 FILLER_31_232 ();
 sg13g2_fill_2 FILLER_31_237 ();
 sg13g2_fill_2 FILLER_31_244 ();
 sg13g2_decap_8 FILLER_31_305 ();
 sg13g2_fill_2 FILLER_31_312 ();
 sg13g2_decap_4 FILLER_31_321 ();
 sg13g2_fill_2 FILLER_31_325 ();
 sg13g2_fill_1 FILLER_31_349 ();
 sg13g2_fill_2 FILLER_31_355 ();
 sg13g2_decap_4 FILLER_31_403 ();
 sg13g2_fill_2 FILLER_31_407 ();
 sg13g2_decap_4 FILLER_32_0 ();
 sg13g2_fill_2 FILLER_32_4 ();
 sg13g2_fill_2 FILLER_32_107 ();
 sg13g2_fill_1 FILLER_32_109 ();
 sg13g2_fill_2 FILLER_32_132 ();
 sg13g2_fill_2 FILLER_32_150 ();
 sg13g2_fill_1 FILLER_32_152 ();
 sg13g2_fill_1 FILLER_32_188 ();
 sg13g2_fill_2 FILLER_32_197 ();
 sg13g2_fill_1 FILLER_32_199 ();
 sg13g2_fill_1 FILLER_32_225 ();
 sg13g2_fill_1 FILLER_32_251 ();
 sg13g2_fill_2 FILLER_32_264 ();
 sg13g2_fill_1 FILLER_32_289 ();
 sg13g2_fill_1 FILLER_32_296 ();
 sg13g2_fill_1 FILLER_32_330 ();
 sg13g2_decap_4 FILLER_32_341 ();
 sg13g2_fill_1 FILLER_32_345 ();
 sg13g2_decap_4 FILLER_32_404 ();
 sg13g2_fill_1 FILLER_32_408 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_4 FILLER_33_7 ();
 sg13g2_fill_1 FILLER_33_65 ();
 sg13g2_decap_8 FILLER_33_140 ();
 sg13g2_decap_8 FILLER_33_147 ();
 sg13g2_decap_4 FILLER_33_154 ();
 sg13g2_fill_2 FILLER_33_194 ();
 sg13g2_fill_2 FILLER_33_215 ();
 sg13g2_decap_4 FILLER_33_228 ();
 sg13g2_fill_2 FILLER_33_232 ();
 sg13g2_decap_8 FILLER_33_242 ();
 sg13g2_fill_2 FILLER_33_270 ();
 sg13g2_fill_1 FILLER_33_272 ();
 sg13g2_fill_1 FILLER_33_293 ();
 sg13g2_fill_2 FILLER_33_326 ();
 sg13g2_fill_2 FILLER_33_345 ();
 sg13g2_fill_2 FILLER_33_352 ();
 sg13g2_fill_1 FILLER_33_354 ();
 sg13g2_fill_1 FILLER_33_365 ();
 sg13g2_fill_2 FILLER_33_371 ();
 sg13g2_fill_1 FILLER_33_408 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_fill_1 FILLER_34_14 ();
 sg13g2_fill_1 FILLER_34_43 ();
 sg13g2_fill_2 FILLER_34_49 ();
 sg13g2_fill_1 FILLER_34_78 ();
 sg13g2_fill_1 FILLER_34_133 ();
 sg13g2_decap_8 FILLER_34_142 ();
 sg13g2_decap_8 FILLER_34_149 ();
 sg13g2_decap_8 FILLER_34_156 ();
 sg13g2_fill_2 FILLER_34_163 ();
 sg13g2_fill_2 FILLER_34_184 ();
 sg13g2_fill_2 FILLER_34_191 ();
 sg13g2_fill_1 FILLER_34_193 ();
 sg13g2_decap_8 FILLER_34_199 ();
 sg13g2_decap_8 FILLER_34_206 ();
 sg13g2_decap_8 FILLER_34_213 ();
 sg13g2_fill_2 FILLER_34_230 ();
 sg13g2_decap_8 FILLER_34_241 ();
 sg13g2_decap_8 FILLER_34_248 ();
 sg13g2_fill_1 FILLER_34_255 ();
 sg13g2_fill_1 FILLER_34_268 ();
 sg13g2_fill_1 FILLER_34_278 ();
 sg13g2_fill_2 FILLER_34_294 ();
 sg13g2_fill_2 FILLER_34_332 ();
 sg13g2_fill_1 FILLER_34_334 ();
 sg13g2_fill_1 FILLER_34_343 ();
 sg13g2_fill_2 FILLER_34_361 ();
 sg13g2_fill_2 FILLER_34_407 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_fill_2 FILLER_35_7 ();
 sg13g2_fill_1 FILLER_35_49 ();
 sg13g2_fill_2 FILLER_35_92 ();
 sg13g2_decap_4 FILLER_35_148 ();
 sg13g2_fill_2 FILLER_35_152 ();
 sg13g2_fill_2 FILLER_35_207 ();
 sg13g2_fill_1 FILLER_35_209 ();
 sg13g2_decap_4 FILLER_35_223 ();
 sg13g2_fill_2 FILLER_35_267 ();
 sg13g2_fill_1 FILLER_35_269 ();
 sg13g2_fill_2 FILLER_35_335 ();
 sg13g2_decap_8 FILLER_35_400 ();
 sg13g2_fill_2 FILLER_35_407 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_fill_1 FILLER_36_14 ();
 sg13g2_fill_2 FILLER_36_132 ();
 sg13g2_fill_2 FILLER_36_143 ();
 sg13g2_fill_1 FILLER_36_145 ();
 sg13g2_fill_1 FILLER_36_209 ();
 sg13g2_fill_1 FILLER_36_265 ();
 sg13g2_decap_8 FILLER_36_401 ();
 sg13g2_fill_1 FILLER_36_408 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_fill_2 FILLER_37_7 ();
 sg13g2_fill_2 FILLER_37_34 ();
 sg13g2_fill_1 FILLER_37_54 ();
 sg13g2_fill_1 FILLER_37_132 ();
 sg13g2_decap_8 FILLER_37_226 ();
 sg13g2_fill_1 FILLER_37_270 ();
 sg13g2_fill_2 FILLER_37_304 ();
 sg13g2_fill_1 FILLER_37_318 ();
 sg13g2_decap_4 FILLER_37_405 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_4 FILLER_38_7 ();
 sg13g2_fill_1 FILLER_38_11 ();
 sg13g2_fill_1 FILLER_38_74 ();
 sg13g2_fill_2 FILLER_38_122 ();
 sg13g2_fill_1 FILLER_38_124 ();
 sg13g2_fill_2 FILLER_38_134 ();
 sg13g2_fill_2 FILLER_38_175 ();
 sg13g2_fill_1 FILLER_38_177 ();
 sg13g2_fill_2 FILLER_38_191 ();
 sg13g2_fill_1 FILLER_38_193 ();
 sg13g2_fill_2 FILLER_38_211 ();
 sg13g2_fill_1 FILLER_38_213 ();
 sg13g2_decap_8 FILLER_38_223 ();
 sg13g2_decap_8 FILLER_38_230 ();
 sg13g2_fill_1 FILLER_38_237 ();
 sg13g2_fill_2 FILLER_38_246 ();
 sg13g2_decap_8 FILLER_38_252 ();
 sg13g2_decap_4 FILLER_38_259 ();
 sg13g2_fill_1 FILLER_38_263 ();
 sg13g2_decap_8 FILLER_38_383 ();
 sg13g2_decap_8 FILLER_38_390 ();
 sg13g2_decap_8 FILLER_38_397 ();
 sg13g2_decap_4 FILLER_38_404 ();
 sg13g2_fill_1 FILLER_38_408 ();
 assign uio_oe[0] = net14;
 assign uio_oe[1] = net15;
 assign uio_oe[2] = net16;
 assign uio_oe[3] = net17;
 assign uio_oe[4] = net18;
 assign uio_oe[5] = net19;
 assign uio_oe[6] = net20;
 assign uio_oe[7] = net21;
 assign uio_out[0] = net22;
 assign uio_out[1] = net23;
 assign uio_out[2] = net24;
 assign uio_out[3] = net25;
 assign uio_out[4] = net26;
 assign uio_out[5] = net27;
 assign uio_out[6] = net28;
 assign uio_out[7] = net29;
endmodule
