module tt_um_ECM24_serv_soc_top (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _00000_;
 wire _00001_;
 wire _00002_;
 wire _00003_;
 wire _00004_;
 wire _00005_;
 wire _00006_;
 wire _00007_;
 wire _00008_;
 wire _00009_;
 wire _00010_;
 wire _00011_;
 wire _00012_;
 wire _00013_;
 wire _00014_;
 wire _00015_;
 wire _00016_;
 wire _00017_;
 wire _00018_;
 wire _00019_;
 wire _00020_;
 wire _00021_;
 wire _00022_;
 wire _00023_;
 wire _00024_;
 wire _00025_;
 wire _00026_;
 wire _00027_;
 wire _00028_;
 wire _00029_;
 wire _00030_;
 wire _00031_;
 wire _00032_;
 wire _00033_;
 wire _00034_;
 wire _00035_;
 wire _00036_;
 wire _00037_;
 wire _00038_;
 wire _00039_;
 wire _00040_;
 wire _00041_;
 wire _00042_;
 wire _00043_;
 wire _00044_;
 wire _00045_;
 wire _00046_;
 wire _00047_;
 wire _00048_;
 wire _00049_;
 wire _00050_;
 wire _00051_;
 wire _00052_;
 wire _00053_;
 wire _00054_;
 wire _00055_;
 wire _00056_;
 wire _00057_;
 wire _00058_;
 wire _00059_;
 wire _00060_;
 wire _00061_;
 wire _00062_;
 wire _00063_;
 wire _00064_;
 wire _00065_;
 wire _00066_;
 wire _00067_;
 wire _00068_;
 wire _00069_;
 wire _00070_;
 wire clk_regs;
 wire _00072_;
 wire _00073_;
 wire _00074_;
 wire _00075_;
 wire _00076_;
 wire _00077_;
 wire _00078_;
 wire _00079_;
 wire _00080_;
 wire _00081_;
 wire _00082_;
 wire _00083_;
 wire _00084_;
 wire _00085_;
 wire _00086_;
 wire _00087_;
 wire _00088_;
 wire _00089_;
 wire _00090_;
 wire _00091_;
 wire _00092_;
 wire _00093_;
 wire _00094_;
 wire _00095_;
 wire _00096_;
 wire _00097_;
 wire _00098_;
 wire _00099_;
 wire _00100_;
 wire _00101_;
 wire _00102_;
 wire _00103_;
 wire _00104_;
 wire _00105_;
 wire _00106_;
 wire _00107_;
 wire _00108_;
 wire _00109_;
 wire _00110_;
 wire _00111_;
 wire _00112_;
 wire _00113_;
 wire _00114_;
 wire _00115_;
 wire _00116_;
 wire _00117_;
 wire _00118_;
 wire _00119_;
 wire _00120_;
 wire _00121_;
 wire _00122_;
 wire _00123_;
 wire _00124_;
 wire _00125_;
 wire _00126_;
 wire _00127_;
 wire _00128_;
 wire _00129_;
 wire _00130_;
 wire _00131_;
 wire _00132_;
 wire _00133_;
 wire _00134_;
 wire _00135_;
 wire _00136_;
 wire _00137_;
 wire _00138_;
 wire _00139_;
 wire _00140_;
 wire _00141_;
 wire _00142_;
 wire _00143_;
 wire _00144_;
 wire _00145_;
 wire _00146_;
 wire _00147_;
 wire _00148_;
 wire _00149_;
 wire _00150_;
 wire _00151_;
 wire _00152_;
 wire _00153_;
 wire _00154_;
 wire _00155_;
 wire _00156_;
 wire _00157_;
 wire _00158_;
 wire _00159_;
 wire _00160_;
 wire _00161_;
 wire _00162_;
 wire _00163_;
 wire _00164_;
 wire _00165_;
 wire _00166_;
 wire _00167_;
 wire _00168_;
 wire _00169_;
 wire _00170_;
 wire _00171_;
 wire _00172_;
 wire _00173_;
 wire _00174_;
 wire _00175_;
 wire _00176_;
 wire _00177_;
 wire _00178_;
 wire _00179_;
 wire _00180_;
 wire _00181_;
 wire _00182_;
 wire _00183_;
 wire _00184_;
 wire _00185_;
 wire _00186_;
 wire _00187_;
 wire _00188_;
 wire _00189_;
 wire _00190_;
 wire _00191_;
 wire _00192_;
 wire _00193_;
 wire _00194_;
 wire _00195_;
 wire _00196_;
 wire _00197_;
 wire _00198_;
 wire _00199_;
 wire _00200_;
 wire _00201_;
 wire _00202_;
 wire _00203_;
 wire _00204_;
 wire _00205_;
 wire _00206_;
 wire _00207_;
 wire _00208_;
 wire _00209_;
 wire _00210_;
 wire _00211_;
 wire _00212_;
 wire _00213_;
 wire _00214_;
 wire _00215_;
 wire _00216_;
 wire _00217_;
 wire _00218_;
 wire _00219_;
 wire _00220_;
 wire _00221_;
 wire _00222_;
 wire _00223_;
 wire _00224_;
 wire _00225_;
 wire _00226_;
 wire _00227_;
 wire _00228_;
 wire _00229_;
 wire _00230_;
 wire _00231_;
 wire _00232_;
 wire _00233_;
 wire _00234_;
 wire _00235_;
 wire _00236_;
 wire _00237_;
 wire _00238_;
 wire _00239_;
 wire _00240_;
 wire _00241_;
 wire _00242_;
 wire _00243_;
 wire _00244_;
 wire _00245_;
 wire _00246_;
 wire _00247_;
 wire _00248_;
 wire _00249_;
 wire _00250_;
 wire _00251_;
 wire _00252_;
 wire _00253_;
 wire _00254_;
 wire _00255_;
 wire _00256_;
 wire _00257_;
 wire _00258_;
 wire _00259_;
 wire _00260_;
 wire _00261_;
 wire _00262_;
 wire _00263_;
 wire _00264_;
 wire _00265_;
 wire _00266_;
 wire _00267_;
 wire _00268_;
 wire _00269_;
 wire _00270_;
 wire _00271_;
 wire _00272_;
 wire _00273_;
 wire _00274_;
 wire _00275_;
 wire _00276_;
 wire _00277_;
 wire _00278_;
 wire _00279_;
 wire _00280_;
 wire _00281_;
 wire _00282_;
 wire _00283_;
 wire _00284_;
 wire _00285_;
 wire _00286_;
 wire _00287_;
 wire _00288_;
 wire _00289_;
 wire _00290_;
 wire _00291_;
 wire _00292_;
 wire _00293_;
 wire _00294_;
 wire _00295_;
 wire _00296_;
 wire _00297_;
 wire _00298_;
 wire _00299_;
 wire _00300_;
 wire _00301_;
 wire _00302_;
 wire _00303_;
 wire _00304_;
 wire _00305_;
 wire _00306_;
 wire _00307_;
 wire _00308_;
 wire _00309_;
 wire _00310_;
 wire _00311_;
 wire _00312_;
 wire _00313_;
 wire _00314_;
 wire _00315_;
 wire _00316_;
 wire _00317_;
 wire _00318_;
 wire _00319_;
 wire _00320_;
 wire _00321_;
 wire _00322_;
 wire _00323_;
 wire _00324_;
 wire _00325_;
 wire _00326_;
 wire _00327_;
 wire _00328_;
 wire _00329_;
 wire _00330_;
 wire _00331_;
 wire _00332_;
 wire _00333_;
 wire _00334_;
 wire _00335_;
 wire _00336_;
 wire _00337_;
 wire _00338_;
 wire _00339_;
 wire _00340_;
 wire _00341_;
 wire _00342_;
 wire _00343_;
 wire _00344_;
 wire _00345_;
 wire _00346_;
 wire _00347_;
 wire _00348_;
 wire _00349_;
 wire _00350_;
 wire _00351_;
 wire _00352_;
 wire _00353_;
 wire _00354_;
 wire _00355_;
 wire _00356_;
 wire _00357_;
 wire _00358_;
 wire _00359_;
 wire _00360_;
 wire _00361_;
 wire _00362_;
 wire _00363_;
 wire _00364_;
 wire _00365_;
 wire _00366_;
 wire _00367_;
 wire _00368_;
 wire _00369_;
 wire _00370_;
 wire _00371_;
 wire _00372_;
 wire _00373_;
 wire _00374_;
 wire _00375_;
 wire _00376_;
 wire _00377_;
 wire _00378_;
 wire _00379_;
 wire _00380_;
 wire _00381_;
 wire _00382_;
 wire _00383_;
 wire _00384_;
 wire _00385_;
 wire _00386_;
 wire _00387_;
 wire _00388_;
 wire _00389_;
 wire _00390_;
 wire _00391_;
 wire _00392_;
 wire _00393_;
 wire _00394_;
 wire _00395_;
 wire _00396_;
 wire _00397_;
 wire _00398_;
 wire _00399_;
 wire _00400_;
 wire _00401_;
 wire _00402_;
 wire _00403_;
 wire _00404_;
 wire _00405_;
 wire _00406_;
 wire _00407_;
 wire _00408_;
 wire _00409_;
 wire _00410_;
 wire _00411_;
 wire _00412_;
 wire _00413_;
 wire _00414_;
 wire _00415_;
 wire _00416_;
 wire _00417_;
 wire _00418_;
 wire _00419_;
 wire _00420_;
 wire _00421_;
 wire _00422_;
 wire _00423_;
 wire _00424_;
 wire _00425_;
 wire _00426_;
 wire _00427_;
 wire _00428_;
 wire _00429_;
 wire _00430_;
 wire _00431_;
 wire _00432_;
 wire _00433_;
 wire _00434_;
 wire _00435_;
 wire _00436_;
 wire _00437_;
 wire _00438_;
 wire _00439_;
 wire _00440_;
 wire _00441_;
 wire _00442_;
 wire _00443_;
 wire _00444_;
 wire _00445_;
 wire _00446_;
 wire _00447_;
 wire _00448_;
 wire _00449_;
 wire _00450_;
 wire _00451_;
 wire _00452_;
 wire _00453_;
 wire _00454_;
 wire _00455_;
 wire _00456_;
 wire _00457_;
 wire _00458_;
 wire _00459_;
 wire _00460_;
 wire _00461_;
 wire _00462_;
 wire _00463_;
 wire _00464_;
 wire _00465_;
 wire _00466_;
 wire _00467_;
 wire _00468_;
 wire _00469_;
 wire _00470_;
 wire _00471_;
 wire _00472_;
 wire _00473_;
 wire _00474_;
 wire _00475_;
 wire _00476_;
 wire _00477_;
 wire _00478_;
 wire _00479_;
 wire _00480_;
 wire _00481_;
 wire _00482_;
 wire _00483_;
 wire _00484_;
 wire _00485_;
 wire _00486_;
 wire _00487_;
 wire _00488_;
 wire _00489_;
 wire _00490_;
 wire _00491_;
 wire _00492_;
 wire _00493_;
 wire _00494_;
 wire _00495_;
 wire _00496_;
 wire _00497_;
 wire _00498_;
 wire _00499_;
 wire _00500_;
 wire _00501_;
 wire _00502_;
 wire _00503_;
 wire _00504_;
 wire _00505_;
 wire _00506_;
 wire _00507_;
 wire _00508_;
 wire _00509_;
 wire _00510_;
 wire _00511_;
 wire _00512_;
 wire _00513_;
 wire _00514_;
 wire _00515_;
 wire _00516_;
 wire _00517_;
 wire _00518_;
 wire _00519_;
 wire _00520_;
 wire _00521_;
 wire _00522_;
 wire _00523_;
 wire _00524_;
 wire _00525_;
 wire _00526_;
 wire _00527_;
 wire _00528_;
 wire _00529_;
 wire _00530_;
 wire _00531_;
 wire _00532_;
 wire _00533_;
 wire _00534_;
 wire _00535_;
 wire _00536_;
 wire _00537_;
 wire _00538_;
 wire _00539_;
 wire _00540_;
 wire _00541_;
 wire _00542_;
 wire _00543_;
 wire _00544_;
 wire _00545_;
 wire _00546_;
 wire _00547_;
 wire _00548_;
 wire _00549_;
 wire _00550_;
 wire _00551_;
 wire _00552_;
 wire _00553_;
 wire _00554_;
 wire _00555_;
 wire _00556_;
 wire _00557_;
 wire _00558_;
 wire _00559_;
 wire _00560_;
 wire _00561_;
 wire _00562_;
 wire _00563_;
 wire _00564_;
 wire _00565_;
 wire _00566_;
 wire _00567_;
 wire _00568_;
 wire _00569_;
 wire _00570_;
 wire _00571_;
 wire _00572_;
 wire _00573_;
 wire _00574_;
 wire _00575_;
 wire _00576_;
 wire _00577_;
 wire _00578_;
 wire _00579_;
 wire _00580_;
 wire _00581_;
 wire _00582_;
 wire _00583_;
 wire _00584_;
 wire _00585_;
 wire _00586_;
 wire _00587_;
 wire _00588_;
 wire _00589_;
 wire _00590_;
 wire _00591_;
 wire _00592_;
 wire _00593_;
 wire _00594_;
 wire _00595_;
 wire _00596_;
 wire _00597_;
 wire _00598_;
 wire _00599_;
 wire _00600_;
 wire _00601_;
 wire _00602_;
 wire _00603_;
 wire _00604_;
 wire _00605_;
 wire _00606_;
 wire _00607_;
 wire _00608_;
 wire _00609_;
 wire _00610_;
 wire _00611_;
 wire _00612_;
 wire _00613_;
 wire _00614_;
 wire _00615_;
 wire _00616_;
 wire _00617_;
 wire _00618_;
 wire _00619_;
 wire _00620_;
 wire _00621_;
 wire _00622_;
 wire _00623_;
 wire _00624_;
 wire _00625_;
 wire _00626_;
 wire _00627_;
 wire _00628_;
 wire _00629_;
 wire _00630_;
 wire _00631_;
 wire _00632_;
 wire _00633_;
 wire _00634_;
 wire _00635_;
 wire _00636_;
 wire _00637_;
 wire _00638_;
 wire _00639_;
 wire _00640_;
 wire _00641_;
 wire _00642_;
 wire _00643_;
 wire _00644_;
 wire _00645_;
 wire _00646_;
 wire _00647_;
 wire _00648_;
 wire _00649_;
 wire _00650_;
 wire _00651_;
 wire _00652_;
 wire _00653_;
 wire _00654_;
 wire _00655_;
 wire _00656_;
 wire _00657_;
 wire _00658_;
 wire _00659_;
 wire _00660_;
 wire _00661_;
 wire _00662_;
 wire _00663_;
 wire _00664_;
 wire _00665_;
 wire _00666_;
 wire _00667_;
 wire _00668_;
 wire _00669_;
 wire _00670_;
 wire _00671_;
 wire _00672_;
 wire _00673_;
 wire _00674_;
 wire _00675_;
 wire _00676_;
 wire _00677_;
 wire _00678_;
 wire _00679_;
 wire _00680_;
 wire _00681_;
 wire _00682_;
 wire _00683_;
 wire _00684_;
 wire _00685_;
 wire _00686_;
 wire _00687_;
 wire _00688_;
 wire _00689_;
 wire _00690_;
 wire _00691_;
 wire _00692_;
 wire _00693_;
 wire _00694_;
 wire _00695_;
 wire _00696_;
 wire _00697_;
 wire _00698_;
 wire _00699_;
 wire _00700_;
 wire _00701_;
 wire _00702_;
 wire _00703_;
 wire _00704_;
 wire _00705_;
 wire _00706_;
 wire _00707_;
 wire _00708_;
 wire _00709_;
 wire _00710_;
 wire _00711_;
 wire _00712_;
 wire _00713_;
 wire _00714_;
 wire _00715_;
 wire _00716_;
 wire _00717_;
 wire _00718_;
 wire _00719_;
 wire _00720_;
 wire _00721_;
 wire _00722_;
 wire _00723_;
 wire _00724_;
 wire _00725_;
 wire _00726_;
 wire _00727_;
 wire _00728_;
 wire _00729_;
 wire _00730_;
 wire _00731_;
 wire _00732_;
 wire _00733_;
 wire _00734_;
 wire _00735_;
 wire _00736_;
 wire _00737_;
 wire _00738_;
 wire _00739_;
 wire _00740_;
 wire _00741_;
 wire _00742_;
 wire _00743_;
 wire _00744_;
 wire _00745_;
 wire _00746_;
 wire _00747_;
 wire _00748_;
 wire _00749_;
 wire _00750_;
 wire _00751_;
 wire _00752_;
 wire _00753_;
 wire _00754_;
 wire _00755_;
 wire _00756_;
 wire _00757_;
 wire _00758_;
 wire _00759_;
 wire _00760_;
 wire _00761_;
 wire _00762_;
 wire _00763_;
 wire _00764_;
 wire _00765_;
 wire _00766_;
 wire _00767_;
 wire _00768_;
 wire _00769_;
 wire _00770_;
 wire _00771_;
 wire _00772_;
 wire _00773_;
 wire _00774_;
 wire _00775_;
 wire _00776_;
 wire _00777_;
 wire _00778_;
 wire _00779_;
 wire _00780_;
 wire _00781_;
 wire _00782_;
 wire _00783_;
 wire _00784_;
 wire _00785_;
 wire _00786_;
 wire _00787_;
 wire _00788_;
 wire _00789_;
 wire _00790_;
 wire _00791_;
 wire _00792_;
 wire _00793_;
 wire _00794_;
 wire _00795_;
 wire _00796_;
 wire _00797_;
 wire _00798_;
 wire _00799_;
 wire _00800_;
 wire _00801_;
 wire _00802_;
 wire _00803_;
 wire _00804_;
 wire _00805_;
 wire _00806_;
 wire _00807_;
 wire _00808_;
 wire _00809_;
 wire _00810_;
 wire _00811_;
 wire _00812_;
 wire _00813_;
 wire _00814_;
 wire _00815_;
 wire _00816_;
 wire _00817_;
 wire _00818_;
 wire _00819_;
 wire _00820_;
 wire _00821_;
 wire _00822_;
 wire _00823_;
 wire _00824_;
 wire _00825_;
 wire _00826_;
 wire _00827_;
 wire _00828_;
 wire _00829_;
 wire _00830_;
 wire _00831_;
 wire _00832_;
 wire _00833_;
 wire _00834_;
 wire _00835_;
 wire _00836_;
 wire _00837_;
 wire _00838_;
 wire _00839_;
 wire _00840_;
 wire _00841_;
 wire _00842_;
 wire _00843_;
 wire _00844_;
 wire _00845_;
 wire _00846_;
 wire _00847_;
 wire _00848_;
 wire _00849_;
 wire _00850_;
 wire _00851_;
 wire _00852_;
 wire _00853_;
 wire _00854_;
 wire _00855_;
 wire _00856_;
 wire _00857_;
 wire _00858_;
 wire _00859_;
 wire _00860_;
 wire _00861_;
 wire _00862_;
 wire _00863_;
 wire _00864_;
 wire _00865_;
 wire _00866_;
 wire _00867_;
 wire _00868_;
 wire _00869_;
 wire _00870_;
 wire _00871_;
 wire _00872_;
 wire _00873_;
 wire _00874_;
 wire _00875_;
 wire _00876_;
 wire _00877_;
 wire _00878_;
 wire _00879_;
 wire _00880_;
 wire _00881_;
 wire _00882_;
 wire _00883_;
 wire _00884_;
 wire _00885_;
 wire _00886_;
 wire _00887_;
 wire _00888_;
 wire _00889_;
 wire _00890_;
 wire _00891_;
 wire _00892_;
 wire _00893_;
 wire _00894_;
 wire _00895_;
 wire _00896_;
 wire _00897_;
 wire _00898_;
 wire _00899_;
 wire _00900_;
 wire _00901_;
 wire _00902_;
 wire _00903_;
 wire _00904_;
 wire _00905_;
 wire _00906_;
 wire _00907_;
 wire _00908_;
 wire _00909_;
 wire _00910_;
 wire _00911_;
 wire _00912_;
 wire _00913_;
 wire _00914_;
 wire _00915_;
 wire _00916_;
 wire _00917_;
 wire _00918_;
 wire _00919_;
 wire _00920_;
 wire _00921_;
 wire _00922_;
 wire _00923_;
 wire _00924_;
 wire _00925_;
 wire _00926_;
 wire _00927_;
 wire _00928_;
 wire _00929_;
 wire _00930_;
 wire _00931_;
 wire _00932_;
 wire _00933_;
 wire _00934_;
 wire _00935_;
 wire _00936_;
 wire _00937_;
 wire _00938_;
 wire _00939_;
 wire _00940_;
 wire _00941_;
 wire _00942_;
 wire _00943_;
 wire _00944_;
 wire _00945_;
 wire _00946_;
 wire _00947_;
 wire _00948_;
 wire _00949_;
 wire _00950_;
 wire _00951_;
 wire _00952_;
 wire _00953_;
 wire _00954_;
 wire _00955_;
 wire _00956_;
 wire _00957_;
 wire _00958_;
 wire _00959_;
 wire _00960_;
 wire _00961_;
 wire _00962_;
 wire _00963_;
 wire _00964_;
 wire _00965_;
 wire _00966_;
 wire _00967_;
 wire _00968_;
 wire _00969_;
 wire _00970_;
 wire _00971_;
 wire _00972_;
 wire _00973_;
 wire _00974_;
 wire _00975_;
 wire _00976_;
 wire _00977_;
 wire _00978_;
 wire _00979_;
 wire _00980_;
 wire _00981_;
 wire _00982_;
 wire _00983_;
 wire _00984_;
 wire _00985_;
 wire _00986_;
 wire _00987_;
 wire _00988_;
 wire _00989_;
 wire _00990_;
 wire _00991_;
 wire _00992_;
 wire _00993_;
 wire _00994_;
 wire _00995_;
 wire _00996_;
 wire _00997_;
 wire _00998_;
 wire _00999_;
 wire _01000_;
 wire _01001_;
 wire _01002_;
 wire _01003_;
 wire _01004_;
 wire _01005_;
 wire _01006_;
 wire _01007_;
 wire _01008_;
 wire _01009_;
 wire _01010_;
 wire _01011_;
 wire _01012_;
 wire _01013_;
 wire _01014_;
 wire _01015_;
 wire _01016_;
 wire _01017_;
 wire _01018_;
 wire _01019_;
 wire _01020_;
 wire _01021_;
 wire _01022_;
 wire _01023_;
 wire _01024_;
 wire _01025_;
 wire _01026_;
 wire _01027_;
 wire _01028_;
 wire _01029_;
 wire _01030_;
 wire _01031_;
 wire _01032_;
 wire _01033_;
 wire _01034_;
 wire _01035_;
 wire _01036_;
 wire _01037_;
 wire _01038_;
 wire _01039_;
 wire _01040_;
 wire _01041_;
 wire _01042_;
 wire _01043_;
 wire _01044_;
 wire _01045_;
 wire _01046_;
 wire _01047_;
 wire _01048_;
 wire _01049_;
 wire _01050_;
 wire _01051_;
 wire _01052_;
 wire _01053_;
 wire _01054_;
 wire _01055_;
 wire _01056_;
 wire _01057_;
 wire _01058_;
 wire _01059_;
 wire _01060_;
 wire _01061_;
 wire _01062_;
 wire _01063_;
 wire _01064_;
 wire _01065_;
 wire _01066_;
 wire _01067_;
 wire _01068_;
 wire _01069_;
 wire _01070_;
 wire _01071_;
 wire _01072_;
 wire _01073_;
 wire _01074_;
 wire _01075_;
 wire _01076_;
 wire _01077_;
 wire _01078_;
 wire _01079_;
 wire _01080_;
 wire _01081_;
 wire _01082_;
 wire _01083_;
 wire _01084_;
 wire _01085_;
 wire _01086_;
 wire _01087_;
 wire _01088_;
 wire _01089_;
 wire _01090_;
 wire _01091_;
 wire _01092_;
 wire _01093_;
 wire _01094_;
 wire _01095_;
 wire _01096_;
 wire _01097_;
 wire _01098_;
 wire _01099_;
 wire _01100_;
 wire _01101_;
 wire _01102_;
 wire _01103_;
 wire _01104_;
 wire _01105_;
 wire _01106_;
 wire _01107_;
 wire _01108_;
 wire _01109_;
 wire _01110_;
 wire _01111_;
 wire _01112_;
 wire _01113_;
 wire _01114_;
 wire _01115_;
 wire _01116_;
 wire _01117_;
 wire _01118_;
 wire _01119_;
 wire _01120_;
 wire _01121_;
 wire _01122_;
 wire _01123_;
 wire _01124_;
 wire _01125_;
 wire _01126_;
 wire _01127_;
 wire _01128_;
 wire _01129_;
 wire _01130_;
 wire _01131_;
 wire _01132_;
 wire _01133_;
 wire _01134_;
 wire _01135_;
 wire _01136_;
 wire _01137_;
 wire _01138_;
 wire _01139_;
 wire _01140_;
 wire _01141_;
 wire _01142_;
 wire _01143_;
 wire _01144_;
 wire _01145_;
 wire _01146_;
 wire _01147_;
 wire _01148_;
 wire _01149_;
 wire _01150_;
 wire _01151_;
 wire _01152_;
 wire _01153_;
 wire _01154_;
 wire _01155_;
 wire _01156_;
 wire _01157_;
 wire _01158_;
 wire _01159_;
 wire _01160_;
 wire _01161_;
 wire _01162_;
 wire _01163_;
 wire _01164_;
 wire _01165_;
 wire _01166_;
 wire _01167_;
 wire _01168_;
 wire _01169_;
 wire _01170_;
 wire _01171_;
 wire _01172_;
 wire _01173_;
 wire _01174_;
 wire _01175_;
 wire _01176_;
 wire _01177_;
 wire _01178_;
 wire _01179_;
 wire _01180_;
 wire _01181_;
 wire _01182_;
 wire _01183_;
 wire _01184_;
 wire _01185_;
 wire _01186_;
 wire _01187_;
 wire _01188_;
 wire _01189_;
 wire _01190_;
 wire _01191_;
 wire _01192_;
 wire _01193_;
 wire _01194_;
 wire _01195_;
 wire _01196_;
 wire _01197_;
 wire _01198_;
 wire _01199_;
 wire _01200_;
 wire _01201_;
 wire _01202_;
 wire _01203_;
 wire _01204_;
 wire _01205_;
 wire _01206_;
 wire _01207_;
 wire _01208_;
 wire _01209_;
 wire _01210_;
 wire _01211_;
 wire _01212_;
 wire _01213_;
 wire _01214_;
 wire _01215_;
 wire _01216_;
 wire _01217_;
 wire _01218_;
 wire _01219_;
 wire _01220_;
 wire _01221_;
 wire _01222_;
 wire _01223_;
 wire _01224_;
 wire _01225_;
 wire _01226_;
 wire _01227_;
 wire _01228_;
 wire _01229_;
 wire _01230_;
 wire _01231_;
 wire _01232_;
 wire _01233_;
 wire _01234_;
 wire _01235_;
 wire _01236_;
 wire _01237_;
 wire _01238_;
 wire _01239_;
 wire _01240_;
 wire _01241_;
 wire _01242_;
 wire _01243_;
 wire _01244_;
 wire _01245_;
 wire _01246_;
 wire _01247_;
 wire _01248_;
 wire _01249_;
 wire _01250_;
 wire _01251_;
 wire _01252_;
 wire _01253_;
 wire _01254_;
 wire _01255_;
 wire _01256_;
 wire _01257_;
 wire _01258_;
 wire _01259_;
 wire _01260_;
 wire _01261_;
 wire _01262_;
 wire _01263_;
 wire _01264_;
 wire _01265_;
 wire _01266_;
 wire _01267_;
 wire _01268_;
 wire _01269_;
 wire _01270_;
 wire _01271_;
 wire _01272_;
 wire _01273_;
 wire _01274_;
 wire _01275_;
 wire _01276_;
 wire _01277_;
 wire _01278_;
 wire _01279_;
 wire _01280_;
 wire _01281_;
 wire _01282_;
 wire _01283_;
 wire _01284_;
 wire _01285_;
 wire _01286_;
 wire _01287_;
 wire _01288_;
 wire _01289_;
 wire _01290_;
 wire _01291_;
 wire _01292_;
 wire _01293_;
 wire _01294_;
 wire _01295_;
 wire _01296_;
 wire _01297_;
 wire _01298_;
 wire _01299_;
 wire _01300_;
 wire _01301_;
 wire _01302_;
 wire _01303_;
 wire _01304_;
 wire _01305_;
 wire _01306_;
 wire _01307_;
 wire _01308_;
 wire _01309_;
 wire _01310_;
 wire _01311_;
 wire _01312_;
 wire _01313_;
 wire _01314_;
 wire _01315_;
 wire _01316_;
 wire _01317_;
 wire _01318_;
 wire _01319_;
 wire _01320_;
 wire _01321_;
 wire _01322_;
 wire _01323_;
 wire _01324_;
 wire _01325_;
 wire _01326_;
 wire _01327_;
 wire _01328_;
 wire _01329_;
 wire _01330_;
 wire _01331_;
 wire _01332_;
 wire _01333_;
 wire _01334_;
 wire _01335_;
 wire _01336_;
 wire _01337_;
 wire _01338_;
 wire _01339_;
 wire _01340_;
 wire _01341_;
 wire _01342_;
 wire _01343_;
 wire _01344_;
 wire _01345_;
 wire _01346_;
 wire _01347_;
 wire _01348_;
 wire _01349_;
 wire _01350_;
 wire _01351_;
 wire _01352_;
 wire _01353_;
 wire _01354_;
 wire _01355_;
 wire _01356_;
 wire _01357_;
 wire _01358_;
 wire _01359_;
 wire _01360_;
 wire _01361_;
 wire _01362_;
 wire _01363_;
 wire _01364_;
 wire _01365_;
 wire _01366_;
 wire _01367_;
 wire _01368_;
 wire _01369_;
 wire _01370_;
 wire _01371_;
 wire _01372_;
 wire _01373_;
 wire _01374_;
 wire _01375_;
 wire _01376_;
 wire _01377_;
 wire _01378_;
 wire _01379_;
 wire _01380_;
 wire _01381_;
 wire _01382_;
 wire _01383_;
 wire _01384_;
 wire _01385_;
 wire _01386_;
 wire _01387_;
 wire _01388_;
 wire _01389_;
 wire _01390_;
 wire _01391_;
 wire _01392_;
 wire _01393_;
 wire _01394_;
 wire _01395_;
 wire _01396_;
 wire _01397_;
 wire _01398_;
 wire _01399_;
 wire _01400_;
 wire _01401_;
 wire _01402_;
 wire _01403_;
 wire _01404_;
 wire _01405_;
 wire _01406_;
 wire _01407_;
 wire _01408_;
 wire _01409_;
 wire _01410_;
 wire _01411_;
 wire _01412_;
 wire _01413_;
 wire _01414_;
 wire _01415_;
 wire _01416_;
 wire _01417_;
 wire _01418_;
 wire _01419_;
 wire _01420_;
 wire _01421_;
 wire _01422_;
 wire _01423_;
 wire _01424_;
 wire _01425_;
 wire _01426_;
 wire _01427_;
 wire _01428_;
 wire _01429_;
 wire _01430_;
 wire _01431_;
 wire _01432_;
 wire _01433_;
 wire _01434_;
 wire _01435_;
 wire _01436_;
 wire _01437_;
 wire _01438_;
 wire _01439_;
 wire _01440_;
 wire _01441_;
 wire _01442_;
 wire _01443_;
 wire _01444_;
 wire _01445_;
 wire _01446_;
 wire _01447_;
 wire _01448_;
 wire _01449_;
 wire _01450_;
 wire _01451_;
 wire _01452_;
 wire _01453_;
 wire _01454_;
 wire _01455_;
 wire _01456_;
 wire _01457_;
 wire _01458_;
 wire _01459_;
 wire _01460_;
 wire _01461_;
 wire _01462_;
 wire _01463_;
 wire _01464_;
 wire _01465_;
 wire _01466_;
 wire _01467_;
 wire _01468_;
 wire _01469_;
 wire _01470_;
 wire _01471_;
 wire _01472_;
 wire _01473_;
 wire _01474_;
 wire _01475_;
 wire _01476_;
 wire _01477_;
 wire _01478_;
 wire _01479_;
 wire _01480_;
 wire _01481_;
 wire _01482_;
 wire _01483_;
 wire _01484_;
 wire _01485_;
 wire _01486_;
 wire _01487_;
 wire _01488_;
 wire _01489_;
 wire _01490_;
 wire _01491_;
 wire _01492_;
 wire _01493_;
 wire _01494_;
 wire _01495_;
 wire _01496_;
 wire _01497_;
 wire _01498_;
 wire _01499_;
 wire _01500_;
 wire _01501_;
 wire _01502_;
 wire _01503_;
 wire _01504_;
 wire _01505_;
 wire _01506_;
 wire _01507_;
 wire _01508_;
 wire _01509_;
 wire _01510_;
 wire _01511_;
 wire _01512_;
 wire _01513_;
 wire _01514_;
 wire _01515_;
 wire _01516_;
 wire _01517_;
 wire _01518_;
 wire _01519_;
 wire _01520_;
 wire _01521_;
 wire _01522_;
 wire _01523_;
 wire _01524_;
 wire _01525_;
 wire _01526_;
 wire _01527_;
 wire _01528_;
 wire _01529_;
 wire _01530_;
 wire _01531_;
 wire _01532_;
 wire _01533_;
 wire _01534_;
 wire _01535_;
 wire _01536_;
 wire _01537_;
 wire _01538_;
 wire _01539_;
 wire _01540_;
 wire _01541_;
 wire _01542_;
 wire _01543_;
 wire _01544_;
 wire _01545_;
 wire _01546_;
 wire _01547_;
 wire _01548_;
 wire _01549_;
 wire _01550_;
 wire _01551_;
 wire _01552_;
 wire _01553_;
 wire _01554_;
 wire _01555_;
 wire _01556_;
 wire _01557_;
 wire _01558_;
 wire _01559_;
 wire _01560_;
 wire _01561_;
 wire _01562_;
 wire _01563_;
 wire _01564_;
 wire _01565_;
 wire _01566_;
 wire _01567_;
 wire _01568_;
 wire _01569_;
 wire _01570_;
 wire _01571_;
 wire _01572_;
 wire _01573_;
 wire _01574_;
 wire _01575_;
 wire _01576_;
 wire _01577_;
 wire _01578_;
 wire _01579_;
 wire _01580_;
 wire _01581_;
 wire _01582_;
 wire _01583_;
 wire _01584_;
 wire _01585_;
 wire _01586_;
 wire _01587_;
 wire _01588_;
 wire _01589_;
 wire _01590_;
 wire _01591_;
 wire _01592_;
 wire _01593_;
 wire _01594_;
 wire _01595_;
 wire _01596_;
 wire _01597_;
 wire _01598_;
 wire _01599_;
 wire _01600_;
 wire _01601_;
 wire _01602_;
 wire _01603_;
 wire _01604_;
 wire _01605_;
 wire _01606_;
 wire _01607_;
 wire _01608_;
 wire _01609_;
 wire _01610_;
 wire _01611_;
 wire _01612_;
 wire _01613_;
 wire _01614_;
 wire _01615_;
 wire _01616_;
 wire _01617_;
 wire _01618_;
 wire _01619_;
 wire _01620_;
 wire _01621_;
 wire _01622_;
 wire _01623_;
 wire _01624_;
 wire _01625_;
 wire _01626_;
 wire _01627_;
 wire _01628_;
 wire _01629_;
 wire _01630_;
 wire _01631_;
 wire _01632_;
 wire _01633_;
 wire _01634_;
 wire _01635_;
 wire _01636_;
 wire _01637_;
 wire _01638_;
 wire _01639_;
 wire _01640_;
 wire _01641_;
 wire _01642_;
 wire _01643_;
 wire _01644_;
 wire _01645_;
 wire _01646_;
 wire _01647_;
 wire _01648_;
 wire _01649_;
 wire _01650_;
 wire _01651_;
 wire _01652_;
 wire _01653_;
 wire _01654_;
 wire _01655_;
 wire _01656_;
 wire _01657_;
 wire _01658_;
 wire _01659_;
 wire _01660_;
 wire _01661_;
 wire _01662_;
 wire _01663_;
 wire _01664_;
 wire _01665_;
 wire _01666_;
 wire _01667_;
 wire _01668_;
 wire _01669_;
 wire _01670_;
 wire _01671_;
 wire _01672_;
 wire _01673_;
 wire _01674_;
 wire _01675_;
 wire _01676_;
 wire _01677_;
 wire _01678_;
 wire _01679_;
 wire _01680_;
 wire _01681_;
 wire _01682_;
 wire _01683_;
 wire _01684_;
 wire _01685_;
 wire _01686_;
 wire _01687_;
 wire _01688_;
 wire _01689_;
 wire _01690_;
 wire _01691_;
 wire _01692_;
 wire _01693_;
 wire _01694_;
 wire _01695_;
 wire _01696_;
 wire _01697_;
 wire _01698_;
 wire _01699_;
 wire _01700_;
 wire _01701_;
 wire _01702_;
 wire _01703_;
 wire _01704_;
 wire _01705_;
 wire _01706_;
 wire _01707_;
 wire _01708_;
 wire _01709_;
 wire _01710_;
 wire _01711_;
 wire _01712_;
 wire _01713_;
 wire _01714_;
 wire _01715_;
 wire _01716_;
 wire _01717_;
 wire _01718_;
 wire _01719_;
 wire _01720_;
 wire _01721_;
 wire _01722_;
 wire _01723_;
 wire _01724_;
 wire _01725_;
 wire _01726_;
 wire _01727_;
 wire _01728_;
 wire _01729_;
 wire _01730_;
 wire _01731_;
 wire _01732_;
 wire _01733_;
 wire _01734_;
 wire _01735_;
 wire _01736_;
 wire _01737_;
 wire _01738_;
 wire _01739_;
 wire _01740_;
 wire _01741_;
 wire _01742_;
 wire _01743_;
 wire _01744_;
 wire _01745_;
 wire _01746_;
 wire _01747_;
 wire _01748_;
 wire _01749_;
 wire _01750_;
 wire _01751_;
 wire _01752_;
 wire _01753_;
 wire _01754_;
 wire _01755_;
 wire _01756_;
 wire _01757_;
 wire _01758_;
 wire _01759_;
 wire _01760_;
 wire _01761_;
 wire _01762_;
 wire _01763_;
 wire _01764_;
 wire _01765_;
 wire _01766_;
 wire _01767_;
 wire _01768_;
 wire _01769_;
 wire _01770_;
 wire _01771_;
 wire _01772_;
 wire _01773_;
 wire _01774_;
 wire _01775_;
 wire _01776_;
 wire _01777_;
 wire _01778_;
 wire _01779_;
 wire _01780_;
 wire _01781_;
 wire _01782_;
 wire _01783_;
 wire _01784_;
 wire _01785_;
 wire _01786_;
 wire _01787_;
 wire _01788_;
 wire _01789_;
 wire _01790_;
 wire _01791_;
 wire _01792_;
 wire _01793_;
 wire _01794_;
 wire _01795_;
 wire _01796_;
 wire _01797_;
 wire _01798_;
 wire _01799_;
 wire _01800_;
 wire _01801_;
 wire _01802_;
 wire _01803_;
 wire _01804_;
 wire _01805_;
 wire _01806_;
 wire _01807_;
 wire _01808_;
 wire _01809_;
 wire _01810_;
 wire _01811_;
 wire _01812_;
 wire _01813_;
 wire _01814_;
 wire _01815_;
 wire _01816_;
 wire _01817_;
 wire _01818_;
 wire _01819_;
 wire _01820_;
 wire _01821_;
 wire _01822_;
 wire _01823_;
 wire _01824_;
 wire _01825_;
 wire _01826_;
 wire _01827_;
 wire _01828_;
 wire _01829_;
 wire _01830_;
 wire _01831_;
 wire _01832_;
 wire _01833_;
 wire _01834_;
 wire _01835_;
 wire _01836_;
 wire _01837_;
 wire _01838_;
 wire _01839_;
 wire _01840_;
 wire _01841_;
 wire _01842_;
 wire _01843_;
 wire _01844_;
 wire _01845_;
 wire _01846_;
 wire _01847_;
 wire _01848_;
 wire _01849_;
 wire _01850_;
 wire _01851_;
 wire _01852_;
 wire _01853_;
 wire _01854_;
 wire _01855_;
 wire _01856_;
 wire _01857_;
 wire _01858_;
 wire _01859_;
 wire _01860_;
 wire _01861_;
 wire _01862_;
 wire _01863_;
 wire _01864_;
 wire _01865_;
 wire _01866_;
 wire _01867_;
 wire _01868_;
 wire _01869_;
 wire _01870_;
 wire _01871_;
 wire _01872_;
 wire _01873_;
 wire _01874_;
 wire _01875_;
 wire _01876_;
 wire _01877_;
 wire _01878_;
 wire _01879_;
 wire _01880_;
 wire _01881_;
 wire _01882_;
 wire _01883_;
 wire _01884_;
 wire _01885_;
 wire _01886_;
 wire _01887_;
 wire _01888_;
 wire _01889_;
 wire _01890_;
 wire _01891_;
 wire _01892_;
 wire _01893_;
 wire _01894_;
 wire _01895_;
 wire _01896_;
 wire _01897_;
 wire _01898_;
 wire _01899_;
 wire _01900_;
 wire _01901_;
 wire _01902_;
 wire _01903_;
 wire _01904_;
 wire _01905_;
 wire _01906_;
 wire _01907_;
 wire _01908_;
 wire _01909_;
 wire _01910_;
 wire _01911_;
 wire _01912_;
 wire _01913_;
 wire _01914_;
 wire _01915_;
 wire _01916_;
 wire _01917_;
 wire _01918_;
 wire _01919_;
 wire _01920_;
 wire _01921_;
 wire _01922_;
 wire _01923_;
 wire _01924_;
 wire _01925_;
 wire _01926_;
 wire _01927_;
 wire _01928_;
 wire _01929_;
 wire _01930_;
 wire _01931_;
 wire _01932_;
 wire _01933_;
 wire _01934_;
 wire _01935_;
 wire _01936_;
 wire _01937_;
 wire _01938_;
 wire _01939_;
 wire _01940_;
 wire _01941_;
 wire _01942_;
 wire _01943_;
 wire _01944_;
 wire _01945_;
 wire _01946_;
 wire _01947_;
 wire _01948_;
 wire _01949_;
 wire _01950_;
 wire _01951_;
 wire _01952_;
 wire _01953_;
 wire _01954_;
 wire _01955_;
 wire _01956_;
 wire _01957_;
 wire _01958_;
 wire _01959_;
 wire _01960_;
 wire _01961_;
 wire _01962_;
 wire _01963_;
 wire _01964_;
 wire _01965_;
 wire _01966_;
 wire _01967_;
 wire _01968_;
 wire _01969_;
 wire _01970_;
 wire _01971_;
 wire _01972_;
 wire _01973_;
 wire _01974_;
 wire _01975_;
 wire _01976_;
 wire _01977_;
 wire _01978_;
 wire _01979_;
 wire _01980_;
 wire _01981_;
 wire _01982_;
 wire _01983_;
 wire _01984_;
 wire _01985_;
 wire _01986_;
 wire _01987_;
 wire _01988_;
 wire _01989_;
 wire _01990_;
 wire _01991_;
 wire _01992_;
 wire _01993_;
 wire _01994_;
 wire _01995_;
 wire _01996_;
 wire _01997_;
 wire _01998_;
 wire _01999_;
 wire _02000_;
 wire _02001_;
 wire _02002_;
 wire _02003_;
 wire _02004_;
 wire _02005_;
 wire _02006_;
 wire _02007_;
 wire _02008_;
 wire _02009_;
 wire _02010_;
 wire _02011_;
 wire _02012_;
 wire _02013_;
 wire _02014_;
 wire _02015_;
 wire _02016_;
 wire _02017_;
 wire _02018_;
 wire _02019_;
 wire _02020_;
 wire _02021_;
 wire _02022_;
 wire _02023_;
 wire _02024_;
 wire _02025_;
 wire _02026_;
 wire _02027_;
 wire _02028_;
 wire _02029_;
 wire _02030_;
 wire _02031_;
 wire _02032_;
 wire _02033_;
 wire _02034_;
 wire _02035_;
 wire _02036_;
 wire _02037_;
 wire _02038_;
 wire _02039_;
 wire _02040_;
 wire _02041_;
 wire _02042_;
 wire _02043_;
 wire _02044_;
 wire _02045_;
 wire _02046_;
 wire _02047_;
 wire _02048_;
 wire _02049_;
 wire _02050_;
 wire _02051_;
 wire _02052_;
 wire _02053_;
 wire _02054_;
 wire _02055_;
 wire _02056_;
 wire _02057_;
 wire _02058_;
 wire _02059_;
 wire _02060_;
 wire _02061_;
 wire _02062_;
 wire _02063_;
 wire _02064_;
 wire _02065_;
 wire _02066_;
 wire _02067_;
 wire _02068_;
 wire _02069_;
 wire _02070_;
 wire _02071_;
 wire _02072_;
 wire _02073_;
 wire _02074_;
 wire _02075_;
 wire _02076_;
 wire _02077_;
 wire _02078_;
 wire _02079_;
 wire _02080_;
 wire _02081_;
 wire _02082_;
 wire _02083_;
 wire _02084_;
 wire _02085_;
 wire _02086_;
 wire _02087_;
 wire _02088_;
 wire _02089_;
 wire _02090_;
 wire _02091_;
 wire _02092_;
 wire _02093_;
 wire _02094_;
 wire _02095_;
 wire _02096_;
 wire _02097_;
 wire _02098_;
 wire _02099_;
 wire _02100_;
 wire _02101_;
 wire _02102_;
 wire _02103_;
 wire _02104_;
 wire _02105_;
 wire _02106_;
 wire _02107_;
 wire _02108_;
 wire _02109_;
 wire _02110_;
 wire _02111_;
 wire _02112_;
 wire _02113_;
 wire _02114_;
 wire _02115_;
 wire _02116_;
 wire _02117_;
 wire _02118_;
 wire _02119_;
 wire _02120_;
 wire _02121_;
 wire _02122_;
 wire _02123_;
 wire _02124_;
 wire _02125_;
 wire _02126_;
 wire _02127_;
 wire _02128_;
 wire _02129_;
 wire _02130_;
 wire _02131_;
 wire _02132_;
 wire _02133_;
 wire _02134_;
 wire _02135_;
 wire _02136_;
 wire _02137_;
 wire _02138_;
 wire _02139_;
 wire _02140_;
 wire _02141_;
 wire _02142_;
 wire _02143_;
 wire _02144_;
 wire _02145_;
 wire _02146_;
 wire _02147_;
 wire _02148_;
 wire _02149_;
 wire _02150_;
 wire _02151_;
 wire _02152_;
 wire _02153_;
 wire _02154_;
 wire _02155_;
 wire _02156_;
 wire _02157_;
 wire _02158_;
 wire _02159_;
 wire _02160_;
 wire _02161_;
 wire _02162_;
 wire _02163_;
 wire _02164_;
 wire _02165_;
 wire _02166_;
 wire _02167_;
 wire _02168_;
 wire _02169_;
 wire _02170_;
 wire _02171_;
 wire _02172_;
 wire _02173_;
 wire _02174_;
 wire _02175_;
 wire _02176_;
 wire _02177_;
 wire _02178_;
 wire _02179_;
 wire _02180_;
 wire _02181_;
 wire _02182_;
 wire _02183_;
 wire _02184_;
 wire _02185_;
 wire _02186_;
 wire _02187_;
 wire _02188_;
 wire _02189_;
 wire _02190_;
 wire _02191_;
 wire _02192_;
 wire _02193_;
 wire _02194_;
 wire _02195_;
 wire _02196_;
 wire _02197_;
 wire _02198_;
 wire _02199_;
 wire _02200_;
 wire _02201_;
 wire _02202_;
 wire _02203_;
 wire _02204_;
 wire _02205_;
 wire _02206_;
 wire _02207_;
 wire _02208_;
 wire _02209_;
 wire _02210_;
 wire _02211_;
 wire _02212_;
 wire _02213_;
 wire _02214_;
 wire _02215_;
 wire _02216_;
 wire _02217_;
 wire _02218_;
 wire _02219_;
 wire _02220_;
 wire _02221_;
 wire _02222_;
 wire _02223_;
 wire _02224_;
 wire _02225_;
 wire _02226_;
 wire _02227_;
 wire _02228_;
 wire _02229_;
 wire _02230_;
 wire _02231_;
 wire _02232_;
 wire _02233_;
 wire _02234_;
 wire _02235_;
 wire _02236_;
 wire _02237_;
 wire _02238_;
 wire _02239_;
 wire _02240_;
 wire _02241_;
 wire _02242_;
 wire _02243_;
 wire _02244_;
 wire _02245_;
 wire _02246_;
 wire _02247_;
 wire _02248_;
 wire _02249_;
 wire _02250_;
 wire _02251_;
 wire _02252_;
 wire _02253_;
 wire _02254_;
 wire _02255_;
 wire _02256_;
 wire _02257_;
 wire _02258_;
 wire _02259_;
 wire _02260_;
 wire _02261_;
 wire _02262_;
 wire _02263_;
 wire _02264_;
 wire _02265_;
 wire _02266_;
 wire _02267_;
 wire _02268_;
 wire _02269_;
 wire _02270_;
 wire _02271_;
 wire _02272_;
 wire _02273_;
 wire _02274_;
 wire _02275_;
 wire _02276_;
 wire _02277_;
 wire _02278_;
 wire _02279_;
 wire _02280_;
 wire _02281_;
 wire _02282_;
 wire _02283_;
 wire _02284_;
 wire _02285_;
 wire _02286_;
 wire _02287_;
 wire _02288_;
 wire _02289_;
 wire _02290_;
 wire _02291_;
 wire _02292_;
 wire _02293_;
 wire _02294_;
 wire _02295_;
 wire _02296_;
 wire _02297_;
 wire _02298_;
 wire _02299_;
 wire _02300_;
 wire _02301_;
 wire _02302_;
 wire _02303_;
 wire _02304_;
 wire _02305_;
 wire _02306_;
 wire _02307_;
 wire _02308_;
 wire _02309_;
 wire _02310_;
 wire _02311_;
 wire _02312_;
 wire _02313_;
 wire _02314_;
 wire _02315_;
 wire _02316_;
 wire _02317_;
 wire _02318_;
 wire _02319_;
 wire _02320_;
 wire _02321_;
 wire _02322_;
 wire _02323_;
 wire _02324_;
 wire _02325_;
 wire _02326_;
 wire _02327_;
 wire _02328_;
 wire _02329_;
 wire _02330_;
 wire _02331_;
 wire _02332_;
 wire _02333_;
 wire _02334_;
 wire _02335_;
 wire _02336_;
 wire _02337_;
 wire _02338_;
 wire _02339_;
 wire _02340_;
 wire _02341_;
 wire _02342_;
 wire _02343_;
 wire _02344_;
 wire _02345_;
 wire _02346_;
 wire _02347_;
 wire _02348_;
 wire _02349_;
 wire _02350_;
 wire _02351_;
 wire _02352_;
 wire _02353_;
 wire _02354_;
 wire _02355_;
 wire _02356_;
 wire _02357_;
 wire _02358_;
 wire _02359_;
 wire _02360_;
 wire _02361_;
 wire _02362_;
 wire _02363_;
 wire _02364_;
 wire _02365_;
 wire _02366_;
 wire _02367_;
 wire _02368_;
 wire _02369_;
 wire _02370_;
 wire _02371_;
 wire _02372_;
 wire _02373_;
 wire _02374_;
 wire _02375_;
 wire _02376_;
 wire _02377_;
 wire _02378_;
 wire _02379_;
 wire _02380_;
 wire _02381_;
 wire _02382_;
 wire _02383_;
 wire _02384_;
 wire _02385_;
 wire _02386_;
 wire _02387_;
 wire _02388_;
 wire _02389_;
 wire _02390_;
 wire _02391_;
 wire _02392_;
 wire _02393_;
 wire _02394_;
 wire _02395_;
 wire _02396_;
 wire _02397_;
 wire _02398_;
 wire _02399_;
 wire _02400_;
 wire _02401_;
 wire _02402_;
 wire _02403_;
 wire _02404_;
 wire _02405_;
 wire _02406_;
 wire _02407_;
 wire _02408_;
 wire _02409_;
 wire _02410_;
 wire _02411_;
 wire _02412_;
 wire _02413_;
 wire _02414_;
 wire _02415_;
 wire _02416_;
 wire _02417_;
 wire _02418_;
 wire _02419_;
 wire _02420_;
 wire _02421_;
 wire _02422_;
 wire _02423_;
 wire _02424_;
 wire _02425_;
 wire _02426_;
 wire _02427_;
 wire _02428_;
 wire _02429_;
 wire _02430_;
 wire _02431_;
 wire _02432_;
 wire _02433_;
 wire _02434_;
 wire _02435_;
 wire _02436_;
 wire _02437_;
 wire _02438_;
 wire _02439_;
 wire _02440_;
 wire _02441_;
 wire _02442_;
 wire _02443_;
 wire _02444_;
 wire _02445_;
 wire _02446_;
 wire _02447_;
 wire _02448_;
 wire _02449_;
 wire _02450_;
 wire _02451_;
 wire _02452_;
 wire _02453_;
 wire _02454_;
 wire _02455_;
 wire _02456_;
 wire _02457_;
 wire _02458_;
 wire _02459_;
 wire _02460_;
 wire _02461_;
 wire _02462_;
 wire _02463_;
 wire _02464_;
 wire _02465_;
 wire _02466_;
 wire _02467_;
 wire _02468_;
 wire _02469_;
 wire _02470_;
 wire _02471_;
 wire _02472_;
 wire _02473_;
 wire _02474_;
 wire _02475_;
 wire _02476_;
 wire _02477_;
 wire _02478_;
 wire _02479_;
 wire _02480_;
 wire _02481_;
 wire _02482_;
 wire _02483_;
 wire _02484_;
 wire _02485_;
 wire _02486_;
 wire _02487_;
 wire _02488_;
 wire _02489_;
 wire _02490_;
 wire _02491_;
 wire _02492_;
 wire _02493_;
 wire _02494_;
 wire _02495_;
 wire _02496_;
 wire _02497_;
 wire _02498_;
 wire _02499_;
 wire _02500_;
 wire _02501_;
 wire _02502_;
 wire _02503_;
 wire _02504_;
 wire _02505_;
 wire _02506_;
 wire _02507_;
 wire _02508_;
 wire _02509_;
 wire _02510_;
 wire _02511_;
 wire _02512_;
 wire _02513_;
 wire _02514_;
 wire _02515_;
 wire _02516_;
 wire _02517_;
 wire _02518_;
 wire _02519_;
 wire _02520_;
 wire _02521_;
 wire _02522_;
 wire _02523_;
 wire _02524_;
 wire _02525_;
 wire _02526_;
 wire _02527_;
 wire _02528_;
 wire _02529_;
 wire _02530_;
 wire _02531_;
 wire _02532_;
 wire _02533_;
 wire _02534_;
 wire _02535_;
 wire _02536_;
 wire _02537_;
 wire _02538_;
 wire _02539_;
 wire _02540_;
 wire _02541_;
 wire _02542_;
 wire _02543_;
 wire _02544_;
 wire _02545_;
 wire _02546_;
 wire _02547_;
 wire _02548_;
 wire _02549_;
 wire _02550_;
 wire _02551_;
 wire _02552_;
 wire _02553_;
 wire _02554_;
 wire _02555_;
 wire _02556_;
 wire _02557_;
 wire _02558_;
 wire _02559_;
 wire _02560_;
 wire _02561_;
 wire _02562_;
 wire _02563_;
 wire _02564_;
 wire _02565_;
 wire _02566_;
 wire _02567_;
 wire _02568_;
 wire _02569_;
 wire _02570_;
 wire _02571_;
 wire _02572_;
 wire _02573_;
 wire _02574_;
 wire _02575_;
 wire _02576_;
 wire _02577_;
 wire _02578_;
 wire _02579_;
 wire _02580_;
 wire _02581_;
 wire _02582_;
 wire _02583_;
 wire _02584_;
 wire _02585_;
 wire _02586_;
 wire _02587_;
 wire _02588_;
 wire _02589_;
 wire _02590_;
 wire _02591_;
 wire _02592_;
 wire _02593_;
 wire _02594_;
 wire _02595_;
 wire _02596_;
 wire _02597_;
 wire _02598_;
 wire _02599_;
 wire _02600_;
 wire _02601_;
 wire _02602_;
 wire _02603_;
 wire _02604_;
 wire _02605_;
 wire _02606_;
 wire _02607_;
 wire _02608_;
 wire _02609_;
 wire _02610_;
 wire _02611_;
 wire _02612_;
 wire _02613_;
 wire _02614_;
 wire _02615_;
 wire _02616_;
 wire _02617_;
 wire _02618_;
 wire _02619_;
 wire _02620_;
 wire _02621_;
 wire _02622_;
 wire _02623_;
 wire _02624_;
 wire _02625_;
 wire _02626_;
 wire _02627_;
 wire _02628_;
 wire _02629_;
 wire _02630_;
 wire _02631_;
 wire _02632_;
 wire _02633_;
 wire _02634_;
 wire _02635_;
 wire _02636_;
 wire _02637_;
 wire _02638_;
 wire _02639_;
 wire _02640_;
 wire _02641_;
 wire _02642_;
 wire _02643_;
 wire _02644_;
 wire _02645_;
 wire _02646_;
 wire _02647_;
 wire _02648_;
 wire _02649_;
 wire _02650_;
 wire _02651_;
 wire _02652_;
 wire _02653_;
 wire _02654_;
 wire _02655_;
 wire _02656_;
 wire _02657_;
 wire _02658_;
 wire _02659_;
 wire _02660_;
 wire _02661_;
 wire _02662_;
 wire _02663_;
 wire _02664_;
 wire _02665_;
 wire _02666_;
 wire _02667_;
 wire _02668_;
 wire _02669_;
 wire _02670_;
 wire _02671_;
 wire _02672_;
 wire _02673_;
 wire _02674_;
 wire _02675_;
 wire _02676_;
 wire _02677_;
 wire _02678_;
 wire _02679_;
 wire _02680_;
 wire _02681_;
 wire _02682_;
 wire _02683_;
 wire _02684_;
 wire _02685_;
 wire _02686_;
 wire _02687_;
 wire _02688_;
 wire _02689_;
 wire _02690_;
 wire _02691_;
 wire _02692_;
 wire _02693_;
 wire _02694_;
 wire _02695_;
 wire _02696_;
 wire _02697_;
 wire _02698_;
 wire _02699_;
 wire _02700_;
 wire _02701_;
 wire _02702_;
 wire _02703_;
 wire _02704_;
 wire _02705_;
 wire _02706_;
 wire _02707_;
 wire _02708_;
 wire _02709_;
 wire _02710_;
 wire _02711_;
 wire _02712_;
 wire _02713_;
 wire _02714_;
 wire _02715_;
 wire _02716_;
 wire _02717_;
 wire _02718_;
 wire _02719_;
 wire _02720_;
 wire _02721_;
 wire _02722_;
 wire _02723_;
 wire _02724_;
 wire _02725_;
 wire _02726_;
 wire _02727_;
 wire _02728_;
 wire _02729_;
 wire _02730_;
 wire _02731_;
 wire _02732_;
 wire _02733_;
 wire _02734_;
 wire _02735_;
 wire _02736_;
 wire _02737_;
 wire _02738_;
 wire _02739_;
 wire _02740_;
 wire _02741_;
 wire _02742_;
 wire _02743_;
 wire _02744_;
 wire _02745_;
 wire _02746_;
 wire _02747_;
 wire _02748_;
 wire _02749_;
 wire _02750_;
 wire _02751_;
 wire _02752_;
 wire _02753_;
 wire _02754_;
 wire _02755_;
 wire _02756_;
 wire _02757_;
 wire _02758_;
 wire _02759_;
 wire _02760_;
 wire _02761_;
 wire _02762_;
 wire _02763_;
 wire _02764_;
 wire _02765_;
 wire _02766_;
 wire _02767_;
 wire _02768_;
 wire _02769_;
 wire _02770_;
 wire _02771_;
 wire _02772_;
 wire _02773_;
 wire _02774_;
 wire _02775_;
 wire _02776_;
 wire _02777_;
 wire _02778_;
 wire _02779_;
 wire _02780_;
 wire _02781_;
 wire _02782_;
 wire _02783_;
 wire _02784_;
 wire _02785_;
 wire _02786_;
 wire _02787_;
 wire _02788_;
 wire _02789_;
 wire _02790_;
 wire _02791_;
 wire _02792_;
 wire _02793_;
 wire _02794_;
 wire _02795_;
 wire _02796_;
 wire _02797_;
 wire _02798_;
 wire _02799_;
 wire _02800_;
 wire _02801_;
 wire _02802_;
 wire _02803_;
 wire _02804_;
 wire _02805_;
 wire _02806_;
 wire _02807_;
 wire _02808_;
 wire _02809_;
 wire _02810_;
 wire _02811_;
 wire _02812_;
 wire _02813_;
 wire _02814_;
 wire _02815_;
 wire _02816_;
 wire _02817_;
 wire _02818_;
 wire _02819_;
 wire _02820_;
 wire _02821_;
 wire _02822_;
 wire _02823_;
 wire _02824_;
 wire _02825_;
 wire _02826_;
 wire _02827_;
 wire _02828_;
 wire _02829_;
 wire _02830_;
 wire _02831_;
 wire _02832_;
 wire _02833_;
 wire _02834_;
 wire _02835_;
 wire _02836_;
 wire _02837_;
 wire _02838_;
 wire _02839_;
 wire _02840_;
 wire _02841_;
 wire _02842_;
 wire _02843_;
 wire _02844_;
 wire _02845_;
 wire _02846_;
 wire _02847_;
 wire _02848_;
 wire _02849_;
 wire _02850_;
 wire _02851_;
 wire _02852_;
 wire _02853_;
 wire _02854_;
 wire _02855_;
 wire _02856_;
 wire _02857_;
 wire _02858_;
 wire _02859_;
 wire _02860_;
 wire _02861_;
 wire _02862_;
 wire _02863_;
 wire _02864_;
 wire _02865_;
 wire _02866_;
 wire _02867_;
 wire _02868_;
 wire _02869_;
 wire _02870_;
 wire _02871_;
 wire _02872_;
 wire _02873_;
 wire _02874_;
 wire _02875_;
 wire _02876_;
 wire _02877_;
 wire _02878_;
 wire _02879_;
 wire _02880_;
 wire _02881_;
 wire _02882_;
 wire _02883_;
 wire _02884_;
 wire _02885_;
 wire _02886_;
 wire _02887_;
 wire _02888_;
 wire _02889_;
 wire _02890_;
 wire _02891_;
 wire _02892_;
 wire _02893_;
 wire _02894_;
 wire _02895_;
 wire _02896_;
 wire _02897_;
 wire _02898_;
 wire _02899_;
 wire _02900_;
 wire _02901_;
 wire _02902_;
 wire _02903_;
 wire _02904_;
 wire _02905_;
 wire _02906_;
 wire _02907_;
 wire _02908_;
 wire _02909_;
 wire _02910_;
 wire _02911_;
 wire _02912_;
 wire _02913_;
 wire _02914_;
 wire _02915_;
 wire _02916_;
 wire _02917_;
 wire _02918_;
 wire _02919_;
 wire _02920_;
 wire _02921_;
 wire _02922_;
 wire _02923_;
 wire _02924_;
 wire _02925_;
 wire _02926_;
 wire _02927_;
 wire _02928_;
 wire _02929_;
 wire _02930_;
 wire _02931_;
 wire _02932_;
 wire _02933_;
 wire _02934_;
 wire _02935_;
 wire _02936_;
 wire _02937_;
 wire _02938_;
 wire _02939_;
 wire _02940_;
 wire _02941_;
 wire _02942_;
 wire _02943_;
 wire _02944_;
 wire _02945_;
 wire _02946_;
 wire _02947_;
 wire _02948_;
 wire _02949_;
 wire _02950_;
 wire _02951_;
 wire _02952_;
 wire _02953_;
 wire _02954_;
 wire _02955_;
 wire _02956_;
 wire _02957_;
 wire _02958_;
 wire _02959_;
 wire _02960_;
 wire _02961_;
 wire _02962_;
 wire _02963_;
 wire _02964_;
 wire _02965_;
 wire _02966_;
 wire _02967_;
 wire _02968_;
 wire _02969_;
 wire _02970_;
 wire _02971_;
 wire _02972_;
 wire _02973_;
 wire _02974_;
 wire _02975_;
 wire _02976_;
 wire _02977_;
 wire _02978_;
 wire _02979_;
 wire _02980_;
 wire _02981_;
 wire _02982_;
 wire _02983_;
 wire _02984_;
 wire _02985_;
 wire _02986_;
 wire _02987_;
 wire _02988_;
 wire _02989_;
 wire _02990_;
 wire _02991_;
 wire _02992_;
 wire _02993_;
 wire _02994_;
 wire _02995_;
 wire _02996_;
 wire _02997_;
 wire _02998_;
 wire _02999_;
 wire _03000_;
 wire _03001_;
 wire _03002_;
 wire _03003_;
 wire _03004_;
 wire _03005_;
 wire _03006_;
 wire _03007_;
 wire _03008_;
 wire _03009_;
 wire _03010_;
 wire _03011_;
 wire _03012_;
 wire _03013_;
 wire _03014_;
 wire _03015_;
 wire _03016_;
 wire _03017_;
 wire _03018_;
 wire _03019_;
 wire _03020_;
 wire _03021_;
 wire _03022_;
 wire _03023_;
 wire _03024_;
 wire _03025_;
 wire _03026_;
 wire _03027_;
 wire _03028_;
 wire _03029_;
 wire _03030_;
 wire _03031_;
 wire _03032_;
 wire _03033_;
 wire _03034_;
 wire _03035_;
 wire _03036_;
 wire _03037_;
 wire _03038_;
 wire _03039_;
 wire _03040_;
 wire _03041_;
 wire _03042_;
 wire _03043_;
 wire _03044_;
 wire _03045_;
 wire _03046_;
 wire _03047_;
 wire _03048_;
 wire _03049_;
 wire _03050_;
 wire _03051_;
 wire _03052_;
 wire _03053_;
 wire _03054_;
 wire _03055_;
 wire _03056_;
 wire _03057_;
 wire _03058_;
 wire _03059_;
 wire _03060_;
 wire _03061_;
 wire _03062_;
 wire _03063_;
 wire _03064_;
 wire _03065_;
 wire _03066_;
 wire _03067_;
 wire _03068_;
 wire _03069_;
 wire _03070_;
 wire _03071_;
 wire _03072_;
 wire _03073_;
 wire _03074_;
 wire _03075_;
 wire _03076_;
 wire _03077_;
 wire _03078_;
 wire _03079_;
 wire _03080_;
 wire _03081_;
 wire _03082_;
 wire _03083_;
 wire _03084_;
 wire _03085_;
 wire _03086_;
 wire _03087_;
 wire _03088_;
 wire _03089_;
 wire _03090_;
 wire _03091_;
 wire _03092_;
 wire _03093_;
 wire _03094_;
 wire _03095_;
 wire _03096_;
 wire _03097_;
 wire _03098_;
 wire _03099_;
 wire _03100_;
 wire _03101_;
 wire _03102_;
 wire _03103_;
 wire _03104_;
 wire _03105_;
 wire _03106_;
 wire _03107_;
 wire _03108_;
 wire _03109_;
 wire _03110_;
 wire _03111_;
 wire _03112_;
 wire _03113_;
 wire _03114_;
 wire _03115_;
 wire _03116_;
 wire _03117_;
 wire _03118_;
 wire _03119_;
 wire _03120_;
 wire _03121_;
 wire _03122_;
 wire _03123_;
 wire _03124_;
 wire _03125_;
 wire _03126_;
 wire _03127_;
 wire _03128_;
 wire _03129_;
 wire _03130_;
 wire _03131_;
 wire _03132_;
 wire _03133_;
 wire _03134_;
 wire _03135_;
 wire _03136_;
 wire _03137_;
 wire _03138_;
 wire _03139_;
 wire _03140_;
 wire _03141_;
 wire _03142_;
 wire _03143_;
 wire _03144_;
 wire _03145_;
 wire _03146_;
 wire _03147_;
 wire _03148_;
 wire _03149_;
 wire _03150_;
 wire _03151_;
 wire _03152_;
 wire _03153_;
 wire _03154_;
 wire _03155_;
 wire _03156_;
 wire _03157_;
 wire _03158_;
 wire _03159_;
 wire _03160_;
 wire _03161_;
 wire _03162_;
 wire _03163_;
 wire _03164_;
 wire _03165_;
 wire _03166_;
 wire _03167_;
 wire _03168_;
 wire _03169_;
 wire _03170_;
 wire _03171_;
 wire _03172_;
 wire _03173_;
 wire _03174_;
 wire _03175_;
 wire _03176_;
 wire _03177_;
 wire _03178_;
 wire _03179_;
 wire _03180_;
 wire _03181_;
 wire _03182_;
 wire _03183_;
 wire _03184_;
 wire _03185_;
 wire _03186_;
 wire _03187_;
 wire _03188_;
 wire _03189_;
 wire _03190_;
 wire _03191_;
 wire _03192_;
 wire _03193_;
 wire _03194_;
 wire _03195_;
 wire _03196_;
 wire _03197_;
 wire _03198_;
 wire _03199_;
 wire _03200_;
 wire _03201_;
 wire _03202_;
 wire _03203_;
 wire _03204_;
 wire _03205_;
 wire _03206_;
 wire _03207_;
 wire _03208_;
 wire _03209_;
 wire _03210_;
 wire _03211_;
 wire _03212_;
 wire _03213_;
 wire _03214_;
 wire _03215_;
 wire _03216_;
 wire _03217_;
 wire _03218_;
 wire _03219_;
 wire _03220_;
 wire _03221_;
 wire _03222_;
 wire _03223_;
 wire _03224_;
 wire _03225_;
 wire _03226_;
 wire _03227_;
 wire _03228_;
 wire _03229_;
 wire _03230_;
 wire _03231_;
 wire _03232_;
 wire _03233_;
 wire _03234_;
 wire _03235_;
 wire _03236_;
 wire _03237_;
 wire _03238_;
 wire _03239_;
 wire _03240_;
 wire _03241_;
 wire _03242_;
 wire _03243_;
 wire _03244_;
 wire _03245_;
 wire _03246_;
 wire _03247_;
 wire _03248_;
 wire _03249_;
 wire _03250_;
 wire _03251_;
 wire _03252_;
 wire _03253_;
 wire _03254_;
 wire _03255_;
 wire _03256_;
 wire _03257_;
 wire _03258_;
 wire _03259_;
 wire _03260_;
 wire _03261_;
 wire _03262_;
 wire _03263_;
 wire _03264_;
 wire _03265_;
 wire _03266_;
 wire _03267_;
 wire _03268_;
 wire _03269_;
 wire _03270_;
 wire _03271_;
 wire _03272_;
 wire _03273_;
 wire _03274_;
 wire _03275_;
 wire _03276_;
 wire _03277_;
 wire _03278_;
 wire _03279_;
 wire _03280_;
 wire _03281_;
 wire _03282_;
 wire _03283_;
 wire _03284_;
 wire _03285_;
 wire _03286_;
 wire _03287_;
 wire _03288_;
 wire _03289_;
 wire _03290_;
 wire _03291_;
 wire _03292_;
 wire _03293_;
 wire _03294_;
 wire _03295_;
 wire _03296_;
 wire _03297_;
 wire _03298_;
 wire _03299_;
 wire _03300_;
 wire _03301_;
 wire _03302_;
 wire _03303_;
 wire _03304_;
 wire _03305_;
 wire _03306_;
 wire _03307_;
 wire _03308_;
 wire _03309_;
 wire _03310_;
 wire _03311_;
 wire _03312_;
 wire _03313_;
 wire _03314_;
 wire _03315_;
 wire _03316_;
 wire _03317_;
 wire _03318_;
 wire _03319_;
 wire _03320_;
 wire _03321_;
 wire _03322_;
 wire _03323_;
 wire _03324_;
 wire _03325_;
 wire _03326_;
 wire _03327_;
 wire _03328_;
 wire _03329_;
 wire _03330_;
 wire _03331_;
 wire _03332_;
 wire _03333_;
 wire _03334_;
 wire _03335_;
 wire _03336_;
 wire _03337_;
 wire _03338_;
 wire _03339_;
 wire _03340_;
 wire _03341_;
 wire _03342_;
 wire _03343_;
 wire _03344_;
 wire _03345_;
 wire _03346_;
 wire _03347_;
 wire _03348_;
 wire _03349_;
 wire _03350_;
 wire _03351_;
 wire _03352_;
 wire _03353_;
 wire _03354_;
 wire _03355_;
 wire _03356_;
 wire _03357_;
 wire _03358_;
 wire _03359_;
 wire _03360_;
 wire _03361_;
 wire _03362_;
 wire _03363_;
 wire _03364_;
 wire _03365_;
 wire _03366_;
 wire _03367_;
 wire _03368_;
 wire _03369_;
 wire _03370_;
 wire _03371_;
 wire _03372_;
 wire _03373_;
 wire _03374_;
 wire _03375_;
 wire _03376_;
 wire _03377_;
 wire _03378_;
 wire _03379_;
 wire _03380_;
 wire _03381_;
 wire _03382_;
 wire _03383_;
 wire _03384_;
 wire _03385_;
 wire _03386_;
 wire _03387_;
 wire _03388_;
 wire _03389_;
 wire _03390_;
 wire _03391_;
 wire _03392_;
 wire _03393_;
 wire _03394_;
 wire _03395_;
 wire _03396_;
 wire _03397_;
 wire _03398_;
 wire _03399_;
 wire _03400_;
 wire _03401_;
 wire _03402_;
 wire _03403_;
 wire _03404_;
 wire _03405_;
 wire _03406_;
 wire _03407_;
 wire _03408_;
 wire _03409_;
 wire _03410_;
 wire _03411_;
 wire _03412_;
 wire _03413_;
 wire _03414_;
 wire _03415_;
 wire _03416_;
 wire _03417_;
 wire _03418_;
 wire _03419_;
 wire _03420_;
 wire _03421_;
 wire _03422_;
 wire _03423_;
 wire _03424_;
 wire _03425_;
 wire _03426_;
 wire _03427_;
 wire _03428_;
 wire _03429_;
 wire _03430_;
 wire _03431_;
 wire _03432_;
 wire _03433_;
 wire _03434_;
 wire _03435_;
 wire _03436_;
 wire _03437_;
 wire _03438_;
 wire _03439_;
 wire _03440_;
 wire _03441_;
 wire _03442_;
 wire _03443_;
 wire _03444_;
 wire _03445_;
 wire _03446_;
 wire _03447_;
 wire _03448_;
 wire _03449_;
 wire _03450_;
 wire _03451_;
 wire _03452_;
 wire _03453_;
 wire _03454_;
 wire _03455_;
 wire _03456_;
 wire _03457_;
 wire _03458_;
 wire _03459_;
 wire _03460_;
 wire _03461_;
 wire _03462_;
 wire _03463_;
 wire _03464_;
 wire _03465_;
 wire _03466_;
 wire _03467_;
 wire _03468_;
 wire _03469_;
 wire _03470_;
 wire _03471_;
 wire _03472_;
 wire _03473_;
 wire _03474_;
 wire _03475_;
 wire _03476_;
 wire _03477_;
 wire _03478_;
 wire _03479_;
 wire _03480_;
 wire _03481_;
 wire _03482_;
 wire _03483_;
 wire _03484_;
 wire _03485_;
 wire _03486_;
 wire _03487_;
 wire _03488_;
 wire _03489_;
 wire _03490_;
 wire _03491_;
 wire _03492_;
 wire _03493_;
 wire _03494_;
 wire _03495_;
 wire _03496_;
 wire _03497_;
 wire _03498_;
 wire _03499_;
 wire _03500_;
 wire _03501_;
 wire _03502_;
 wire _03503_;
 wire _03504_;
 wire _03505_;
 wire _03506_;
 wire _03507_;
 wire _03508_;
 wire _03509_;
 wire _03510_;
 wire _03511_;
 wire _03512_;
 wire _03513_;
 wire _03514_;
 wire _03515_;
 wire _03516_;
 wire _03517_;
 wire _03518_;
 wire _03519_;
 wire _03520_;
 wire _03521_;
 wire _03522_;
 wire _03523_;
 wire _03524_;
 wire _03525_;
 wire _03526_;
 wire _03527_;
 wire _03528_;
 wire _03529_;
 wire _03530_;
 wire _03531_;
 wire _03532_;
 wire _03533_;
 wire _03534_;
 wire _03535_;
 wire _03536_;
 wire _03537_;
 wire _03538_;
 wire _03539_;
 wire _03540_;
 wire _03541_;
 wire _03542_;
 wire _03543_;
 wire _03544_;
 wire _03545_;
 wire _03546_;
 wire _03547_;
 wire _03548_;
 wire _03549_;
 wire _03550_;
 wire _03551_;
 wire _03552_;
 wire _03553_;
 wire _03554_;
 wire _03555_;
 wire _03556_;
 wire _03557_;
 wire _03558_;
 wire _03559_;
 wire _03560_;
 wire _03561_;
 wire _03562_;
 wire _03563_;
 wire _03564_;
 wire _03565_;
 wire _03566_;
 wire _03567_;
 wire _03568_;
 wire _03569_;
 wire _03570_;
 wire _03571_;
 wire _03572_;
 wire _03573_;
 wire _03574_;
 wire _03575_;
 wire _03576_;
 wire _03577_;
 wire _03578_;
 wire _03579_;
 wire _03580_;
 wire _03581_;
 wire _03582_;
 wire _03583_;
 wire _03584_;
 wire _03585_;
 wire _03586_;
 wire _03587_;
 wire _03588_;
 wire _03589_;
 wire _03590_;
 wire _03591_;
 wire _03592_;
 wire _03593_;
 wire _03594_;
 wire _03595_;
 wire _03596_;
 wire _03597_;
 wire _03598_;
 wire _03599_;
 wire _03600_;
 wire _03601_;
 wire _03602_;
 wire _03603_;
 wire _03604_;
 wire _03605_;
 wire _03606_;
 wire _03607_;
 wire _03608_;
 wire _03609_;
 wire _03610_;
 wire _03611_;
 wire _03612_;
 wire _03613_;
 wire _03614_;
 wire _03615_;
 wire _03616_;
 wire _03617_;
 wire _03618_;
 wire _03619_;
 wire _03620_;
 wire _03621_;
 wire _03622_;
 wire _03623_;
 wire _03624_;
 wire _03625_;
 wire _03626_;
 wire _03627_;
 wire _03628_;
 wire _03629_;
 wire _03630_;
 wire _03631_;
 wire _03632_;
 wire _03633_;
 wire _03634_;
 wire _03635_;
 wire _03636_;
 wire _03637_;
 wire _03638_;
 wire _03639_;
 wire _03640_;
 wire _03641_;
 wire _03642_;
 wire _03643_;
 wire _03644_;
 wire _03645_;
 wire _03646_;
 wire _03647_;
 wire _03648_;
 wire _03649_;
 wire _03650_;
 wire _03651_;
 wire _03652_;
 wire _03653_;
 wire _03654_;
 wire _03655_;
 wire _03656_;
 wire _03657_;
 wire _03658_;
 wire _03659_;
 wire _03660_;
 wire _03661_;
 wire _03662_;
 wire _03663_;
 wire _03664_;
 wire _03665_;
 wire _03666_;
 wire _03667_;
 wire _03668_;
 wire _03669_;
 wire _03670_;
 wire _03671_;
 wire _03672_;
 wire _03673_;
 wire _03674_;
 wire _03675_;
 wire _03676_;
 wire _03677_;
 wire _03678_;
 wire _03679_;
 wire _03680_;
 wire _03681_;
 wire _03682_;
 wire _03683_;
 wire _03684_;
 wire _03685_;
 wire _03686_;
 wire _03687_;
 wire _03688_;
 wire _03689_;
 wire _03690_;
 wire _03691_;
 wire _03692_;
 wire _03693_;
 wire _03694_;
 wire _03695_;
 wire _03696_;
 wire _03697_;
 wire _03698_;
 wire _03699_;
 wire _03700_;
 wire _03701_;
 wire _03702_;
 wire _03703_;
 wire _03704_;
 wire _03705_;
 wire _03706_;
 wire _03707_;
 wire _03708_;
 wire _03709_;
 wire _03710_;
 wire _03711_;
 wire _03712_;
 wire _03713_;
 wire _03714_;
 wire _03715_;
 wire _03716_;
 wire _03717_;
 wire _03718_;
 wire _03719_;
 wire _03720_;
 wire _03721_;
 wire _03722_;
 wire _03723_;
 wire _03724_;
 wire _03725_;
 wire _03726_;
 wire _03727_;
 wire _03728_;
 wire _03729_;
 wire _03730_;
 wire _03731_;
 wire _03732_;
 wire _03733_;
 wire _03734_;
 wire _03735_;
 wire _03736_;
 wire _03737_;
 wire _03738_;
 wire _03739_;
 wire _03740_;
 wire _03741_;
 wire _03742_;
 wire _03743_;
 wire _03744_;
 wire _03745_;
 wire _03746_;
 wire _03747_;
 wire _03748_;
 wire _03749_;
 wire _03750_;
 wire _03751_;
 wire _03752_;
 wire _03753_;
 wire _03754_;
 wire _03755_;
 wire _03756_;
 wire _03757_;
 wire _03758_;
 wire _03759_;
 wire _03760_;
 wire _03761_;
 wire _03762_;
 wire _03763_;
 wire _03764_;
 wire _03765_;
 wire _03766_;
 wire _03767_;
 wire _03768_;
 wire _03769_;
 wire _03770_;
 wire _03771_;
 wire _03772_;
 wire _03773_;
 wire _03774_;
 wire _03775_;
 wire _03776_;
 wire _03777_;
 wire _03778_;
 wire _03779_;
 wire _03780_;
 wire _03781_;
 wire _03782_;
 wire _03783_;
 wire _03784_;
 wire _03785_;
 wire _03786_;
 wire _03787_;
 wire _03788_;
 wire _03789_;
 wire _03790_;
 wire _03791_;
 wire _03792_;
 wire _03793_;
 wire _03794_;
 wire _03795_;
 wire _03796_;
 wire _03797_;
 wire _03798_;
 wire _03799_;
 wire _03800_;
 wire _03801_;
 wire _03802_;
 wire _03803_;
 wire _03804_;
 wire _03805_;
 wire _03806_;
 wire _03807_;
 wire _03808_;
 wire _03809_;
 wire _03810_;
 wire _03811_;
 wire _03812_;
 wire _03813_;
 wire _03814_;
 wire _03815_;
 wire _03816_;
 wire _03817_;
 wire _03818_;
 wire _03819_;
 wire _03820_;
 wire _03821_;
 wire _03822_;
 wire _03823_;
 wire _03824_;
 wire _03825_;
 wire _03826_;
 wire _03827_;
 wire _03828_;
 wire _03829_;
 wire _03830_;
 wire _03831_;
 wire _03832_;
 wire _03833_;
 wire _03834_;
 wire _03835_;
 wire _03836_;
 wire _03837_;
 wire _03838_;
 wire _03839_;
 wire _03840_;
 wire _03841_;
 wire _03842_;
 wire _03843_;
 wire _03844_;
 wire _03845_;
 wire _03846_;
 wire _03847_;
 wire _03848_;
 wire _03849_;
 wire _03850_;
 wire _03851_;
 wire _03852_;
 wire _03853_;
 wire _03854_;
 wire _03855_;
 wire _03856_;
 wire _03857_;
 wire _03858_;
 wire _03859_;
 wire _03860_;
 wire _03861_;
 wire _03862_;
 wire _03863_;
 wire _03864_;
 wire _03865_;
 wire _03866_;
 wire _03867_;
 wire _03868_;
 wire _03869_;
 wire _03870_;
 wire _03871_;
 wire _03872_;
 wire _03873_;
 wire _03874_;
 wire _03875_;
 wire _03876_;
 wire _03877_;
 wire _03878_;
 wire _03879_;
 wire _03880_;
 wire _03881_;
 wire _03882_;
 wire _03883_;
 wire _03884_;
 wire _03885_;
 wire _03886_;
 wire _03887_;
 wire _03888_;
 wire _03889_;
 wire _03890_;
 wire _03891_;
 wire _03892_;
 wire _03893_;
 wire _03894_;
 wire _03895_;
 wire _03896_;
 wire _03897_;
 wire _03898_;
 wire _03899_;
 wire _03900_;
 wire _03901_;
 wire _03902_;
 wire _03903_;
 wire _03904_;
 wire _03905_;
 wire _03906_;
 wire _03907_;
 wire _03908_;
 wire _03909_;
 wire _03910_;
 wire _03911_;
 wire _03912_;
 wire _03913_;
 wire _03914_;
 wire _03915_;
 wire _03916_;
 wire _03917_;
 wire _03918_;
 wire _03919_;
 wire _03920_;
 wire _03921_;
 wire _03922_;
 wire _03923_;
 wire _03924_;
 wire _03925_;
 wire _03926_;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net865;
 wire net866;
 wire net867;
 wire net868;
 wire net869;
 wire net870;
 wire net871;
 wire net872;
 wire net873;
 wire net874;
 wire net875;
 wire net876;
 wire net877;
 wire net878;
 wire net879;
 wire net880;
 wire net881;
 wire net882;
 wire net883;
 wire net884;
 wire net885;
 wire net886;
 wire net887;
 wire net888;
 wire net889;
 wire net890;
 wire net891;
 wire net892;
 wire net893;
 wire net894;
 wire net895;
 wire net896;
 wire net897;
 wire net898;
 wire net899;
 wire net900;
 wire net901;
 wire net902;
 wire net903;
 wire net904;
 wire net905;
 wire net906;
 wire net907;
 wire net908;
 wire net909;
 wire net910;
 wire net911;
 wire net912;
 wire net913;
 wire net914;
 wire net915;
 wire net916;
 wire net917;
 wire net918;
 wire net919;
 wire net920;
 wire net921;
 wire net922;
 wire net923;
 wire net924;
 wire net925;
 wire net926;
 wire net927;
 wire net928;
 wire net929;
 wire net930;
 wire net931;
 wire net932;
 wire net933;
 wire net934;
 wire net935;
 wire net936;
 wire net937;
 wire net938;
 wire net939;
 wire net940;
 wire net941;
 wire net942;
 wire net943;
 wire net944;
 wire net945;
 wire net946;
 wire net947;
 wire net948;
 wire net949;
 wire net950;
 wire net951;
 wire net952;
 wire net953;
 wire net954;
 wire net955;
 wire net956;
 wire net957;
 wire net958;
 wire net959;
 wire net960;
 wire net961;
 wire net962;
 wire net963;
 wire net964;
 wire net965;
 wire net966;
 wire net967;
 wire net968;
 wire net969;
 wire net970;
 wire net971;
 wire net972;
 wire net973;
 wire net974;
 wire net975;
 wire net976;
 wire net977;
 wire net978;
 wire net979;
 wire net980;
 wire net981;
 wire net982;
 wire net983;
 wire net984;
 wire net985;
 wire net986;
 wire net987;
 wire net988;
 wire net989;
 wire net990;
 wire net991;
 wire net992;
 wire net993;
 wire net994;
 wire net995;
 wire net996;
 wire net997;
 wire net998;
 wire net999;
 wire net1000;
 wire net1001;
 wire net1002;
 wire net1003;
 wire net1004;
 wire net1005;
 wire net1006;
 wire net1007;
 wire net1008;
 wire net1009;
 wire net1010;
 wire net1011;
 wire net1012;
 wire net1013;
 wire net1014;
 wire net1015;
 wire net1016;
 wire net1017;
 wire net1018;
 wire net1019;
 wire net1020;
 wire net1021;
 wire net1022;
 wire net1023;
 wire net1024;
 wire net1025;
 wire net1026;
 wire net1027;
 wire net1028;
 wire net1029;
 wire net1030;
 wire net1031;
 wire net1032;
 wire net1033;
 wire net1034;
 wire net1035;
 wire net1036;
 wire net1037;
 wire net1038;
 wire net1039;
 wire net1040;
 wire net1041;
 wire net1042;
 wire net1043;
 wire net1044;
 wire net1045;
 wire net1046;
 wire net1047;
 wire net1048;
 wire net1049;
 wire net1050;
 wire net1051;
 wire net1052;
 wire net1053;
 wire net1054;
 wire net1055;
 wire net1056;
 wire net1057;
 wire net1058;
 wire net1059;
 wire net1060;
 wire net1061;
 wire net1062;
 wire net1063;
 wire net1064;
 wire net1065;
 wire net1066;
 wire net1067;
 wire net1068;
 wire net1069;
 wire net1070;
 wire net1071;
 wire net1072;
 wire net1073;
 wire net1074;
 wire net1075;
 wire net1076;
 wire net1077;
 wire net1078;
 wire net1079;
 wire net1080;
 wire net1081;
 wire net1082;
 wire net1083;
 wire net1084;
 wire net1085;
 wire net1086;
 wire net1087;
 wire net1088;
 wire net1089;
 wire net1090;
 wire net1091;
 wire net1092;
 wire net1093;
 wire net1094;
 wire net1095;
 wire net1096;
 wire net1097;
 wire net1098;
 wire net1099;
 wire net1100;
 wire net1101;
 wire net1102;
 wire net1103;
 wire net1104;
 wire net1105;
 wire net1106;
 wire net1107;
 wire net1108;
 wire net1109;
 wire net1110;
 wire net1111;
 wire net1112;
 wire net1113;
 wire net1114;
 wire net1115;
 wire net1116;
 wire net1117;
 wire net1118;
 wire net1119;
 wire net1120;
 wire net1121;
 wire net1122;
 wire net1123;
 wire net1124;
 wire net1125;
 wire net1126;
 wire net1127;
 wire net1128;
 wire net1129;
 wire net1130;
 wire net1131;
 wire net1132;
 wire net1133;
 wire net1134;
 wire net1135;
 wire net1136;
 wire net1137;
 wire net1138;
 wire net1139;
 wire net1140;
 wire net1141;
 wire net1142;
 wire net1143;
 wire net1144;
 wire net1145;
 wire net1146;
 wire net1147;
 wire net1148;
 wire net1149;
 wire net1150;
 wire net1151;
 wire net1152;
 wire net1153;
 wire net1154;
 wire net1155;
 wire net1156;
 wire net1157;
 wire net1158;
 wire net1159;
 wire net1160;
 wire net1161;
 wire net1162;
 wire net1163;
 wire net1164;
 wire net1165;
 wire net1166;
 wire net1167;
 wire net1168;
 wire net1169;
 wire net1170;
 wire net1171;
 wire net1172;
 wire net1173;
 wire net1174;
 wire net1175;
 wire net1176;
 wire net1177;
 wire net1178;
 wire net1179;
 wire net1180;
 wire net1181;
 wire net1182;
 wire net1183;
 wire net1184;
 wire net1185;
 wire net1186;
 wire net1187;
 wire net1188;
 wire net1189;
 wire net1190;
 wire net1191;
 wire net1192;
 wire net1193;
 wire net1194;
 wire net1195;
 wire net1196;
 wire net1197;
 wire net1198;
 wire net1199;
 wire net1200;
 wire net1201;
 wire net1202;
 wire net1203;
 wire net1204;
 wire net1205;
 wire net1206;
 wire net1207;
 wire net1208;
 wire net1209;
 wire net1210;
 wire net1211;
 wire net1212;
 wire net1213;
 wire net1214;
 wire net1215;
 wire net1216;
 wire net1217;
 wire net1218;
 wire net1219;
 wire net1220;
 wire net1221;
 wire net1222;
 wire net1223;
 wire net1224;
 wire net1225;
 wire net1226;
 wire net1227;
 wire net1228;
 wire net1229;
 wire net1230;
 wire net1231;
 wire net1232;
 wire net1233;
 wire net1234;
 wire net1235;
 wire net1236;
 wire net1237;
 wire net1238;
 wire net1239;
 wire net1240;
 wire net1241;
 wire net1242;
 wire net1243;
 wire net1244;
 wire net1245;
 wire net1246;
 wire net1247;
 wire net1248;
 wire net1249;
 wire net1250;
 wire net1251;
 wire net1252;
 wire net1253;
 wire net1254;
 wire net1255;
 wire net1256;
 wire net1257;
 wire net1258;
 wire net1259;
 wire net1260;
 wire net1261;
 wire net1262;
 wire net1263;
 wire net1264;
 wire net1265;
 wire net1266;
 wire net1267;
 wire net1268;
 wire net1269;
 wire net1270;
 wire net1271;
 wire net1272;
 wire net1273;
 wire net1274;
 wire net1275;
 wire net1276;
 wire net1277;
 wire net1278;
 wire net1279;
 wire net1280;
 wire net1281;
 wire net1282;
 wire net1283;
 wire net1284;
 wire net1285;
 wire net1286;
 wire net1287;
 wire net1288;
 wire net1289;
 wire net1290;
 wire net1291;
 wire net1292;
 wire net1293;
 wire net1294;
 wire net1295;
 wire net1296;
 wire net1297;
 wire net1298;
 wire net1299;
 wire net1300;
 wire net1301;
 wire net1302;
 wire net1303;
 wire net1304;
 wire net1305;
 wire net1306;
 wire net1307;
 wire net1308;
 wire net1309;
 wire net1310;
 wire net1311;
 wire net1312;
 wire net1313;
 wire net1314;
 wire net1315;
 wire net1316;
 wire net1317;
 wire net1318;
 wire net1319;
 wire net1320;
 wire net1321;
 wire net1322;
 wire net1323;
 wire net1324;
 wire net1325;
 wire net1326;
 wire net1327;
 wire net1328;
 wire net1329;
 wire net1330;
 wire net1331;
 wire net1332;
 wire net1333;
 wire net1334;
 wire net1335;
 wire net1336;
 wire net1337;
 wire net1338;
 wire net1339;
 wire net1340;
 wire net1341;
 wire net1342;
 wire net1343;
 wire net1344;
 wire net1345;
 wire net1346;
 wire net1347;
 wire net1348;
 wire net1349;
 wire net1350;
 wire net1351;
 wire net1352;
 wire net1353;
 wire net1354;
 wire net1355;
 wire net1356;
 wire net1357;
 wire net1358;
 wire net1359;
 wire net1360;
 wire net1361;
 wire net1362;
 wire net1363;
 wire net1364;
 wire net1365;
 wire net1366;
 wire net1367;
 wire net1368;
 wire net1369;
 wire net1370;
 wire net1371;
 wire net1372;
 wire net1373;
 wire net1374;
 wire \cpu.arbiter.i_wb_cpu_dbus_adr[10] ;
 wire \cpu.arbiter.i_wb_cpu_dbus_adr[11] ;
 wire \cpu.arbiter.i_wb_cpu_dbus_adr[12] ;
 wire \cpu.arbiter.i_wb_cpu_dbus_adr[13] ;
 wire \cpu.arbiter.i_wb_cpu_dbus_adr[14] ;
 wire \cpu.arbiter.i_wb_cpu_dbus_adr[15] ;
 wire \cpu.arbiter.i_wb_cpu_dbus_adr[16] ;
 wire \cpu.arbiter.i_wb_cpu_dbus_adr[17] ;
 wire \cpu.arbiter.i_wb_cpu_dbus_adr[18] ;
 wire \cpu.arbiter.i_wb_cpu_dbus_adr[19] ;
 wire \cpu.arbiter.i_wb_cpu_dbus_adr[20] ;
 wire \cpu.arbiter.i_wb_cpu_dbus_adr[21] ;
 wire \cpu.arbiter.i_wb_cpu_dbus_adr[22] ;
 wire \cpu.arbiter.i_wb_cpu_dbus_adr[23] ;
 wire \cpu.arbiter.i_wb_cpu_dbus_adr[24] ;
 wire \cpu.arbiter.i_wb_cpu_dbus_adr[25] ;
 wire \cpu.arbiter.i_wb_cpu_dbus_adr[26] ;
 wire \cpu.arbiter.i_wb_cpu_dbus_adr[27] ;
 wire \cpu.arbiter.i_wb_cpu_dbus_adr[28] ;
 wire \cpu.arbiter.i_wb_cpu_dbus_adr[29] ;
 wire \cpu.arbiter.i_wb_cpu_dbus_adr[2] ;
 wire \cpu.arbiter.i_wb_cpu_dbus_adr[30] ;
 wire \cpu.arbiter.i_wb_cpu_dbus_adr[31] ;
 wire \cpu.arbiter.i_wb_cpu_dbus_adr[3] ;
 wire \cpu.arbiter.i_wb_cpu_dbus_adr[4] ;
 wire \cpu.arbiter.i_wb_cpu_dbus_adr[5] ;
 wire \cpu.arbiter.i_wb_cpu_dbus_adr[6] ;
 wire \cpu.arbiter.i_wb_cpu_dbus_adr[7] ;
 wire \cpu.arbiter.i_wb_cpu_dbus_adr[8] ;
 wire \cpu.arbiter.i_wb_cpu_dbus_adr[9] ;
 wire \cpu.arbiter.i_wb_cpu_dbus_dat[0] ;
 wire \cpu.arbiter.i_wb_cpu_dbus_dat[10] ;
 wire \cpu.arbiter.i_wb_cpu_dbus_dat[11] ;
 wire \cpu.arbiter.i_wb_cpu_dbus_dat[12] ;
 wire \cpu.arbiter.i_wb_cpu_dbus_dat[13] ;
 wire \cpu.arbiter.i_wb_cpu_dbus_dat[14] ;
 wire \cpu.arbiter.i_wb_cpu_dbus_dat[15] ;
 wire \cpu.arbiter.i_wb_cpu_dbus_dat[16] ;
 wire \cpu.arbiter.i_wb_cpu_dbus_dat[17] ;
 wire \cpu.arbiter.i_wb_cpu_dbus_dat[18] ;
 wire \cpu.arbiter.i_wb_cpu_dbus_dat[19] ;
 wire \cpu.arbiter.i_wb_cpu_dbus_dat[1] ;
 wire \cpu.arbiter.i_wb_cpu_dbus_dat[20] ;
 wire \cpu.arbiter.i_wb_cpu_dbus_dat[21] ;
 wire \cpu.arbiter.i_wb_cpu_dbus_dat[22] ;
 wire \cpu.arbiter.i_wb_cpu_dbus_dat[23] ;
 wire \cpu.arbiter.i_wb_cpu_dbus_dat[24] ;
 wire \cpu.arbiter.i_wb_cpu_dbus_dat[25] ;
 wire \cpu.arbiter.i_wb_cpu_dbus_dat[26] ;
 wire \cpu.arbiter.i_wb_cpu_dbus_dat[27] ;
 wire \cpu.arbiter.i_wb_cpu_dbus_dat[28] ;
 wire \cpu.arbiter.i_wb_cpu_dbus_dat[29] ;
 wire \cpu.arbiter.i_wb_cpu_dbus_dat[2] ;
 wire \cpu.arbiter.i_wb_cpu_dbus_dat[30] ;
 wire \cpu.arbiter.i_wb_cpu_dbus_dat[31] ;
 wire \cpu.arbiter.i_wb_cpu_dbus_dat[3] ;
 wire \cpu.arbiter.i_wb_cpu_dbus_dat[4] ;
 wire \cpu.arbiter.i_wb_cpu_dbus_dat[5] ;
 wire \cpu.arbiter.i_wb_cpu_dbus_dat[6] ;
 wire \cpu.arbiter.i_wb_cpu_dbus_dat[7] ;
 wire \cpu.arbiter.i_wb_cpu_dbus_dat[8] ;
 wire \cpu.arbiter.i_wb_cpu_dbus_dat[9] ;
 wire \cpu.arbiter.i_wb_cpu_dbus_we ;
 wire \cpu.arbiter.i_wb_cpu_ibus_adr[10] ;
 wire \cpu.arbiter.i_wb_cpu_ibus_adr[11] ;
 wire \cpu.arbiter.i_wb_cpu_ibus_adr[12] ;
 wire \cpu.arbiter.i_wb_cpu_ibus_adr[13] ;
 wire \cpu.arbiter.i_wb_cpu_ibus_adr[14] ;
 wire \cpu.arbiter.i_wb_cpu_ibus_adr[15] ;
 wire \cpu.arbiter.i_wb_cpu_ibus_adr[16] ;
 wire \cpu.arbiter.i_wb_cpu_ibus_adr[17] ;
 wire \cpu.arbiter.i_wb_cpu_ibus_adr[18] ;
 wire \cpu.arbiter.i_wb_cpu_ibus_adr[19] ;
 wire \cpu.arbiter.i_wb_cpu_ibus_adr[1] ;
 wire \cpu.arbiter.i_wb_cpu_ibus_adr[20] ;
 wire \cpu.arbiter.i_wb_cpu_ibus_adr[21] ;
 wire \cpu.arbiter.i_wb_cpu_ibus_adr[22] ;
 wire \cpu.arbiter.i_wb_cpu_ibus_adr[23] ;
 wire \cpu.arbiter.i_wb_cpu_ibus_adr[24] ;
 wire \cpu.arbiter.i_wb_cpu_ibus_adr[25] ;
 wire \cpu.arbiter.i_wb_cpu_ibus_adr[26] ;
 wire \cpu.arbiter.i_wb_cpu_ibus_adr[27] ;
 wire \cpu.arbiter.i_wb_cpu_ibus_adr[28] ;
 wire \cpu.arbiter.i_wb_cpu_ibus_adr[29] ;
 wire \cpu.arbiter.i_wb_cpu_ibus_adr[2] ;
 wire \cpu.arbiter.i_wb_cpu_ibus_adr[30] ;
 wire \cpu.arbiter.i_wb_cpu_ibus_adr[31] ;
 wire \cpu.arbiter.i_wb_cpu_ibus_adr[3] ;
 wire \cpu.arbiter.i_wb_cpu_ibus_adr[4] ;
 wire \cpu.arbiter.i_wb_cpu_ibus_adr[5] ;
 wire \cpu.arbiter.i_wb_cpu_ibus_adr[6] ;
 wire \cpu.arbiter.i_wb_cpu_ibus_adr[7] ;
 wire \cpu.arbiter.i_wb_cpu_ibus_adr[8] ;
 wire \cpu.arbiter.i_wb_cpu_ibus_adr[9] ;
 wire \cpu.arbiter.i_wb_mem_rdt[0] ;
 wire \cpu.arbiter.i_wb_mem_rdt[10] ;
 wire \cpu.arbiter.i_wb_mem_rdt[11] ;
 wire \cpu.arbiter.i_wb_mem_rdt[12] ;
 wire \cpu.arbiter.i_wb_mem_rdt[13] ;
 wire \cpu.arbiter.i_wb_mem_rdt[14] ;
 wire \cpu.arbiter.i_wb_mem_rdt[15] ;
 wire \cpu.arbiter.i_wb_mem_rdt[16] ;
 wire \cpu.arbiter.i_wb_mem_rdt[17] ;
 wire \cpu.arbiter.i_wb_mem_rdt[18] ;
 wire \cpu.arbiter.i_wb_mem_rdt[19] ;
 wire \cpu.arbiter.i_wb_mem_rdt[1] ;
 wire \cpu.arbiter.i_wb_mem_rdt[20] ;
 wire \cpu.arbiter.i_wb_mem_rdt[21] ;
 wire \cpu.arbiter.i_wb_mem_rdt[22] ;
 wire \cpu.arbiter.i_wb_mem_rdt[23] ;
 wire \cpu.arbiter.i_wb_mem_rdt[24] ;
 wire \cpu.arbiter.i_wb_mem_rdt[25] ;
 wire \cpu.arbiter.i_wb_mem_rdt[26] ;
 wire \cpu.arbiter.i_wb_mem_rdt[27] ;
 wire \cpu.arbiter.i_wb_mem_rdt[28] ;
 wire \cpu.arbiter.i_wb_mem_rdt[29] ;
 wire \cpu.arbiter.i_wb_mem_rdt[2] ;
 wire \cpu.arbiter.i_wb_mem_rdt[30] ;
 wire \cpu.arbiter.i_wb_mem_rdt[31] ;
 wire \cpu.arbiter.i_wb_mem_rdt[3] ;
 wire \cpu.arbiter.i_wb_mem_rdt[4] ;
 wire \cpu.arbiter.i_wb_mem_rdt[5] ;
 wire \cpu.arbiter.i_wb_mem_rdt[6] ;
 wire \cpu.arbiter.i_wb_mem_rdt[7] ;
 wire \cpu.arbiter.i_wb_mem_rdt[8] ;
 wire \cpu.arbiter.i_wb_mem_rdt[9] ;
 wire \cpu.cpu.alu.cmp_r ;
 wire \cpu.cpu.bne_or_bge ;
 wire \cpu.cpu.branch_op ;
 wire \cpu.cpu.bufreg.data[0] ;
 wire \cpu.cpu.bufreg.data[1] ;
 wire \cpu.cpu.bufreg.i_right_shift_op ;
 wire \cpu.cpu.bufreg.i_sh_signed ;
 wire \cpu.cpu.bufreg2.i_bytecnt[0] ;
 wire \cpu.cpu.bufreg2.i_bytecnt[1] ;
 wire \cpu.cpu.ctrl.i_jump ;
 wire \cpu.cpu.decode.co_ebreak ;
 wire \cpu.cpu.decode.co_mem_word ;
 wire \cpu.cpu.decode.opcode[0] ;
 wire \cpu.cpu.decode.opcode[1] ;
 wire \cpu.cpu.decode.opcode[2] ;
 wire \cpu.cpu.immdec.gen_immdec_w_eq_1.imm11_7[0] ;
 wire \cpu.cpu.immdec.gen_immdec_w_eq_1.imm11_7[1] ;
 wire \cpu.cpu.immdec.gen_immdec_w_eq_1.imm11_7[2] ;
 wire \cpu.cpu.immdec.gen_immdec_w_eq_1.imm11_7[3] ;
 wire \cpu.cpu.immdec.gen_immdec_w_eq_1.imm11_7[4] ;
 wire \cpu.cpu.immdec.gen_immdec_w_eq_1.imm19_12_20[0] ;
 wire \cpu.cpu.immdec.gen_immdec_w_eq_1.imm19_12_20[1] ;
 wire \cpu.cpu.immdec.gen_immdec_w_eq_1.imm19_12_20[2] ;
 wire \cpu.cpu.immdec.gen_immdec_w_eq_1.imm19_12_20[3] ;
 wire \cpu.cpu.immdec.gen_immdec_w_eq_1.imm19_12_20[5] ;
 wire \cpu.cpu.immdec.gen_immdec_w_eq_1.imm19_12_20[6] ;
 wire \cpu.cpu.immdec.gen_immdec_w_eq_1.imm19_12_20[7] ;
 wire \cpu.cpu.immdec.gen_immdec_w_eq_1.imm19_12_20[8] ;
 wire \cpu.cpu.immdec.gen_immdec_w_eq_1.imm24_20[0] ;
 wire \cpu.cpu.immdec.gen_immdec_w_eq_1.imm24_20[1] ;
 wire \cpu.cpu.immdec.gen_immdec_w_eq_1.imm24_20[2] ;
 wire \cpu.cpu.immdec.gen_immdec_w_eq_1.imm24_20[3] ;
 wire \cpu.cpu.immdec.gen_immdec_w_eq_1.imm24_20[4] ;
 wire \cpu.cpu.immdec.gen_immdec_w_eq_1.imm30_25[0] ;
 wire \cpu.cpu.immdec.gen_immdec_w_eq_1.imm30_25[1] ;
 wire \cpu.cpu.immdec.gen_immdec_w_eq_1.imm30_25[2] ;
 wire \cpu.cpu.immdec.gen_immdec_w_eq_1.imm30_25[3] ;
 wire \cpu.cpu.immdec.gen_immdec_w_eq_1.imm30_25[4] ;
 wire \cpu.cpu.immdec.gen_immdec_w_eq_1.imm30_25[5] ;
 wire \cpu.cpu.immdec.gen_immdec_w_eq_1.imm31 ;
 wire \cpu.cpu.immdec.gen_immdec_w_eq_1.imm7 ;
 wire \cpu.cpu.mem_if.signbit ;
 wire \cpu.cpu.state.cnt_r[0] ;
 wire \cpu.cpu.state.cnt_r[1] ;
 wire \cpu.cpu.state.cnt_r[2] ;
 wire \cpu.cpu.state.cnt_r[3] ;
 wire \cpu.cpu.state.ibus_cyc ;
 wire \cpu.cpu.state.init_done ;
 wire \cpu.cpu.state.o_cnt[2] ;
 wire \cpu.i_rf_rdata[0] ;
 wire \cpu.i_rf_rdata[10] ;
 wire \cpu.i_rf_rdata[11] ;
 wire \cpu.i_rf_rdata[12] ;
 wire \cpu.i_rf_rdata[13] ;
 wire \cpu.i_rf_rdata[14] ;
 wire \cpu.i_rf_rdata[15] ;
 wire \cpu.i_rf_rdata[16] ;
 wire \cpu.i_rf_rdata[17] ;
 wire \cpu.i_rf_rdata[18] ;
 wire \cpu.i_rf_rdata[19] ;
 wire \cpu.i_rf_rdata[1] ;
 wire \cpu.i_rf_rdata[20] ;
 wire \cpu.i_rf_rdata[21] ;
 wire \cpu.i_rf_rdata[22] ;
 wire \cpu.i_rf_rdata[23] ;
 wire \cpu.i_rf_rdata[24] ;
 wire \cpu.i_rf_rdata[25] ;
 wire \cpu.i_rf_rdata[26] ;
 wire \cpu.i_rf_rdata[27] ;
 wire \cpu.i_rf_rdata[28] ;
 wire \cpu.i_rf_rdata[29] ;
 wire \cpu.i_rf_rdata[2] ;
 wire \cpu.i_rf_rdata[30] ;
 wire \cpu.i_rf_rdata[31] ;
 wire \cpu.i_rf_rdata[3] ;
 wire \cpu.i_rf_rdata[4] ;
 wire \cpu.i_rf_rdata[5] ;
 wire \cpu.i_rf_rdata[6] ;
 wire \cpu.i_rf_rdata[7] ;
 wire \cpu.i_rf_rdata[8] ;
 wire \cpu.i_rf_rdata[9] ;
 wire \cpu.i_wb_ext_rdt[0] ;
 wire \cpu.i_wb_ext_rdt[1] ;
 wire \cpu.i_wb_ext_rdt[2] ;
 wire \cpu.i_wb_ext_rdt[3] ;
 wire \cpu.i_wb_ext_rdt[4] ;
 wire \cpu.i_wb_ext_rdt[5] ;
 wire \cpu.i_wb_ext_rdt[6] ;
 wire \cpu.i_wb_ext_rdt[7] ;
 wire \cpu.rf_ram_if.gen_wtrig_ratio_neq_2.wtrig0_r ;
 wire \cpu.rf_ram_if.rcnt[0] ;
 wire \cpu.rf_ram_if.rcnt[1] ;
 wire \cpu.rf_ram_if.rcnt[2] ;
 wire \cpu.rf_ram_if.rcnt[3] ;
 wire \cpu.rf_ram_if.rcnt[4] ;
 wire \cpu.rf_ram_if.rdata0[10] ;
 wire \cpu.rf_ram_if.rdata0[11] ;
 wire \cpu.rf_ram_if.rdata0[12] ;
 wire \cpu.rf_ram_if.rdata0[13] ;
 wire \cpu.rf_ram_if.rdata0[14] ;
 wire \cpu.rf_ram_if.rdata0[15] ;
 wire \cpu.rf_ram_if.rdata0[16] ;
 wire \cpu.rf_ram_if.rdata0[17] ;
 wire \cpu.rf_ram_if.rdata0[18] ;
 wire \cpu.rf_ram_if.rdata0[19] ;
 wire \cpu.rf_ram_if.rdata0[1] ;
 wire \cpu.rf_ram_if.rdata0[20] ;
 wire \cpu.rf_ram_if.rdata0[21] ;
 wire \cpu.rf_ram_if.rdata0[22] ;
 wire \cpu.rf_ram_if.rdata0[23] ;
 wire \cpu.rf_ram_if.rdata0[24] ;
 wire \cpu.rf_ram_if.rdata0[25] ;
 wire \cpu.rf_ram_if.rdata0[26] ;
 wire \cpu.rf_ram_if.rdata0[27] ;
 wire \cpu.rf_ram_if.rdata0[28] ;
 wire \cpu.rf_ram_if.rdata0[29] ;
 wire \cpu.rf_ram_if.rdata0[2] ;
 wire \cpu.rf_ram_if.rdata0[30] ;
 wire \cpu.rf_ram_if.rdata0[31] ;
 wire \cpu.rf_ram_if.rdata0[3] ;
 wire \cpu.rf_ram_if.rdata0[4] ;
 wire \cpu.rf_ram_if.rdata0[5] ;
 wire \cpu.rf_ram_if.rdata0[6] ;
 wire \cpu.rf_ram_if.rdata0[7] ;
 wire \cpu.rf_ram_if.rdata0[8] ;
 wire \cpu.rf_ram_if.rdata0[9] ;
 wire \cpu.rf_ram_if.rdata1[0] ;
 wire \cpu.rf_ram_if.rdata1[10] ;
 wire \cpu.rf_ram_if.rdata1[11] ;
 wire \cpu.rf_ram_if.rdata1[12] ;
 wire \cpu.rf_ram_if.rdata1[13] ;
 wire \cpu.rf_ram_if.rdata1[14] ;
 wire \cpu.rf_ram_if.rdata1[15] ;
 wire \cpu.rf_ram_if.rdata1[16] ;
 wire \cpu.rf_ram_if.rdata1[17] ;
 wire \cpu.rf_ram_if.rdata1[18] ;
 wire \cpu.rf_ram_if.rdata1[19] ;
 wire \cpu.rf_ram_if.rdata1[1] ;
 wire \cpu.rf_ram_if.rdata1[20] ;
 wire \cpu.rf_ram_if.rdata1[21] ;
 wire \cpu.rf_ram_if.rdata1[22] ;
 wire \cpu.rf_ram_if.rdata1[23] ;
 wire \cpu.rf_ram_if.rdata1[24] ;
 wire \cpu.rf_ram_if.rdata1[25] ;
 wire \cpu.rf_ram_if.rdata1[26] ;
 wire \cpu.rf_ram_if.rdata1[27] ;
 wire \cpu.rf_ram_if.rdata1[28] ;
 wire \cpu.rf_ram_if.rdata1[29] ;
 wire \cpu.rf_ram_if.rdata1[2] ;
 wire \cpu.rf_ram_if.rdata1[30] ;
 wire \cpu.rf_ram_if.rdata1[3] ;
 wire \cpu.rf_ram_if.rdata1[4] ;
 wire \cpu.rf_ram_if.rdata1[5] ;
 wire \cpu.rf_ram_if.rdata1[6] ;
 wire \cpu.rf_ram_if.rdata1[7] ;
 wire \cpu.rf_ram_if.rdata1[8] ;
 wire \cpu.rf_ram_if.rdata1[9] ;
 wire \cpu.rf_ram_if.rgate ;
 wire \cpu.rf_ram_if.rgnt ;
 wire \cpu.rf_ram_if.rreq_r ;
 wire \cpu.rf_ram_if.rtrig0 ;
 wire \cpu.rf_ram_if.rtrig1 ;
 wire \cpu.rf_ram_if.wdata0_r[0] ;
 wire \cpu.rf_ram_if.wdata0_r[10] ;
 wire \cpu.rf_ram_if.wdata0_r[11] ;
 wire \cpu.rf_ram_if.wdata0_r[12] ;
 wire \cpu.rf_ram_if.wdata0_r[13] ;
 wire \cpu.rf_ram_if.wdata0_r[14] ;
 wire \cpu.rf_ram_if.wdata0_r[15] ;
 wire \cpu.rf_ram_if.wdata0_r[16] ;
 wire \cpu.rf_ram_if.wdata0_r[17] ;
 wire \cpu.rf_ram_if.wdata0_r[18] ;
 wire \cpu.rf_ram_if.wdata0_r[19] ;
 wire \cpu.rf_ram_if.wdata0_r[1] ;
 wire \cpu.rf_ram_if.wdata0_r[20] ;
 wire \cpu.rf_ram_if.wdata0_r[21] ;
 wire \cpu.rf_ram_if.wdata0_r[22] ;
 wire \cpu.rf_ram_if.wdata0_r[23] ;
 wire \cpu.rf_ram_if.wdata0_r[24] ;
 wire \cpu.rf_ram_if.wdata0_r[25] ;
 wire \cpu.rf_ram_if.wdata0_r[26] ;
 wire \cpu.rf_ram_if.wdata0_r[27] ;
 wire \cpu.rf_ram_if.wdata0_r[28] ;
 wire \cpu.rf_ram_if.wdata0_r[29] ;
 wire \cpu.rf_ram_if.wdata0_r[2] ;
 wire \cpu.rf_ram_if.wdata0_r[30] ;
 wire \cpu.rf_ram_if.wdata0_r[31] ;
 wire \cpu.rf_ram_if.wdata0_r[3] ;
 wire \cpu.rf_ram_if.wdata0_r[4] ;
 wire \cpu.rf_ram_if.wdata0_r[5] ;
 wire \cpu.rf_ram_if.wdata0_r[6] ;
 wire \cpu.rf_ram_if.wdata0_r[7] ;
 wire \cpu.rf_ram_if.wdata0_r[8] ;
 wire \cpu.rf_ram_if.wdata0_r[9] ;
 wire \cpu.rf_ram_if.wen0_r ;
 wire \ram_spi_if.cycle_counter[0] ;
 wire \ram_spi_if.cycle_counter[1] ;
 wire \ram_spi_if.cycle_counter[2] ;
 wire \ram_spi_if.cycle_counter[3] ;
 wire \ram_spi_if.cycle_counter[4] ;
 wire \ram_spi_if.cycle_counter[5] ;
 wire \ram_spi_if.spi_clk ;
 wire \ram_spi_if.spi_cs_n ;
 wire \ram_spi_if.spi_mosi ;
 wire \ram_spi_if.state_reg[0] ;
 wire \ram_spi_if.state_reg[1] ;
 wire \ram_spi_if.state_reg[2] ;
 wire \ram_spi_if.state_reg[3] ;
 wire \rf_ram.RAM[0][0] ;
 wire \rf_ram.RAM[0][10] ;
 wire \rf_ram.RAM[0][11] ;
 wire \rf_ram.RAM[0][12] ;
 wire \rf_ram.RAM[0][13] ;
 wire \rf_ram.RAM[0][14] ;
 wire \rf_ram.RAM[0][15] ;
 wire \rf_ram.RAM[0][16] ;
 wire \rf_ram.RAM[0][17] ;
 wire \rf_ram.RAM[0][18] ;
 wire \rf_ram.RAM[0][19] ;
 wire \rf_ram.RAM[0][1] ;
 wire \rf_ram.RAM[0][20] ;
 wire \rf_ram.RAM[0][21] ;
 wire \rf_ram.RAM[0][22] ;
 wire \rf_ram.RAM[0][23] ;
 wire \rf_ram.RAM[0][24] ;
 wire \rf_ram.RAM[0][25] ;
 wire \rf_ram.RAM[0][26] ;
 wire \rf_ram.RAM[0][27] ;
 wire \rf_ram.RAM[0][28] ;
 wire \rf_ram.RAM[0][29] ;
 wire \rf_ram.RAM[0][2] ;
 wire \rf_ram.RAM[0][30] ;
 wire \rf_ram.RAM[0][31] ;
 wire \rf_ram.RAM[0][3] ;
 wire \rf_ram.RAM[0][4] ;
 wire \rf_ram.RAM[0][5] ;
 wire \rf_ram.RAM[0][6] ;
 wire \rf_ram.RAM[0][7] ;
 wire \rf_ram.RAM[0][8] ;
 wire \rf_ram.RAM[0][9] ;
 wire \rf_ram.RAM[10][0] ;
 wire \rf_ram.RAM[10][10] ;
 wire \rf_ram.RAM[10][11] ;
 wire \rf_ram.RAM[10][12] ;
 wire \rf_ram.RAM[10][13] ;
 wire \rf_ram.RAM[10][14] ;
 wire \rf_ram.RAM[10][15] ;
 wire \rf_ram.RAM[10][16] ;
 wire \rf_ram.RAM[10][17] ;
 wire \rf_ram.RAM[10][18] ;
 wire \rf_ram.RAM[10][19] ;
 wire \rf_ram.RAM[10][1] ;
 wire \rf_ram.RAM[10][20] ;
 wire \rf_ram.RAM[10][21] ;
 wire \rf_ram.RAM[10][22] ;
 wire \rf_ram.RAM[10][23] ;
 wire \rf_ram.RAM[10][24] ;
 wire \rf_ram.RAM[10][25] ;
 wire \rf_ram.RAM[10][26] ;
 wire \rf_ram.RAM[10][27] ;
 wire \rf_ram.RAM[10][28] ;
 wire \rf_ram.RAM[10][29] ;
 wire \rf_ram.RAM[10][2] ;
 wire \rf_ram.RAM[10][30] ;
 wire \rf_ram.RAM[10][31] ;
 wire \rf_ram.RAM[10][3] ;
 wire \rf_ram.RAM[10][4] ;
 wire \rf_ram.RAM[10][5] ;
 wire \rf_ram.RAM[10][6] ;
 wire \rf_ram.RAM[10][7] ;
 wire \rf_ram.RAM[10][8] ;
 wire \rf_ram.RAM[10][9] ;
 wire \rf_ram.RAM[11][0] ;
 wire \rf_ram.RAM[11][10] ;
 wire \rf_ram.RAM[11][11] ;
 wire \rf_ram.RAM[11][12] ;
 wire \rf_ram.RAM[11][13] ;
 wire \rf_ram.RAM[11][14] ;
 wire \rf_ram.RAM[11][15] ;
 wire \rf_ram.RAM[11][16] ;
 wire \rf_ram.RAM[11][17] ;
 wire \rf_ram.RAM[11][18] ;
 wire \rf_ram.RAM[11][19] ;
 wire \rf_ram.RAM[11][1] ;
 wire \rf_ram.RAM[11][20] ;
 wire \rf_ram.RAM[11][21] ;
 wire \rf_ram.RAM[11][22] ;
 wire \rf_ram.RAM[11][23] ;
 wire \rf_ram.RAM[11][24] ;
 wire \rf_ram.RAM[11][25] ;
 wire \rf_ram.RAM[11][26] ;
 wire \rf_ram.RAM[11][27] ;
 wire \rf_ram.RAM[11][28] ;
 wire \rf_ram.RAM[11][29] ;
 wire \rf_ram.RAM[11][2] ;
 wire \rf_ram.RAM[11][30] ;
 wire \rf_ram.RAM[11][31] ;
 wire \rf_ram.RAM[11][3] ;
 wire \rf_ram.RAM[11][4] ;
 wire \rf_ram.RAM[11][5] ;
 wire \rf_ram.RAM[11][6] ;
 wire \rf_ram.RAM[11][7] ;
 wire \rf_ram.RAM[11][8] ;
 wire \rf_ram.RAM[11][9] ;
 wire \rf_ram.RAM[12][0] ;
 wire \rf_ram.RAM[12][10] ;
 wire \rf_ram.RAM[12][11] ;
 wire \rf_ram.RAM[12][12] ;
 wire \rf_ram.RAM[12][13] ;
 wire \rf_ram.RAM[12][14] ;
 wire \rf_ram.RAM[12][15] ;
 wire \rf_ram.RAM[12][16] ;
 wire \rf_ram.RAM[12][17] ;
 wire \rf_ram.RAM[12][18] ;
 wire \rf_ram.RAM[12][19] ;
 wire \rf_ram.RAM[12][1] ;
 wire \rf_ram.RAM[12][20] ;
 wire \rf_ram.RAM[12][21] ;
 wire \rf_ram.RAM[12][22] ;
 wire \rf_ram.RAM[12][23] ;
 wire \rf_ram.RAM[12][24] ;
 wire \rf_ram.RAM[12][25] ;
 wire \rf_ram.RAM[12][26] ;
 wire \rf_ram.RAM[12][27] ;
 wire \rf_ram.RAM[12][28] ;
 wire \rf_ram.RAM[12][29] ;
 wire \rf_ram.RAM[12][2] ;
 wire \rf_ram.RAM[12][30] ;
 wire \rf_ram.RAM[12][31] ;
 wire \rf_ram.RAM[12][3] ;
 wire \rf_ram.RAM[12][4] ;
 wire \rf_ram.RAM[12][5] ;
 wire \rf_ram.RAM[12][6] ;
 wire \rf_ram.RAM[12][7] ;
 wire \rf_ram.RAM[12][8] ;
 wire \rf_ram.RAM[12][9] ;
 wire \rf_ram.RAM[13][0] ;
 wire \rf_ram.RAM[13][10] ;
 wire \rf_ram.RAM[13][11] ;
 wire \rf_ram.RAM[13][12] ;
 wire \rf_ram.RAM[13][13] ;
 wire \rf_ram.RAM[13][14] ;
 wire \rf_ram.RAM[13][15] ;
 wire \rf_ram.RAM[13][16] ;
 wire \rf_ram.RAM[13][17] ;
 wire \rf_ram.RAM[13][18] ;
 wire \rf_ram.RAM[13][19] ;
 wire \rf_ram.RAM[13][1] ;
 wire \rf_ram.RAM[13][20] ;
 wire \rf_ram.RAM[13][21] ;
 wire \rf_ram.RAM[13][22] ;
 wire \rf_ram.RAM[13][23] ;
 wire \rf_ram.RAM[13][24] ;
 wire \rf_ram.RAM[13][25] ;
 wire \rf_ram.RAM[13][26] ;
 wire \rf_ram.RAM[13][27] ;
 wire \rf_ram.RAM[13][28] ;
 wire \rf_ram.RAM[13][29] ;
 wire \rf_ram.RAM[13][2] ;
 wire \rf_ram.RAM[13][30] ;
 wire \rf_ram.RAM[13][31] ;
 wire \rf_ram.RAM[13][3] ;
 wire \rf_ram.RAM[13][4] ;
 wire \rf_ram.RAM[13][5] ;
 wire \rf_ram.RAM[13][6] ;
 wire \rf_ram.RAM[13][7] ;
 wire \rf_ram.RAM[13][8] ;
 wire \rf_ram.RAM[13][9] ;
 wire \rf_ram.RAM[14][0] ;
 wire \rf_ram.RAM[14][10] ;
 wire \rf_ram.RAM[14][11] ;
 wire \rf_ram.RAM[14][12] ;
 wire \rf_ram.RAM[14][13] ;
 wire \rf_ram.RAM[14][14] ;
 wire \rf_ram.RAM[14][15] ;
 wire \rf_ram.RAM[14][16] ;
 wire \rf_ram.RAM[14][17] ;
 wire \rf_ram.RAM[14][18] ;
 wire \rf_ram.RAM[14][19] ;
 wire \rf_ram.RAM[14][1] ;
 wire \rf_ram.RAM[14][20] ;
 wire \rf_ram.RAM[14][21] ;
 wire \rf_ram.RAM[14][22] ;
 wire \rf_ram.RAM[14][23] ;
 wire \rf_ram.RAM[14][24] ;
 wire \rf_ram.RAM[14][25] ;
 wire \rf_ram.RAM[14][26] ;
 wire \rf_ram.RAM[14][27] ;
 wire \rf_ram.RAM[14][28] ;
 wire \rf_ram.RAM[14][29] ;
 wire \rf_ram.RAM[14][2] ;
 wire \rf_ram.RAM[14][30] ;
 wire \rf_ram.RAM[14][31] ;
 wire \rf_ram.RAM[14][3] ;
 wire \rf_ram.RAM[14][4] ;
 wire \rf_ram.RAM[14][5] ;
 wire \rf_ram.RAM[14][6] ;
 wire \rf_ram.RAM[14][7] ;
 wire \rf_ram.RAM[14][8] ;
 wire \rf_ram.RAM[14][9] ;
 wire \rf_ram.RAM[15][0] ;
 wire \rf_ram.RAM[15][10] ;
 wire \rf_ram.RAM[15][11] ;
 wire \rf_ram.RAM[15][12] ;
 wire \rf_ram.RAM[15][13] ;
 wire \rf_ram.RAM[15][14] ;
 wire \rf_ram.RAM[15][15] ;
 wire \rf_ram.RAM[15][16] ;
 wire \rf_ram.RAM[15][17] ;
 wire \rf_ram.RAM[15][18] ;
 wire \rf_ram.RAM[15][19] ;
 wire \rf_ram.RAM[15][1] ;
 wire \rf_ram.RAM[15][20] ;
 wire \rf_ram.RAM[15][21] ;
 wire \rf_ram.RAM[15][22] ;
 wire \rf_ram.RAM[15][23] ;
 wire \rf_ram.RAM[15][24] ;
 wire \rf_ram.RAM[15][25] ;
 wire \rf_ram.RAM[15][26] ;
 wire \rf_ram.RAM[15][27] ;
 wire \rf_ram.RAM[15][28] ;
 wire \rf_ram.RAM[15][29] ;
 wire \rf_ram.RAM[15][2] ;
 wire \rf_ram.RAM[15][30] ;
 wire \rf_ram.RAM[15][31] ;
 wire \rf_ram.RAM[15][3] ;
 wire \rf_ram.RAM[15][4] ;
 wire \rf_ram.RAM[15][5] ;
 wire \rf_ram.RAM[15][6] ;
 wire \rf_ram.RAM[15][7] ;
 wire \rf_ram.RAM[15][8] ;
 wire \rf_ram.RAM[15][9] ;
 wire \rf_ram.RAM[16][0] ;
 wire \rf_ram.RAM[16][10] ;
 wire \rf_ram.RAM[16][11] ;
 wire \rf_ram.RAM[16][12] ;
 wire \rf_ram.RAM[16][13] ;
 wire \rf_ram.RAM[16][14] ;
 wire \rf_ram.RAM[16][15] ;
 wire \rf_ram.RAM[16][16] ;
 wire \rf_ram.RAM[16][17] ;
 wire \rf_ram.RAM[16][18] ;
 wire \rf_ram.RAM[16][19] ;
 wire \rf_ram.RAM[16][1] ;
 wire \rf_ram.RAM[16][20] ;
 wire \rf_ram.RAM[16][21] ;
 wire \rf_ram.RAM[16][22] ;
 wire \rf_ram.RAM[16][23] ;
 wire \rf_ram.RAM[16][24] ;
 wire \rf_ram.RAM[16][25] ;
 wire \rf_ram.RAM[16][26] ;
 wire \rf_ram.RAM[16][27] ;
 wire \rf_ram.RAM[16][28] ;
 wire \rf_ram.RAM[16][29] ;
 wire \rf_ram.RAM[16][2] ;
 wire \rf_ram.RAM[16][30] ;
 wire \rf_ram.RAM[16][31] ;
 wire \rf_ram.RAM[16][3] ;
 wire \rf_ram.RAM[16][4] ;
 wire \rf_ram.RAM[16][5] ;
 wire \rf_ram.RAM[16][6] ;
 wire \rf_ram.RAM[16][7] ;
 wire \rf_ram.RAM[16][8] ;
 wire \rf_ram.RAM[16][9] ;
 wire \rf_ram.RAM[17][0] ;
 wire \rf_ram.RAM[17][10] ;
 wire \rf_ram.RAM[17][11] ;
 wire \rf_ram.RAM[17][12] ;
 wire \rf_ram.RAM[17][13] ;
 wire \rf_ram.RAM[17][14] ;
 wire \rf_ram.RAM[17][15] ;
 wire \rf_ram.RAM[17][16] ;
 wire \rf_ram.RAM[17][17] ;
 wire \rf_ram.RAM[17][18] ;
 wire \rf_ram.RAM[17][19] ;
 wire \rf_ram.RAM[17][1] ;
 wire \rf_ram.RAM[17][20] ;
 wire \rf_ram.RAM[17][21] ;
 wire \rf_ram.RAM[17][22] ;
 wire \rf_ram.RAM[17][23] ;
 wire \rf_ram.RAM[17][24] ;
 wire \rf_ram.RAM[17][25] ;
 wire \rf_ram.RAM[17][26] ;
 wire \rf_ram.RAM[17][27] ;
 wire \rf_ram.RAM[17][28] ;
 wire \rf_ram.RAM[17][29] ;
 wire \rf_ram.RAM[17][2] ;
 wire \rf_ram.RAM[17][30] ;
 wire \rf_ram.RAM[17][31] ;
 wire \rf_ram.RAM[17][3] ;
 wire \rf_ram.RAM[17][4] ;
 wire \rf_ram.RAM[17][5] ;
 wire \rf_ram.RAM[17][6] ;
 wire \rf_ram.RAM[17][7] ;
 wire \rf_ram.RAM[17][8] ;
 wire \rf_ram.RAM[17][9] ;
 wire \rf_ram.RAM[18][0] ;
 wire \rf_ram.RAM[18][10] ;
 wire \rf_ram.RAM[18][11] ;
 wire \rf_ram.RAM[18][12] ;
 wire \rf_ram.RAM[18][13] ;
 wire \rf_ram.RAM[18][14] ;
 wire \rf_ram.RAM[18][15] ;
 wire \rf_ram.RAM[18][16] ;
 wire \rf_ram.RAM[18][17] ;
 wire \rf_ram.RAM[18][18] ;
 wire \rf_ram.RAM[18][19] ;
 wire \rf_ram.RAM[18][1] ;
 wire \rf_ram.RAM[18][20] ;
 wire \rf_ram.RAM[18][21] ;
 wire \rf_ram.RAM[18][22] ;
 wire \rf_ram.RAM[18][23] ;
 wire \rf_ram.RAM[18][24] ;
 wire \rf_ram.RAM[18][25] ;
 wire \rf_ram.RAM[18][26] ;
 wire \rf_ram.RAM[18][27] ;
 wire \rf_ram.RAM[18][28] ;
 wire \rf_ram.RAM[18][29] ;
 wire \rf_ram.RAM[18][2] ;
 wire \rf_ram.RAM[18][30] ;
 wire \rf_ram.RAM[18][31] ;
 wire \rf_ram.RAM[18][3] ;
 wire \rf_ram.RAM[18][4] ;
 wire \rf_ram.RAM[18][5] ;
 wire \rf_ram.RAM[18][6] ;
 wire \rf_ram.RAM[18][7] ;
 wire \rf_ram.RAM[18][8] ;
 wire \rf_ram.RAM[18][9] ;
 wire \rf_ram.RAM[19][0] ;
 wire \rf_ram.RAM[19][10] ;
 wire \rf_ram.RAM[19][11] ;
 wire \rf_ram.RAM[19][12] ;
 wire \rf_ram.RAM[19][13] ;
 wire \rf_ram.RAM[19][14] ;
 wire \rf_ram.RAM[19][15] ;
 wire \rf_ram.RAM[19][16] ;
 wire \rf_ram.RAM[19][17] ;
 wire \rf_ram.RAM[19][18] ;
 wire \rf_ram.RAM[19][19] ;
 wire \rf_ram.RAM[19][1] ;
 wire \rf_ram.RAM[19][20] ;
 wire \rf_ram.RAM[19][21] ;
 wire \rf_ram.RAM[19][22] ;
 wire \rf_ram.RAM[19][23] ;
 wire \rf_ram.RAM[19][24] ;
 wire \rf_ram.RAM[19][25] ;
 wire \rf_ram.RAM[19][26] ;
 wire \rf_ram.RAM[19][27] ;
 wire \rf_ram.RAM[19][28] ;
 wire \rf_ram.RAM[19][29] ;
 wire \rf_ram.RAM[19][2] ;
 wire \rf_ram.RAM[19][30] ;
 wire \rf_ram.RAM[19][31] ;
 wire \rf_ram.RAM[19][3] ;
 wire \rf_ram.RAM[19][4] ;
 wire \rf_ram.RAM[19][5] ;
 wire \rf_ram.RAM[19][6] ;
 wire \rf_ram.RAM[19][7] ;
 wire \rf_ram.RAM[19][8] ;
 wire \rf_ram.RAM[19][9] ;
 wire \rf_ram.RAM[1][0] ;
 wire \rf_ram.RAM[1][10] ;
 wire \rf_ram.RAM[1][11] ;
 wire \rf_ram.RAM[1][12] ;
 wire \rf_ram.RAM[1][13] ;
 wire \rf_ram.RAM[1][14] ;
 wire \rf_ram.RAM[1][15] ;
 wire \rf_ram.RAM[1][16] ;
 wire \rf_ram.RAM[1][17] ;
 wire \rf_ram.RAM[1][18] ;
 wire \rf_ram.RAM[1][19] ;
 wire \rf_ram.RAM[1][1] ;
 wire \rf_ram.RAM[1][20] ;
 wire \rf_ram.RAM[1][21] ;
 wire \rf_ram.RAM[1][22] ;
 wire \rf_ram.RAM[1][23] ;
 wire \rf_ram.RAM[1][24] ;
 wire \rf_ram.RAM[1][25] ;
 wire \rf_ram.RAM[1][26] ;
 wire \rf_ram.RAM[1][27] ;
 wire \rf_ram.RAM[1][28] ;
 wire \rf_ram.RAM[1][29] ;
 wire \rf_ram.RAM[1][2] ;
 wire \rf_ram.RAM[1][30] ;
 wire \rf_ram.RAM[1][31] ;
 wire \rf_ram.RAM[1][3] ;
 wire \rf_ram.RAM[1][4] ;
 wire \rf_ram.RAM[1][5] ;
 wire \rf_ram.RAM[1][6] ;
 wire \rf_ram.RAM[1][7] ;
 wire \rf_ram.RAM[1][8] ;
 wire \rf_ram.RAM[1][9] ;
 wire \rf_ram.RAM[20][0] ;
 wire \rf_ram.RAM[20][10] ;
 wire \rf_ram.RAM[20][11] ;
 wire \rf_ram.RAM[20][12] ;
 wire \rf_ram.RAM[20][13] ;
 wire \rf_ram.RAM[20][14] ;
 wire \rf_ram.RAM[20][15] ;
 wire \rf_ram.RAM[20][16] ;
 wire \rf_ram.RAM[20][17] ;
 wire \rf_ram.RAM[20][18] ;
 wire \rf_ram.RAM[20][19] ;
 wire \rf_ram.RAM[20][1] ;
 wire \rf_ram.RAM[20][20] ;
 wire \rf_ram.RAM[20][21] ;
 wire \rf_ram.RAM[20][22] ;
 wire \rf_ram.RAM[20][23] ;
 wire \rf_ram.RAM[20][24] ;
 wire \rf_ram.RAM[20][25] ;
 wire \rf_ram.RAM[20][26] ;
 wire \rf_ram.RAM[20][27] ;
 wire \rf_ram.RAM[20][28] ;
 wire \rf_ram.RAM[20][29] ;
 wire \rf_ram.RAM[20][2] ;
 wire \rf_ram.RAM[20][30] ;
 wire \rf_ram.RAM[20][31] ;
 wire \rf_ram.RAM[20][3] ;
 wire \rf_ram.RAM[20][4] ;
 wire \rf_ram.RAM[20][5] ;
 wire \rf_ram.RAM[20][6] ;
 wire \rf_ram.RAM[20][7] ;
 wire \rf_ram.RAM[20][8] ;
 wire \rf_ram.RAM[20][9] ;
 wire \rf_ram.RAM[21][0] ;
 wire \rf_ram.RAM[21][10] ;
 wire \rf_ram.RAM[21][11] ;
 wire \rf_ram.RAM[21][12] ;
 wire \rf_ram.RAM[21][13] ;
 wire \rf_ram.RAM[21][14] ;
 wire \rf_ram.RAM[21][15] ;
 wire \rf_ram.RAM[21][16] ;
 wire \rf_ram.RAM[21][17] ;
 wire \rf_ram.RAM[21][18] ;
 wire \rf_ram.RAM[21][19] ;
 wire \rf_ram.RAM[21][1] ;
 wire \rf_ram.RAM[21][20] ;
 wire \rf_ram.RAM[21][21] ;
 wire \rf_ram.RAM[21][22] ;
 wire \rf_ram.RAM[21][23] ;
 wire \rf_ram.RAM[21][24] ;
 wire \rf_ram.RAM[21][25] ;
 wire \rf_ram.RAM[21][26] ;
 wire \rf_ram.RAM[21][27] ;
 wire \rf_ram.RAM[21][28] ;
 wire \rf_ram.RAM[21][29] ;
 wire \rf_ram.RAM[21][2] ;
 wire \rf_ram.RAM[21][30] ;
 wire \rf_ram.RAM[21][31] ;
 wire \rf_ram.RAM[21][3] ;
 wire \rf_ram.RAM[21][4] ;
 wire \rf_ram.RAM[21][5] ;
 wire \rf_ram.RAM[21][6] ;
 wire \rf_ram.RAM[21][7] ;
 wire \rf_ram.RAM[21][8] ;
 wire \rf_ram.RAM[21][9] ;
 wire \rf_ram.RAM[22][0] ;
 wire \rf_ram.RAM[22][10] ;
 wire \rf_ram.RAM[22][11] ;
 wire \rf_ram.RAM[22][12] ;
 wire \rf_ram.RAM[22][13] ;
 wire \rf_ram.RAM[22][14] ;
 wire \rf_ram.RAM[22][15] ;
 wire \rf_ram.RAM[22][16] ;
 wire \rf_ram.RAM[22][17] ;
 wire \rf_ram.RAM[22][18] ;
 wire \rf_ram.RAM[22][19] ;
 wire \rf_ram.RAM[22][1] ;
 wire \rf_ram.RAM[22][20] ;
 wire \rf_ram.RAM[22][21] ;
 wire \rf_ram.RAM[22][22] ;
 wire \rf_ram.RAM[22][23] ;
 wire \rf_ram.RAM[22][24] ;
 wire \rf_ram.RAM[22][25] ;
 wire \rf_ram.RAM[22][26] ;
 wire \rf_ram.RAM[22][27] ;
 wire \rf_ram.RAM[22][28] ;
 wire \rf_ram.RAM[22][29] ;
 wire \rf_ram.RAM[22][2] ;
 wire \rf_ram.RAM[22][30] ;
 wire \rf_ram.RAM[22][31] ;
 wire \rf_ram.RAM[22][3] ;
 wire \rf_ram.RAM[22][4] ;
 wire \rf_ram.RAM[22][5] ;
 wire \rf_ram.RAM[22][6] ;
 wire \rf_ram.RAM[22][7] ;
 wire \rf_ram.RAM[22][8] ;
 wire \rf_ram.RAM[22][9] ;
 wire \rf_ram.RAM[23][0] ;
 wire \rf_ram.RAM[23][10] ;
 wire \rf_ram.RAM[23][11] ;
 wire \rf_ram.RAM[23][12] ;
 wire \rf_ram.RAM[23][13] ;
 wire \rf_ram.RAM[23][14] ;
 wire \rf_ram.RAM[23][15] ;
 wire \rf_ram.RAM[23][16] ;
 wire \rf_ram.RAM[23][17] ;
 wire \rf_ram.RAM[23][18] ;
 wire \rf_ram.RAM[23][19] ;
 wire \rf_ram.RAM[23][1] ;
 wire \rf_ram.RAM[23][20] ;
 wire \rf_ram.RAM[23][21] ;
 wire \rf_ram.RAM[23][22] ;
 wire \rf_ram.RAM[23][23] ;
 wire \rf_ram.RAM[23][24] ;
 wire \rf_ram.RAM[23][25] ;
 wire \rf_ram.RAM[23][26] ;
 wire \rf_ram.RAM[23][27] ;
 wire \rf_ram.RAM[23][28] ;
 wire \rf_ram.RAM[23][29] ;
 wire \rf_ram.RAM[23][2] ;
 wire \rf_ram.RAM[23][30] ;
 wire \rf_ram.RAM[23][31] ;
 wire \rf_ram.RAM[23][3] ;
 wire \rf_ram.RAM[23][4] ;
 wire \rf_ram.RAM[23][5] ;
 wire \rf_ram.RAM[23][6] ;
 wire \rf_ram.RAM[23][7] ;
 wire \rf_ram.RAM[23][8] ;
 wire \rf_ram.RAM[23][9] ;
 wire \rf_ram.RAM[24][0] ;
 wire \rf_ram.RAM[24][10] ;
 wire \rf_ram.RAM[24][11] ;
 wire \rf_ram.RAM[24][12] ;
 wire \rf_ram.RAM[24][13] ;
 wire \rf_ram.RAM[24][14] ;
 wire \rf_ram.RAM[24][15] ;
 wire \rf_ram.RAM[24][16] ;
 wire \rf_ram.RAM[24][17] ;
 wire \rf_ram.RAM[24][18] ;
 wire \rf_ram.RAM[24][19] ;
 wire \rf_ram.RAM[24][1] ;
 wire \rf_ram.RAM[24][20] ;
 wire \rf_ram.RAM[24][21] ;
 wire \rf_ram.RAM[24][22] ;
 wire \rf_ram.RAM[24][23] ;
 wire \rf_ram.RAM[24][24] ;
 wire \rf_ram.RAM[24][25] ;
 wire \rf_ram.RAM[24][26] ;
 wire \rf_ram.RAM[24][27] ;
 wire \rf_ram.RAM[24][28] ;
 wire \rf_ram.RAM[24][29] ;
 wire \rf_ram.RAM[24][2] ;
 wire \rf_ram.RAM[24][30] ;
 wire \rf_ram.RAM[24][31] ;
 wire \rf_ram.RAM[24][3] ;
 wire \rf_ram.RAM[24][4] ;
 wire \rf_ram.RAM[24][5] ;
 wire \rf_ram.RAM[24][6] ;
 wire \rf_ram.RAM[24][7] ;
 wire \rf_ram.RAM[24][8] ;
 wire \rf_ram.RAM[24][9] ;
 wire \rf_ram.RAM[25][0] ;
 wire \rf_ram.RAM[25][10] ;
 wire \rf_ram.RAM[25][11] ;
 wire \rf_ram.RAM[25][12] ;
 wire \rf_ram.RAM[25][13] ;
 wire \rf_ram.RAM[25][14] ;
 wire \rf_ram.RAM[25][15] ;
 wire \rf_ram.RAM[25][16] ;
 wire \rf_ram.RAM[25][17] ;
 wire \rf_ram.RAM[25][18] ;
 wire \rf_ram.RAM[25][19] ;
 wire \rf_ram.RAM[25][1] ;
 wire \rf_ram.RAM[25][20] ;
 wire \rf_ram.RAM[25][21] ;
 wire \rf_ram.RAM[25][22] ;
 wire \rf_ram.RAM[25][23] ;
 wire \rf_ram.RAM[25][24] ;
 wire \rf_ram.RAM[25][25] ;
 wire \rf_ram.RAM[25][26] ;
 wire \rf_ram.RAM[25][27] ;
 wire \rf_ram.RAM[25][28] ;
 wire \rf_ram.RAM[25][29] ;
 wire \rf_ram.RAM[25][2] ;
 wire \rf_ram.RAM[25][30] ;
 wire \rf_ram.RAM[25][31] ;
 wire \rf_ram.RAM[25][3] ;
 wire \rf_ram.RAM[25][4] ;
 wire \rf_ram.RAM[25][5] ;
 wire \rf_ram.RAM[25][6] ;
 wire \rf_ram.RAM[25][7] ;
 wire \rf_ram.RAM[25][8] ;
 wire \rf_ram.RAM[25][9] ;
 wire \rf_ram.RAM[26][0] ;
 wire \rf_ram.RAM[26][10] ;
 wire \rf_ram.RAM[26][11] ;
 wire \rf_ram.RAM[26][12] ;
 wire \rf_ram.RAM[26][13] ;
 wire \rf_ram.RAM[26][14] ;
 wire \rf_ram.RAM[26][15] ;
 wire \rf_ram.RAM[26][16] ;
 wire \rf_ram.RAM[26][17] ;
 wire \rf_ram.RAM[26][18] ;
 wire \rf_ram.RAM[26][19] ;
 wire \rf_ram.RAM[26][1] ;
 wire \rf_ram.RAM[26][20] ;
 wire \rf_ram.RAM[26][21] ;
 wire \rf_ram.RAM[26][22] ;
 wire \rf_ram.RAM[26][23] ;
 wire \rf_ram.RAM[26][24] ;
 wire \rf_ram.RAM[26][25] ;
 wire \rf_ram.RAM[26][26] ;
 wire \rf_ram.RAM[26][27] ;
 wire \rf_ram.RAM[26][28] ;
 wire \rf_ram.RAM[26][29] ;
 wire \rf_ram.RAM[26][2] ;
 wire \rf_ram.RAM[26][30] ;
 wire \rf_ram.RAM[26][31] ;
 wire \rf_ram.RAM[26][3] ;
 wire \rf_ram.RAM[26][4] ;
 wire \rf_ram.RAM[26][5] ;
 wire \rf_ram.RAM[26][6] ;
 wire \rf_ram.RAM[26][7] ;
 wire \rf_ram.RAM[26][8] ;
 wire \rf_ram.RAM[26][9] ;
 wire \rf_ram.RAM[27][0] ;
 wire \rf_ram.RAM[27][10] ;
 wire \rf_ram.RAM[27][11] ;
 wire \rf_ram.RAM[27][12] ;
 wire \rf_ram.RAM[27][13] ;
 wire \rf_ram.RAM[27][14] ;
 wire \rf_ram.RAM[27][15] ;
 wire \rf_ram.RAM[27][16] ;
 wire \rf_ram.RAM[27][17] ;
 wire \rf_ram.RAM[27][18] ;
 wire \rf_ram.RAM[27][19] ;
 wire \rf_ram.RAM[27][1] ;
 wire \rf_ram.RAM[27][20] ;
 wire \rf_ram.RAM[27][21] ;
 wire \rf_ram.RAM[27][22] ;
 wire \rf_ram.RAM[27][23] ;
 wire \rf_ram.RAM[27][24] ;
 wire \rf_ram.RAM[27][25] ;
 wire \rf_ram.RAM[27][26] ;
 wire \rf_ram.RAM[27][27] ;
 wire \rf_ram.RAM[27][28] ;
 wire \rf_ram.RAM[27][29] ;
 wire \rf_ram.RAM[27][2] ;
 wire \rf_ram.RAM[27][30] ;
 wire \rf_ram.RAM[27][31] ;
 wire \rf_ram.RAM[27][3] ;
 wire \rf_ram.RAM[27][4] ;
 wire \rf_ram.RAM[27][5] ;
 wire \rf_ram.RAM[27][6] ;
 wire \rf_ram.RAM[27][7] ;
 wire \rf_ram.RAM[27][8] ;
 wire \rf_ram.RAM[27][9] ;
 wire \rf_ram.RAM[28][0] ;
 wire \rf_ram.RAM[28][10] ;
 wire \rf_ram.RAM[28][11] ;
 wire \rf_ram.RAM[28][12] ;
 wire \rf_ram.RAM[28][13] ;
 wire \rf_ram.RAM[28][14] ;
 wire \rf_ram.RAM[28][15] ;
 wire \rf_ram.RAM[28][16] ;
 wire \rf_ram.RAM[28][17] ;
 wire \rf_ram.RAM[28][18] ;
 wire \rf_ram.RAM[28][19] ;
 wire \rf_ram.RAM[28][1] ;
 wire \rf_ram.RAM[28][20] ;
 wire \rf_ram.RAM[28][21] ;
 wire \rf_ram.RAM[28][22] ;
 wire \rf_ram.RAM[28][23] ;
 wire \rf_ram.RAM[28][24] ;
 wire \rf_ram.RAM[28][25] ;
 wire \rf_ram.RAM[28][26] ;
 wire \rf_ram.RAM[28][27] ;
 wire \rf_ram.RAM[28][28] ;
 wire \rf_ram.RAM[28][29] ;
 wire \rf_ram.RAM[28][2] ;
 wire \rf_ram.RAM[28][30] ;
 wire \rf_ram.RAM[28][31] ;
 wire \rf_ram.RAM[28][3] ;
 wire \rf_ram.RAM[28][4] ;
 wire \rf_ram.RAM[28][5] ;
 wire \rf_ram.RAM[28][6] ;
 wire \rf_ram.RAM[28][7] ;
 wire \rf_ram.RAM[28][8] ;
 wire \rf_ram.RAM[28][9] ;
 wire \rf_ram.RAM[29][0] ;
 wire \rf_ram.RAM[29][10] ;
 wire \rf_ram.RAM[29][11] ;
 wire \rf_ram.RAM[29][12] ;
 wire \rf_ram.RAM[29][13] ;
 wire \rf_ram.RAM[29][14] ;
 wire \rf_ram.RAM[29][15] ;
 wire \rf_ram.RAM[29][16] ;
 wire \rf_ram.RAM[29][17] ;
 wire \rf_ram.RAM[29][18] ;
 wire \rf_ram.RAM[29][19] ;
 wire \rf_ram.RAM[29][1] ;
 wire \rf_ram.RAM[29][20] ;
 wire \rf_ram.RAM[29][21] ;
 wire \rf_ram.RAM[29][22] ;
 wire \rf_ram.RAM[29][23] ;
 wire \rf_ram.RAM[29][24] ;
 wire \rf_ram.RAM[29][25] ;
 wire \rf_ram.RAM[29][26] ;
 wire \rf_ram.RAM[29][27] ;
 wire \rf_ram.RAM[29][28] ;
 wire \rf_ram.RAM[29][29] ;
 wire \rf_ram.RAM[29][2] ;
 wire \rf_ram.RAM[29][30] ;
 wire \rf_ram.RAM[29][31] ;
 wire \rf_ram.RAM[29][3] ;
 wire \rf_ram.RAM[29][4] ;
 wire \rf_ram.RAM[29][5] ;
 wire \rf_ram.RAM[29][6] ;
 wire \rf_ram.RAM[29][7] ;
 wire \rf_ram.RAM[29][8] ;
 wire \rf_ram.RAM[29][9] ;
 wire \rf_ram.RAM[2][0] ;
 wire \rf_ram.RAM[2][10] ;
 wire \rf_ram.RAM[2][11] ;
 wire \rf_ram.RAM[2][12] ;
 wire \rf_ram.RAM[2][13] ;
 wire \rf_ram.RAM[2][14] ;
 wire \rf_ram.RAM[2][15] ;
 wire \rf_ram.RAM[2][16] ;
 wire \rf_ram.RAM[2][17] ;
 wire \rf_ram.RAM[2][18] ;
 wire \rf_ram.RAM[2][19] ;
 wire \rf_ram.RAM[2][1] ;
 wire \rf_ram.RAM[2][20] ;
 wire \rf_ram.RAM[2][21] ;
 wire \rf_ram.RAM[2][22] ;
 wire \rf_ram.RAM[2][23] ;
 wire \rf_ram.RAM[2][24] ;
 wire \rf_ram.RAM[2][25] ;
 wire \rf_ram.RAM[2][26] ;
 wire \rf_ram.RAM[2][27] ;
 wire \rf_ram.RAM[2][28] ;
 wire \rf_ram.RAM[2][29] ;
 wire \rf_ram.RAM[2][2] ;
 wire \rf_ram.RAM[2][30] ;
 wire \rf_ram.RAM[2][31] ;
 wire \rf_ram.RAM[2][3] ;
 wire \rf_ram.RAM[2][4] ;
 wire \rf_ram.RAM[2][5] ;
 wire \rf_ram.RAM[2][6] ;
 wire \rf_ram.RAM[2][7] ;
 wire \rf_ram.RAM[2][8] ;
 wire \rf_ram.RAM[2][9] ;
 wire \rf_ram.RAM[30][0] ;
 wire \rf_ram.RAM[30][10] ;
 wire \rf_ram.RAM[30][11] ;
 wire \rf_ram.RAM[30][12] ;
 wire \rf_ram.RAM[30][13] ;
 wire \rf_ram.RAM[30][14] ;
 wire \rf_ram.RAM[30][15] ;
 wire \rf_ram.RAM[30][16] ;
 wire \rf_ram.RAM[30][17] ;
 wire \rf_ram.RAM[30][18] ;
 wire \rf_ram.RAM[30][19] ;
 wire \rf_ram.RAM[30][1] ;
 wire \rf_ram.RAM[30][20] ;
 wire \rf_ram.RAM[30][21] ;
 wire \rf_ram.RAM[30][22] ;
 wire \rf_ram.RAM[30][23] ;
 wire \rf_ram.RAM[30][24] ;
 wire \rf_ram.RAM[30][25] ;
 wire \rf_ram.RAM[30][26] ;
 wire \rf_ram.RAM[30][27] ;
 wire \rf_ram.RAM[30][28] ;
 wire \rf_ram.RAM[30][29] ;
 wire \rf_ram.RAM[30][2] ;
 wire \rf_ram.RAM[30][30] ;
 wire \rf_ram.RAM[30][31] ;
 wire \rf_ram.RAM[30][3] ;
 wire \rf_ram.RAM[30][4] ;
 wire \rf_ram.RAM[30][5] ;
 wire \rf_ram.RAM[30][6] ;
 wire \rf_ram.RAM[30][7] ;
 wire \rf_ram.RAM[30][8] ;
 wire \rf_ram.RAM[30][9] ;
 wire \rf_ram.RAM[31][0] ;
 wire \rf_ram.RAM[31][10] ;
 wire \rf_ram.RAM[31][11] ;
 wire \rf_ram.RAM[31][12] ;
 wire \rf_ram.RAM[31][13] ;
 wire \rf_ram.RAM[31][14] ;
 wire \rf_ram.RAM[31][15] ;
 wire \rf_ram.RAM[31][16] ;
 wire \rf_ram.RAM[31][17] ;
 wire \rf_ram.RAM[31][18] ;
 wire \rf_ram.RAM[31][19] ;
 wire \rf_ram.RAM[31][1] ;
 wire \rf_ram.RAM[31][20] ;
 wire \rf_ram.RAM[31][21] ;
 wire \rf_ram.RAM[31][22] ;
 wire \rf_ram.RAM[31][23] ;
 wire \rf_ram.RAM[31][24] ;
 wire \rf_ram.RAM[31][25] ;
 wire \rf_ram.RAM[31][26] ;
 wire \rf_ram.RAM[31][27] ;
 wire \rf_ram.RAM[31][28] ;
 wire \rf_ram.RAM[31][29] ;
 wire \rf_ram.RAM[31][2] ;
 wire \rf_ram.RAM[31][30] ;
 wire \rf_ram.RAM[31][31] ;
 wire \rf_ram.RAM[31][3] ;
 wire \rf_ram.RAM[31][4] ;
 wire \rf_ram.RAM[31][5] ;
 wire \rf_ram.RAM[31][6] ;
 wire \rf_ram.RAM[31][7] ;
 wire \rf_ram.RAM[31][8] ;
 wire \rf_ram.RAM[31][9] ;
 wire \rf_ram.RAM[3][0] ;
 wire \rf_ram.RAM[3][10] ;
 wire \rf_ram.RAM[3][11] ;
 wire \rf_ram.RAM[3][12] ;
 wire \rf_ram.RAM[3][13] ;
 wire \rf_ram.RAM[3][14] ;
 wire \rf_ram.RAM[3][15] ;
 wire \rf_ram.RAM[3][16] ;
 wire \rf_ram.RAM[3][17] ;
 wire \rf_ram.RAM[3][18] ;
 wire \rf_ram.RAM[3][19] ;
 wire \rf_ram.RAM[3][1] ;
 wire \rf_ram.RAM[3][20] ;
 wire \rf_ram.RAM[3][21] ;
 wire \rf_ram.RAM[3][22] ;
 wire \rf_ram.RAM[3][23] ;
 wire \rf_ram.RAM[3][24] ;
 wire \rf_ram.RAM[3][25] ;
 wire \rf_ram.RAM[3][26] ;
 wire \rf_ram.RAM[3][27] ;
 wire \rf_ram.RAM[3][28] ;
 wire \rf_ram.RAM[3][29] ;
 wire \rf_ram.RAM[3][2] ;
 wire \rf_ram.RAM[3][30] ;
 wire \rf_ram.RAM[3][31] ;
 wire \rf_ram.RAM[3][3] ;
 wire \rf_ram.RAM[3][4] ;
 wire \rf_ram.RAM[3][5] ;
 wire \rf_ram.RAM[3][6] ;
 wire \rf_ram.RAM[3][7] ;
 wire \rf_ram.RAM[3][8] ;
 wire \rf_ram.RAM[3][9] ;
 wire \rf_ram.RAM[4][0] ;
 wire \rf_ram.RAM[4][10] ;
 wire \rf_ram.RAM[4][11] ;
 wire \rf_ram.RAM[4][12] ;
 wire \rf_ram.RAM[4][13] ;
 wire \rf_ram.RAM[4][14] ;
 wire \rf_ram.RAM[4][15] ;
 wire \rf_ram.RAM[4][16] ;
 wire \rf_ram.RAM[4][17] ;
 wire \rf_ram.RAM[4][18] ;
 wire \rf_ram.RAM[4][19] ;
 wire \rf_ram.RAM[4][1] ;
 wire \rf_ram.RAM[4][20] ;
 wire \rf_ram.RAM[4][21] ;
 wire \rf_ram.RAM[4][22] ;
 wire \rf_ram.RAM[4][23] ;
 wire \rf_ram.RAM[4][24] ;
 wire \rf_ram.RAM[4][25] ;
 wire \rf_ram.RAM[4][26] ;
 wire \rf_ram.RAM[4][27] ;
 wire \rf_ram.RAM[4][28] ;
 wire \rf_ram.RAM[4][29] ;
 wire \rf_ram.RAM[4][2] ;
 wire \rf_ram.RAM[4][30] ;
 wire \rf_ram.RAM[4][31] ;
 wire \rf_ram.RAM[4][3] ;
 wire \rf_ram.RAM[4][4] ;
 wire \rf_ram.RAM[4][5] ;
 wire \rf_ram.RAM[4][6] ;
 wire \rf_ram.RAM[4][7] ;
 wire \rf_ram.RAM[4][8] ;
 wire \rf_ram.RAM[4][9] ;
 wire \rf_ram.RAM[5][0] ;
 wire \rf_ram.RAM[5][10] ;
 wire \rf_ram.RAM[5][11] ;
 wire \rf_ram.RAM[5][12] ;
 wire \rf_ram.RAM[5][13] ;
 wire \rf_ram.RAM[5][14] ;
 wire \rf_ram.RAM[5][15] ;
 wire \rf_ram.RAM[5][16] ;
 wire \rf_ram.RAM[5][17] ;
 wire \rf_ram.RAM[5][18] ;
 wire \rf_ram.RAM[5][19] ;
 wire \rf_ram.RAM[5][1] ;
 wire \rf_ram.RAM[5][20] ;
 wire \rf_ram.RAM[5][21] ;
 wire \rf_ram.RAM[5][22] ;
 wire \rf_ram.RAM[5][23] ;
 wire \rf_ram.RAM[5][24] ;
 wire \rf_ram.RAM[5][25] ;
 wire \rf_ram.RAM[5][26] ;
 wire \rf_ram.RAM[5][27] ;
 wire \rf_ram.RAM[5][28] ;
 wire \rf_ram.RAM[5][29] ;
 wire \rf_ram.RAM[5][2] ;
 wire \rf_ram.RAM[5][30] ;
 wire \rf_ram.RAM[5][31] ;
 wire \rf_ram.RAM[5][3] ;
 wire \rf_ram.RAM[5][4] ;
 wire \rf_ram.RAM[5][5] ;
 wire \rf_ram.RAM[5][6] ;
 wire \rf_ram.RAM[5][7] ;
 wire \rf_ram.RAM[5][8] ;
 wire \rf_ram.RAM[5][9] ;
 wire \rf_ram.RAM[6][0] ;
 wire \rf_ram.RAM[6][10] ;
 wire \rf_ram.RAM[6][11] ;
 wire \rf_ram.RAM[6][12] ;
 wire \rf_ram.RAM[6][13] ;
 wire \rf_ram.RAM[6][14] ;
 wire \rf_ram.RAM[6][15] ;
 wire \rf_ram.RAM[6][16] ;
 wire \rf_ram.RAM[6][17] ;
 wire \rf_ram.RAM[6][18] ;
 wire \rf_ram.RAM[6][19] ;
 wire \rf_ram.RAM[6][1] ;
 wire \rf_ram.RAM[6][20] ;
 wire \rf_ram.RAM[6][21] ;
 wire \rf_ram.RAM[6][22] ;
 wire \rf_ram.RAM[6][23] ;
 wire \rf_ram.RAM[6][24] ;
 wire \rf_ram.RAM[6][25] ;
 wire \rf_ram.RAM[6][26] ;
 wire \rf_ram.RAM[6][27] ;
 wire \rf_ram.RAM[6][28] ;
 wire \rf_ram.RAM[6][29] ;
 wire \rf_ram.RAM[6][2] ;
 wire \rf_ram.RAM[6][30] ;
 wire \rf_ram.RAM[6][31] ;
 wire \rf_ram.RAM[6][3] ;
 wire \rf_ram.RAM[6][4] ;
 wire \rf_ram.RAM[6][5] ;
 wire \rf_ram.RAM[6][6] ;
 wire \rf_ram.RAM[6][7] ;
 wire \rf_ram.RAM[6][8] ;
 wire \rf_ram.RAM[6][9] ;
 wire \rf_ram.RAM[7][0] ;
 wire \rf_ram.RAM[7][10] ;
 wire \rf_ram.RAM[7][11] ;
 wire \rf_ram.RAM[7][12] ;
 wire \rf_ram.RAM[7][13] ;
 wire \rf_ram.RAM[7][14] ;
 wire \rf_ram.RAM[7][15] ;
 wire \rf_ram.RAM[7][16] ;
 wire \rf_ram.RAM[7][17] ;
 wire \rf_ram.RAM[7][18] ;
 wire \rf_ram.RAM[7][19] ;
 wire \rf_ram.RAM[7][1] ;
 wire \rf_ram.RAM[7][20] ;
 wire \rf_ram.RAM[7][21] ;
 wire \rf_ram.RAM[7][22] ;
 wire \rf_ram.RAM[7][23] ;
 wire \rf_ram.RAM[7][24] ;
 wire \rf_ram.RAM[7][25] ;
 wire \rf_ram.RAM[7][26] ;
 wire \rf_ram.RAM[7][27] ;
 wire \rf_ram.RAM[7][28] ;
 wire \rf_ram.RAM[7][29] ;
 wire \rf_ram.RAM[7][2] ;
 wire \rf_ram.RAM[7][30] ;
 wire \rf_ram.RAM[7][31] ;
 wire \rf_ram.RAM[7][3] ;
 wire \rf_ram.RAM[7][4] ;
 wire \rf_ram.RAM[7][5] ;
 wire \rf_ram.RAM[7][6] ;
 wire \rf_ram.RAM[7][7] ;
 wire \rf_ram.RAM[7][8] ;
 wire \rf_ram.RAM[7][9] ;
 wire \rf_ram.RAM[8][0] ;
 wire \rf_ram.RAM[8][10] ;
 wire \rf_ram.RAM[8][11] ;
 wire \rf_ram.RAM[8][12] ;
 wire \rf_ram.RAM[8][13] ;
 wire \rf_ram.RAM[8][14] ;
 wire \rf_ram.RAM[8][15] ;
 wire \rf_ram.RAM[8][16] ;
 wire \rf_ram.RAM[8][17] ;
 wire \rf_ram.RAM[8][18] ;
 wire \rf_ram.RAM[8][19] ;
 wire \rf_ram.RAM[8][1] ;
 wire \rf_ram.RAM[8][20] ;
 wire \rf_ram.RAM[8][21] ;
 wire \rf_ram.RAM[8][22] ;
 wire \rf_ram.RAM[8][23] ;
 wire \rf_ram.RAM[8][24] ;
 wire \rf_ram.RAM[8][25] ;
 wire \rf_ram.RAM[8][26] ;
 wire \rf_ram.RAM[8][27] ;
 wire \rf_ram.RAM[8][28] ;
 wire \rf_ram.RAM[8][29] ;
 wire \rf_ram.RAM[8][2] ;
 wire \rf_ram.RAM[8][30] ;
 wire \rf_ram.RAM[8][31] ;
 wire \rf_ram.RAM[8][3] ;
 wire \rf_ram.RAM[8][4] ;
 wire \rf_ram.RAM[8][5] ;
 wire \rf_ram.RAM[8][6] ;
 wire \rf_ram.RAM[8][7] ;
 wire \rf_ram.RAM[8][8] ;
 wire \rf_ram.RAM[8][9] ;
 wire \rf_ram.RAM[9][0] ;
 wire \rf_ram.RAM[9][10] ;
 wire \rf_ram.RAM[9][11] ;
 wire \rf_ram.RAM[9][12] ;
 wire \rf_ram.RAM[9][13] ;
 wire \rf_ram.RAM[9][14] ;
 wire \rf_ram.RAM[9][15] ;
 wire \rf_ram.RAM[9][16] ;
 wire \rf_ram.RAM[9][17] ;
 wire \rf_ram.RAM[9][18] ;
 wire \rf_ram.RAM[9][19] ;
 wire \rf_ram.RAM[9][1] ;
 wire \rf_ram.RAM[9][20] ;
 wire \rf_ram.RAM[9][21] ;
 wire \rf_ram.RAM[9][22] ;
 wire \rf_ram.RAM[9][23] ;
 wire \rf_ram.RAM[9][24] ;
 wire \rf_ram.RAM[9][25] ;
 wire \rf_ram.RAM[9][26] ;
 wire \rf_ram.RAM[9][27] ;
 wire \rf_ram.RAM[9][28] ;
 wire \rf_ram.RAM[9][29] ;
 wire \rf_ram.RAM[9][2] ;
 wire \rf_ram.RAM[9][30] ;
 wire \rf_ram.RAM[9][31] ;
 wire \rf_ram.RAM[9][3] ;
 wire \rf_ram.RAM[9][4] ;
 wire \rf_ram.RAM[9][5] ;
 wire \rf_ram.RAM[9][6] ;
 wire \rf_ram.RAM[9][7] ;
 wire \rf_ram.RAM[9][8] ;
 wire \rf_ram.RAM[9][9] ;
 wire net1375;
 wire net1376;
 wire net8;
 wire net1377;
 wire net1378;
 wire net1379;
 wire net9;
 wire net10;
 wire net11;
 wire net1380;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net1749;
 wire net1750;
 wire net1751;
 wire net1752;
 wire net1753;
 wire net1754;
 wire net1755;
 wire net1756;
 wire net1757;
 wire net1758;
 wire net1759;
 wire net1760;
 wire net1761;
 wire net1762;
 wire net1763;
 wire net1764;
 wire net1765;
 wire net1766;
 wire net1767;
 wire net1768;
 wire net1769;
 wire net1770;
 wire net1771;
 wire net1772;
 wire net1773;
 wire net1774;
 wire net1775;
 wire net1776;
 wire net1777;
 wire net1778;
 wire net1779;
 wire net1780;
 wire net1781;
 wire net1782;
 wire net1783;
 wire net1784;
 wire net1785;
 wire net1786;
 wire net1787;
 wire net1788;
 wire net1789;
 wire net1790;
 wire net1791;
 wire net1792;
 wire net1793;
 wire net1794;
 wire net1795;
 wire net1796;
 wire net1797;
 wire net1798;
 wire net1799;
 wire net1800;
 wire net1801;
 wire net1802;
 wire net1803;
 wire net1804;
 wire net1805;
 wire net1806;
 wire net1807;
 wire net1808;
 wire net1809;
 wire net1810;
 wire net1811;
 wire net1812;
 wire net1813;
 wire net1814;
 wire net1815;
 wire net1816;
 wire net1817;
 wire net1818;
 wire net1819;
 wire net1820;
 wire net1821;
 wire net1822;
 wire net1823;
 wire net1824;
 wire net1825;
 wire net1826;
 wire net1827;
 wire net1828;
 wire net1829;
 wire net1830;
 wire net1831;
 wire net1832;
 wire net1833;
 wire net1834;
 wire net1835;
 wire net1836;
 wire net1837;
 wire net1838;
 wire net1839;
 wire net1840;
 wire net1841;
 wire net1842;
 wire net1843;
 wire net1844;
 wire net1845;
 wire net1846;
 wire net1847;
 wire net1848;
 wire net1849;
 wire net1850;
 wire net1851;
 wire net1852;
 wire net1853;
 wire net1854;
 wire net1855;
 wire net1856;
 wire net1857;
 wire net1858;
 wire net1859;
 wire net1860;
 wire net1861;
 wire net1862;
 wire net1863;
 wire net1864;
 wire net1865;
 wire net1866;
 wire net1867;
 wire net1868;
 wire net1869;
 wire net1870;
 wire net1871;
 wire net1872;
 wire net1873;
 wire net1874;
 wire net1875;
 wire net1876;
 wire net1877;
 wire net1878;
 wire net1879;
 wire net1880;
 wire net1881;
 wire net1882;
 wire net1883;
 wire net1884;
 wire net1885;
 wire net1886;
 wire net1887;
 wire net1888;
 wire net1889;
 wire net1890;
 wire net1891;
 wire net1892;
 wire net1893;
 wire net1894;
 wire net1895;
 wire net1896;
 wire net1897;
 wire net1898;
 wire net1899;
 wire net1900;
 wire net1901;
 wire net1902;
 wire net1903;
 wire net1904;
 wire net1905;
 wire net1906;
 wire net1907;
 wire net1908;
 wire net1909;
 wire net1910;
 wire net1911;
 wire net1912;
 wire net1913;
 wire net1914;
 wire net1915;
 wire net1916;
 wire net1917;
 wire net1918;
 wire net1919;
 wire net1920;
 wire net1921;
 wire net1922;
 wire net1923;
 wire net1924;
 wire net1925;
 wire net1926;
 wire net1927;
 wire net1928;
 wire net1929;
 wire net1930;
 wire net1931;
 wire net1932;
 wire net1933;
 wire net1934;
 wire net1935;
 wire net1936;
 wire net1937;
 wire net1938;
 wire net1939;
 wire net1940;
 wire net1941;
 wire net1942;
 wire net1943;
 wire net1944;
 wire net1945;
 wire net1946;
 wire net1947;
 wire net1948;
 wire net1949;
 wire net1950;
 wire net1951;
 wire net1952;
 wire net1953;
 wire net1954;
 wire net1955;
 wire net1956;
 wire net1957;
 wire net1958;
 wire net1959;
 wire net1960;
 wire net1961;
 wire net1962;
 wire net1963;
 wire net1964;
 wire net1965;
 wire net1966;
 wire net1967;
 wire net1968;
 wire net1969;
 wire net1970;
 wire net1971;
 wire net1972;
 wire net1973;
 wire net1974;
 wire net1975;
 wire net1976;
 wire net1977;
 wire net1978;
 wire net1979;
 wire net1980;
 wire net1981;
 wire net1982;
 wire net1983;
 wire net1984;
 wire net1985;
 wire net1986;
 wire net1987;
 wire net1988;
 wire net1989;
 wire net1990;
 wire net1991;
 wire net1992;
 wire net1993;
 wire net1994;
 wire net1995;
 wire net1996;
 wire net1997;
 wire net1998;
 wire net1999;
 wire net2000;
 wire net2001;
 wire net2002;
 wire net2003;
 wire net2004;
 wire net2005;
 wire net2006;
 wire net2007;
 wire net2008;
 wire net2009;
 wire net2010;
 wire net2011;
 wire net2012;
 wire net2013;
 wire net2014;
 wire net2015;
 wire net2016;
 wire net2017;
 wire net2018;
 wire net2019;
 wire net2020;
 wire net2021;
 wire net2022;
 wire net2023;
 wire net2024;
 wire net2025;
 wire net2026;
 wire net2027;
 wire net2028;
 wire net2029;
 wire net2030;
 wire net2031;
 wire net2032;
 wire net2033;
 wire net2034;
 wire net2035;
 wire net2036;
 wire net2037;
 wire net2038;
 wire net2039;
 wire net2040;
 wire net2041;
 wire net2042;
 wire net2043;
 wire net2044;
 wire net2045;
 wire net2046;
 wire net2047;
 wire net2048;
 wire net2049;
 wire net2050;
 wire net2051;
 wire net2052;
 wire net2053;
 wire net2054;
 wire net2055;
 wire net2056;
 wire net2057;
 wire net2058;
 wire net2059;
 wire net2060;
 wire net2061;
 wire net2062;
 wire net2063;
 wire net2064;
 wire net2065;
 wire net2066;
 wire net2067;
 wire net2068;
 wire net2069;
 wire net2070;
 wire net2071;
 wire net2072;
 wire net2073;
 wire net2074;
 wire net2075;
 wire net2076;
 wire net2077;
 wire net2078;
 wire net2079;
 wire net2080;
 wire net2081;
 wire net2082;
 wire net2083;
 wire net2084;
 wire net2085;
 wire net2086;
 wire net2087;
 wire net2088;
 wire net2089;
 wire net2090;
 wire net2091;
 wire net2092;
 wire net2093;
 wire net2094;
 wire net2095;
 wire net2096;
 wire net2097;
 wire net2098;
 wire net2099;
 wire net2100;
 wire net2101;
 wire net2102;
 wire net2103;
 wire net2104;
 wire net2105;
 wire net2106;
 wire net2107;
 wire net2108;
 wire net2109;
 wire net2110;
 wire net2111;
 wire net2112;
 wire net2113;
 wire net2114;
 wire net2115;
 wire net2116;
 wire net2117;
 wire net2118;
 wire net2119;
 wire net2120;
 wire net2121;
 wire net2122;
 wire net2123;
 wire net2124;
 wire net2125;
 wire net2126;
 wire net2127;
 wire net2128;
 wire net2129;
 wire net2130;
 wire net2131;
 wire net2132;
 wire net2133;
 wire net2134;
 wire net2135;
 wire net2136;
 wire net2137;
 wire net2138;
 wire net2139;
 wire net2140;
 wire net2141;
 wire net2142;
 wire net2143;
 wire net2144;
 wire net2145;
 wire net2146;
 wire net2147;
 wire net2148;
 wire net2149;
 wire net2150;
 wire net2151;
 wire net2152;
 wire net2153;
 wire net2154;
 wire net2155;
 wire net2156;
 wire net2157;
 wire net2158;
 wire net2159;
 wire net2160;
 wire net2161;
 wire net2162;
 wire net2163;
 wire net2164;
 wire net2165;
 wire net2166;
 wire net2167;
 wire net2168;
 wire net2169;
 wire net2170;
 wire net2171;
 wire net2172;
 wire net2173;
 wire net2174;
 wire net2175;
 wire net2176;
 wire net2177;
 wire net2178;
 wire net2179;
 wire net2180;
 wire net2181;
 wire net2182;
 wire net2183;
 wire net2184;
 wire net2185;
 wire net2186;
 wire net2187;
 wire net2188;
 wire net2189;
 wire net2190;
 wire net2191;
 wire net2192;
 wire net2193;
 wire net2194;
 wire net2195;
 wire net2196;
 wire net2197;
 wire net2198;
 wire net2199;
 wire net2200;
 wire net2201;
 wire net2202;
 wire net2203;
 wire net2204;
 wire net2205;
 wire net2206;
 wire net2207;
 wire net2208;
 wire net2209;
 wire net2210;
 wire net2211;
 wire net2212;
 wire net2213;
 wire net2214;
 wire net2215;
 wire net2216;
 wire net2217;
 wire net2218;
 wire net2219;
 wire net2220;
 wire net2221;
 wire net2222;
 wire net2223;
 wire net2224;
 wire net2225;
 wire net2226;
 wire net2227;
 wire net2228;
 wire net2229;
 wire net2230;
 wire net2231;
 wire net2232;
 wire net2233;
 wire net2234;
 wire net2235;
 wire net2236;
 wire net2237;
 wire net2238;
 wire net2239;
 wire net2240;
 wire net2241;
 wire net2242;
 wire net2243;
 wire net2244;
 wire net2245;
 wire net2246;
 wire net2247;
 wire net2248;
 wire net2249;
 wire net2250;
 wire net2251;
 wire net2252;
 wire net2253;
 wire net2254;
 wire net2255;
 wire net2256;
 wire net2257;
 wire net2258;
 wire net2259;
 wire net2260;
 wire net2261;
 wire net2262;
 wire net2263;
 wire net2264;
 wire net2265;
 wire net2266;
 wire net2267;
 wire net2268;
 wire net2269;
 wire net2270;
 wire net2271;
 wire net2272;
 wire net2273;
 wire net2274;
 wire net2275;
 wire net2276;
 wire net2277;
 wire net2278;
 wire net2279;
 wire net2280;
 wire net2281;
 wire net2282;
 wire net2283;
 wire net2284;
 wire net2285;
 wire net2286;
 wire net2287;
 wire net2288;
 wire net2289;
 wire net2290;
 wire net2291;
 wire net2292;
 wire net2293;
 wire net2294;
 wire net2295;
 wire net2296;
 wire net2297;
 wire net2298;
 wire net2299;
 wire net2300;
 wire net2301;
 wire net2302;
 wire net2303;
 wire net2304;
 wire net2305;
 wire net2306;
 wire net2307;
 wire net2308;
 wire net2309;
 wire net2310;
 wire net2311;
 wire net2312;
 wire net2313;
 wire net2314;
 wire net2315;
 wire net2316;
 wire net2317;
 wire net2318;
 wire net2319;
 wire net2320;
 wire net2321;
 wire net2322;
 wire net2323;
 wire net2324;
 wire net2325;
 wire net2326;
 wire net2327;
 wire net2328;
 wire net2329;
 wire net2330;
 wire net2331;
 wire net2332;
 wire net2333;
 wire net2334;
 wire net2335;
 wire net2336;
 wire net2337;
 wire net2338;
 wire net2339;
 wire net2340;
 wire net2341;
 wire net2342;
 wire net2343;
 wire net2344;
 wire net2345;
 wire net2346;
 wire net2347;
 wire net2348;
 wire net2349;
 wire net2350;
 wire net2351;
 wire net2352;
 wire net2353;
 wire net2354;
 wire net2355;
 wire net2356;
 wire net2357;
 wire net2358;
 wire net2359;
 wire net2360;
 wire net2361;
 wire net2362;
 wire net2363;
 wire net2364;
 wire net2365;
 wire net2366;
 wire net2367;
 wire net2368;
 wire net2369;
 wire net2370;
 wire net2371;
 wire net2372;
 wire net2373;
 wire net2374;
 wire net2375;
 wire net2376;
 wire net2377;
 wire net2378;
 wire net2379;
 wire net2380;
 wire net2381;
 wire net2382;
 wire net2383;
 wire net2384;
 wire net2385;
 wire net2386;
 wire net2387;
 wire net2388;
 wire net2389;
 wire net2390;
 wire net2391;
 wire net2392;
 wire net2393;
 wire net2394;
 wire net2395;
 wire net2396;
 wire net2397;
 wire net2398;
 wire net2399;
 wire net2400;
 wire net2401;
 wire net2402;
 wire net2403;
 wire net2404;
 wire net2405;
 wire net2406;
 wire net2407;
 wire net2408;
 wire net2409;
 wire net2410;
 wire net2411;
 wire net2412;
 wire net2413;
 wire net2414;
 wire net2415;
 wire net2416;
 wire net2417;
 wire net2418;
 wire net2419;
 wire net2420;
 wire net2421;
 wire net2422;
 wire net2423;
 wire net2424;
 wire net2425;
 wire net2426;
 wire net2427;
 wire net2428;
 wire net2429;
 wire net2430;
 wire net2431;
 wire net2432;
 wire net2433;
 wire net2434;
 wire net2435;
 wire net2436;
 wire net2437;
 wire net2438;
 wire net2439;
 wire net2440;
 wire net2441;
 wire net2442;
 wire net2443;
 wire net2444;
 wire net2445;
 wire net2446;
 wire net2447;
 wire net2448;
 wire net2449;
 wire net2450;
 wire net2451;
 wire net2452;
 wire net2453;
 wire net2454;
 wire net2455;
 wire net2456;
 wire net2457;
 wire net2458;
 wire net2459;
 wire net2460;
 wire net2461;
 wire net2462;
 wire net2463;
 wire net2464;
 wire net2465;
 wire net2466;
 wire net2467;
 wire net2468;
 wire net2469;
 wire net2470;
 wire net2471;
 wire net2472;
 wire net2473;
 wire net2474;
 wire net2475;
 wire net2476;
 wire net2477;
 wire net2478;
 wire net2479;
 wire net2480;
 wire net2481;
 wire net2482;
 wire net2483;
 wire net2484;
 wire net2485;
 wire net2486;
 wire net2487;
 wire net2488;
 wire net2489;
 wire net2490;
 wire net2491;
 wire net2492;
 wire net2493;
 wire net2494;
 wire net2495;
 wire net2496;
 wire net2497;
 wire net2498;
 wire net2499;
 wire net2500;
 wire net2501;
 wire net2502;
 wire net2503;
 wire net2504;
 wire net2505;
 wire net2506;
 wire net2507;
 wire net2508;
 wire net2509;
 wire net2510;
 wire net2511;
 wire net2512;
 wire net2513;
 wire net2514;
 wire net2515;
 wire net2516;
 wire net2517;
 wire net2518;
 wire net2519;
 wire net2520;
 wire net2521;
 wire net2522;
 wire net2523;
 wire net2524;
 wire net2525;
 wire net2526;
 wire net2527;
 wire net2528;
 wire net2529;
 wire net2530;
 wire net2531;
 wire net2532;
 wire net2533;
 wire net2534;
 wire net2535;
 wire net2536;
 wire net2537;
 wire net2538;
 wire net2539;
 wire net2540;
 wire net2541;
 wire net2542;
 wire net2543;
 wire net2544;
 wire net2545;
 wire net2546;
 wire net2547;
 wire net2548;
 wire net2549;
 wire net2550;
 wire net2551;
 wire net2552;
 wire net2553;
 wire net2554;
 wire net2555;
 wire net2556;
 wire net2557;
 wire net2558;
 wire net2559;
 wire net2560;
 wire net2561;
 wire net2562;
 wire net2563;
 wire net2564;
 wire net2565;
 wire net2566;
 wire net2567;
 wire net2568;
 wire net2569;
 wire net2570;
 wire net2571;
 wire net2572;
 wire net2573;
 wire net2574;
 wire net2575;
 wire net2576;
 wire net2577;
 wire net2578;
 wire net2579;
 wire net2580;
 wire net2581;
 wire net2582;
 wire net2583;
 wire net2584;
 wire net2585;
 wire net2586;
 wire net2587;
 wire net2588;
 wire net2589;
 wire net2590;
 wire net2591;
 wire net2592;
 wire net2593;
 wire net2594;
 wire net2595;
 wire net2596;
 wire net2597;
 wire net2598;
 wire net2599;
 wire net2600;
 wire net2601;
 wire net2602;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire clknet_0_clk;
 wire clknet_1_0__leaf_clk;
 wire clknet_1_1__leaf_clk;
 wire clknet_leaf_0_clk_regs;
 wire clknet_leaf_1_clk_regs;
 wire clknet_leaf_2_clk_regs;
 wire clknet_leaf_3_clk_regs;
 wire clknet_leaf_4_clk_regs;
 wire clknet_leaf_5_clk_regs;
 wire clknet_leaf_6_clk_regs;
 wire clknet_leaf_7_clk_regs;
 wire clknet_leaf_8_clk_regs;
 wire clknet_leaf_9_clk_regs;
 wire clknet_leaf_10_clk_regs;
 wire clknet_leaf_11_clk_regs;
 wire clknet_leaf_12_clk_regs;
 wire clknet_leaf_13_clk_regs;
 wire clknet_leaf_14_clk_regs;
 wire clknet_leaf_15_clk_regs;
 wire clknet_leaf_16_clk_regs;
 wire clknet_leaf_17_clk_regs;
 wire clknet_leaf_18_clk_regs;
 wire clknet_leaf_19_clk_regs;
 wire clknet_leaf_20_clk_regs;
 wire clknet_leaf_21_clk_regs;
 wire clknet_leaf_22_clk_regs;
 wire clknet_leaf_23_clk_regs;
 wire clknet_leaf_24_clk_regs;
 wire clknet_leaf_25_clk_regs;
 wire clknet_leaf_26_clk_regs;
 wire clknet_leaf_27_clk_regs;
 wire clknet_leaf_28_clk_regs;
 wire clknet_leaf_29_clk_regs;
 wire clknet_leaf_30_clk_regs;
 wire clknet_leaf_31_clk_regs;
 wire clknet_leaf_32_clk_regs;
 wire clknet_leaf_33_clk_regs;
 wire clknet_leaf_34_clk_regs;
 wire clknet_leaf_35_clk_regs;
 wire clknet_leaf_36_clk_regs;
 wire clknet_leaf_37_clk_regs;
 wire clknet_leaf_38_clk_regs;
 wire clknet_leaf_39_clk_regs;
 wire clknet_leaf_40_clk_regs;
 wire clknet_leaf_41_clk_regs;
 wire clknet_leaf_42_clk_regs;
 wire clknet_leaf_43_clk_regs;
 wire clknet_leaf_44_clk_regs;
 wire clknet_leaf_45_clk_regs;
 wire clknet_leaf_46_clk_regs;
 wire clknet_leaf_47_clk_regs;
 wire clknet_leaf_48_clk_regs;
 wire clknet_leaf_49_clk_regs;
 wire clknet_leaf_50_clk_regs;
 wire clknet_leaf_51_clk_regs;
 wire clknet_leaf_52_clk_regs;
 wire clknet_leaf_53_clk_regs;
 wire clknet_leaf_54_clk_regs;
 wire clknet_leaf_55_clk_regs;
 wire clknet_leaf_56_clk_regs;
 wire clknet_leaf_57_clk_regs;
 wire clknet_leaf_58_clk_regs;
 wire clknet_leaf_59_clk_regs;
 wire clknet_leaf_60_clk_regs;
 wire clknet_leaf_61_clk_regs;
 wire clknet_leaf_62_clk_regs;
 wire clknet_leaf_63_clk_regs;
 wire clknet_leaf_64_clk_regs;
 wire clknet_leaf_65_clk_regs;
 wire clknet_leaf_66_clk_regs;
 wire clknet_leaf_67_clk_regs;
 wire clknet_leaf_68_clk_regs;
 wire clknet_leaf_69_clk_regs;
 wire clknet_leaf_70_clk_regs;
 wire clknet_leaf_71_clk_regs;
 wire clknet_leaf_72_clk_regs;
 wire clknet_leaf_73_clk_regs;
 wire clknet_leaf_74_clk_regs;
 wire clknet_leaf_75_clk_regs;
 wire clknet_leaf_76_clk_regs;
 wire clknet_leaf_77_clk_regs;
 wire clknet_leaf_78_clk_regs;
 wire clknet_leaf_79_clk_regs;
 wire clknet_leaf_80_clk_regs;
 wire clknet_leaf_81_clk_regs;
 wire clknet_leaf_82_clk_regs;
 wire clknet_leaf_83_clk_regs;
 wire clknet_leaf_84_clk_regs;
 wire clknet_leaf_85_clk_regs;
 wire clknet_leaf_86_clk_regs;
 wire clknet_leaf_87_clk_regs;
 wire clknet_leaf_88_clk_regs;
 wire clknet_leaf_89_clk_regs;
 wire clknet_leaf_90_clk_regs;
 wire clknet_leaf_91_clk_regs;
 wire clknet_leaf_92_clk_regs;
 wire clknet_leaf_93_clk_regs;
 wire clknet_leaf_94_clk_regs;
 wire clknet_leaf_95_clk_regs;
 wire clknet_leaf_96_clk_regs;
 wire clknet_leaf_97_clk_regs;
 wire clknet_leaf_98_clk_regs;
 wire clknet_leaf_99_clk_regs;
 wire clknet_leaf_100_clk_regs;
 wire clknet_leaf_101_clk_regs;
 wire clknet_leaf_102_clk_regs;
 wire clknet_leaf_103_clk_regs;
 wire clknet_leaf_104_clk_regs;
 wire clknet_leaf_105_clk_regs;
 wire clknet_leaf_107_clk_regs;
 wire clknet_leaf_108_clk_regs;
 wire clknet_leaf_109_clk_regs;
 wire clknet_leaf_110_clk_regs;
 wire clknet_leaf_111_clk_regs;
 wire clknet_leaf_112_clk_regs;
 wire clknet_leaf_113_clk_regs;
 wire clknet_leaf_114_clk_regs;
 wire clknet_leaf_115_clk_regs;
 wire clknet_leaf_116_clk_regs;
 wire clknet_leaf_117_clk_regs;
 wire clknet_leaf_118_clk_regs;
 wire clknet_leaf_119_clk_regs;
 wire clknet_leaf_120_clk_regs;
 wire clknet_leaf_121_clk_regs;
 wire clknet_leaf_122_clk_regs;
 wire clknet_leaf_123_clk_regs;
 wire clknet_leaf_124_clk_regs;
 wire clknet_leaf_125_clk_regs;
 wire clknet_leaf_126_clk_regs;
 wire clknet_leaf_127_clk_regs;
 wire clknet_leaf_128_clk_regs;
 wire clknet_leaf_129_clk_regs;
 wire clknet_leaf_130_clk_regs;
 wire clknet_leaf_131_clk_regs;
 wire clknet_leaf_132_clk_regs;
 wire clknet_leaf_133_clk_regs;
 wire clknet_leaf_134_clk_regs;
 wire clknet_leaf_135_clk_regs;
 wire clknet_leaf_136_clk_regs;
 wire clknet_leaf_137_clk_regs;
 wire clknet_leaf_138_clk_regs;
 wire clknet_leaf_139_clk_regs;
 wire clknet_leaf_140_clk_regs;
 wire clknet_leaf_141_clk_regs;
 wire clknet_leaf_142_clk_regs;
 wire clknet_leaf_143_clk_regs;
 wire clknet_leaf_144_clk_regs;
 wire clknet_leaf_145_clk_regs;
 wire clknet_leaf_146_clk_regs;
 wire clknet_leaf_147_clk_regs;
 wire clknet_leaf_148_clk_regs;
 wire clknet_leaf_149_clk_regs;
 wire clknet_leaf_150_clk_regs;
 wire clknet_leaf_151_clk_regs;
 wire clknet_leaf_152_clk_regs;
 wire clknet_leaf_153_clk_regs;
 wire clknet_leaf_154_clk_regs;
 wire clknet_leaf_155_clk_regs;
 wire clknet_leaf_156_clk_regs;
 wire clknet_leaf_157_clk_regs;
 wire clknet_leaf_158_clk_regs;
 wire clknet_leaf_159_clk_regs;
 wire clknet_leaf_160_clk_regs;
 wire clknet_leaf_161_clk_regs;
 wire clknet_leaf_162_clk_regs;
 wire clknet_leaf_163_clk_regs;
 wire clknet_leaf_164_clk_regs;
 wire clknet_leaf_165_clk_regs;
 wire clknet_leaf_166_clk_regs;
 wire clknet_leaf_167_clk_regs;
 wire clknet_leaf_168_clk_regs;
 wire clknet_leaf_169_clk_regs;
 wire clknet_leaf_170_clk_regs;
 wire clknet_leaf_171_clk_regs;
 wire clknet_leaf_172_clk_regs;
 wire clknet_0_clk_regs;
 wire clknet_4_0_0_clk_regs;
 wire clknet_4_1_0_clk_regs;
 wire clknet_4_2_0_clk_regs;
 wire clknet_4_3_0_clk_regs;
 wire clknet_4_4_0_clk_regs;
 wire clknet_4_5_0_clk_regs;
 wire clknet_4_6_0_clk_regs;
 wire clknet_4_7_0_clk_regs;
 wire clknet_4_8_0_clk_regs;
 wire clknet_4_9_0_clk_regs;
 wire clknet_4_10_0_clk_regs;
 wire clknet_4_11_0_clk_regs;
 wire clknet_4_12_0_clk_regs;
 wire clknet_4_13_0_clk_regs;
 wire clknet_4_14_0_clk_regs;
 wire clknet_4_15_0_clk_regs;
 wire clknet_5_0__leaf_clk_regs;
 wire clknet_5_1__leaf_clk_regs;
 wire clknet_5_2__leaf_clk_regs;
 wire clknet_5_3__leaf_clk_regs;
 wire clknet_5_4__leaf_clk_regs;
 wire clknet_5_5__leaf_clk_regs;
 wire clknet_5_6__leaf_clk_regs;
 wire clknet_5_7__leaf_clk_regs;
 wire clknet_5_8__leaf_clk_regs;
 wire clknet_5_9__leaf_clk_regs;
 wire clknet_5_10__leaf_clk_regs;
 wire clknet_5_11__leaf_clk_regs;
 wire clknet_5_12__leaf_clk_regs;
 wire clknet_5_13__leaf_clk_regs;
 wire clknet_5_14__leaf_clk_regs;
 wire clknet_5_15__leaf_clk_regs;
 wire clknet_5_16__leaf_clk_regs;
 wire clknet_5_17__leaf_clk_regs;
 wire clknet_5_18__leaf_clk_regs;
 wire clknet_5_19__leaf_clk_regs;
 wire clknet_5_20__leaf_clk_regs;
 wire clknet_5_21__leaf_clk_regs;
 wire clknet_5_22__leaf_clk_regs;
 wire clknet_5_23__leaf_clk_regs;
 wire clknet_5_24__leaf_clk_regs;
 wire clknet_5_25__leaf_clk_regs;
 wire clknet_5_26__leaf_clk_regs;
 wire clknet_5_27__leaf_clk_regs;
 wire clknet_5_28__leaf_clk_regs;
 wire clknet_5_29__leaf_clk_regs;
 wire clknet_5_30__leaf_clk_regs;
 wire clknet_5_31__leaf_clk_regs;
 wire delaynet_0_clk;
 wire net1381;
 wire net1382;
 wire net1383;
 wire net1384;
 wire net1385;
 wire net1386;
 wire net1387;
 wire net1388;
 wire net1389;
 wire net1390;
 wire net1391;
 wire net1392;
 wire net1393;
 wire net1394;
 wire net1395;
 wire net1396;
 wire net1397;
 wire net1398;
 wire net1399;
 wire net1400;
 wire net1401;
 wire net1402;
 wire net1403;
 wire net1404;
 wire net1405;
 wire net1406;
 wire net1407;
 wire net1408;
 wire net1409;
 wire net1410;
 wire net1411;
 wire net1412;
 wire net1413;
 wire net1414;
 wire net1415;
 wire net1416;
 wire net1417;
 wire net1418;
 wire net1419;
 wire net1420;
 wire net1421;
 wire net1422;
 wire net1423;
 wire net1424;
 wire net1425;
 wire net1426;
 wire net1427;
 wire net1428;
 wire net1429;
 wire net1430;
 wire net1431;
 wire net1432;
 wire net1433;
 wire net1434;
 wire net1435;
 wire net1436;
 wire net1437;
 wire net1438;
 wire net1439;
 wire net1440;
 wire net1441;
 wire net1442;
 wire net1443;
 wire net1444;
 wire net1445;
 wire net1446;
 wire net1447;
 wire net1448;
 wire net1449;
 wire net1450;
 wire net1451;
 wire net1452;
 wire net1453;
 wire net1454;
 wire net1455;
 wire net1456;
 wire net1457;
 wire net1458;
 wire net1459;
 wire net1460;
 wire net1461;
 wire net1462;
 wire net1463;
 wire net1464;
 wire net1465;
 wire net1466;
 wire net1467;
 wire net1468;
 wire net1469;
 wire net1470;
 wire net1471;
 wire net1472;
 wire net1473;
 wire net1474;
 wire net1475;
 wire net1476;
 wire net1477;
 wire net1478;
 wire net1479;
 wire net1480;
 wire net1481;
 wire net1482;
 wire net1483;
 wire net1484;
 wire net1485;
 wire net1486;
 wire net1487;
 wire net1488;
 wire net1489;
 wire net1490;
 wire net1491;
 wire net1492;
 wire net1493;
 wire net1494;
 wire net1495;
 wire net1496;
 wire net1497;
 wire net1498;
 wire net1499;
 wire net1500;
 wire net1501;
 wire net1502;
 wire net1503;
 wire net1504;
 wire net1505;
 wire net1506;
 wire net1507;
 wire net1508;
 wire net1509;
 wire net1510;
 wire net1511;
 wire net1512;
 wire net1513;
 wire net1514;
 wire net1515;
 wire net1516;
 wire net1517;
 wire net1518;
 wire net1519;
 wire net1520;
 wire net1521;
 wire net1522;
 wire net1523;
 wire net1524;
 wire net1525;
 wire net1526;
 wire net1527;
 wire net1528;
 wire net1529;
 wire net1530;
 wire net1531;
 wire net1532;
 wire net1533;
 wire net1534;
 wire net1535;
 wire net1536;
 wire net1537;
 wire net1538;
 wire net1539;
 wire net1540;
 wire net1541;
 wire net1542;
 wire net1543;
 wire net1544;
 wire net1545;
 wire net1546;
 wire net1547;
 wire net1548;
 wire net1549;
 wire net1550;
 wire net1551;
 wire net1552;
 wire net1553;
 wire net1554;
 wire net1555;
 wire net1556;
 wire net1557;
 wire net1558;
 wire net1559;
 wire net1560;
 wire net1561;
 wire net1562;
 wire net1563;
 wire net1564;
 wire net1565;
 wire net1566;
 wire net1567;
 wire net1568;
 wire net1569;
 wire net1570;
 wire net1571;
 wire net1572;
 wire net1573;
 wire net1574;
 wire net1575;
 wire net1576;
 wire net1577;
 wire net1578;
 wire net1579;
 wire net1580;
 wire net1581;
 wire net1582;
 wire net1583;
 wire net1584;
 wire net1585;
 wire net1586;
 wire net1587;
 wire net1588;
 wire net1589;
 wire net1590;
 wire net1591;
 wire net1592;
 wire net1593;
 wire net1594;
 wire net1595;
 wire net1596;
 wire net1597;
 wire net1598;
 wire net1599;
 wire net1600;
 wire net1601;
 wire net1602;
 wire net1603;
 wire net1604;
 wire net1605;
 wire net1606;
 wire net1607;
 wire net1608;
 wire net1609;
 wire net1610;
 wire net1611;
 wire net1612;
 wire net1613;
 wire net1614;
 wire net1615;
 wire net1616;
 wire net1617;
 wire net1618;
 wire net1619;
 wire net1620;
 wire net1621;
 wire net1622;
 wire net1623;
 wire net1624;
 wire net1625;
 wire net1626;
 wire net1627;
 wire net1628;
 wire net1629;
 wire net1630;
 wire net1631;
 wire net1632;
 wire net1633;
 wire net1634;
 wire net1635;
 wire net1636;
 wire net1637;
 wire net1638;
 wire net1639;
 wire net1640;
 wire net1641;
 wire net1642;
 wire net1643;
 wire net1644;
 wire net1645;
 wire net1646;
 wire net1647;
 wire net1648;
 wire net1649;
 wire net1650;
 wire net1651;
 wire net1652;
 wire net1653;
 wire net1654;
 wire net1655;
 wire net1656;
 wire net1657;
 wire net1658;
 wire net1659;
 wire net1660;
 wire net1661;
 wire net1662;
 wire net1663;
 wire net1664;
 wire net1665;
 wire net1666;
 wire net1667;
 wire net1668;
 wire net1669;
 wire net1670;
 wire net1671;
 wire net1672;
 wire net1673;
 wire net1674;
 wire net1675;
 wire net1676;
 wire net1677;
 wire net1678;
 wire net1679;
 wire net1680;
 wire net1681;
 wire net1682;
 wire net1683;
 wire net1684;
 wire net1685;
 wire net1686;
 wire net1687;
 wire net1688;
 wire net1689;
 wire net1690;
 wire net1691;
 wire net1692;
 wire net1693;
 wire net1694;
 wire net1695;
 wire net1696;
 wire net1697;
 wire net1698;
 wire net1699;
 wire net1700;
 wire net1701;
 wire net1702;
 wire net1703;
 wire net1704;
 wire net1705;
 wire net1706;
 wire net1707;
 wire net1708;
 wire net1709;
 wire net1710;
 wire net1711;
 wire net1712;
 wire net1713;
 wire net1714;
 wire net1715;
 wire net1716;
 wire net1717;
 wire net1718;
 wire net1719;
 wire net1720;
 wire net1721;
 wire net1722;
 wire net1723;
 wire net1724;
 wire net1725;
 wire net1726;
 wire net1727;
 wire net1728;
 wire net1729;
 wire net1730;
 wire net1731;
 wire net1732;
 wire net1733;
 wire net1734;
 wire net1735;
 wire net1736;
 wire net1737;
 wire net1738;
 wire net1739;
 wire net1740;
 wire net1741;
 wire net1742;
 wire net1743;
 wire net1744;
 wire net1745;
 wire net1746;
 wire net1747;
 wire net1748;
 wire net2603;
 wire net2604;
 wire net2605;
 wire net2606;
 wire net2607;
 wire net2608;
 wire net2609;
 wire net2610;
 wire net2611;
 wire net2612;
 wire net2613;
 wire net2614;
 wire net2615;
 wire net2616;
 wire net2617;
 wire net2618;
 wire net2619;
 wire net2620;
 wire net2621;
 wire net2622;
 wire net2623;
 wire net2624;
 wire net2625;
 wire net2626;
 wire net2627;
 wire net2628;
 wire net2629;
 wire net2630;
 wire net2631;
 wire net2632;
 wire net2633;
 wire net2634;
 wire net2635;
 wire net2636;
 wire net2637;
 wire net2638;
 wire net2639;
 wire net2640;
 wire net2641;
 wire net2642;
 wire net2643;
 wire net2644;
 wire net2645;
 wire net2646;
 wire net2647;
 wire net2648;
 wire net2649;
 wire net2650;
 wire net2651;
 wire net2652;
 wire net2653;
 wire net2654;
 wire net2655;
 wire net2656;
 wire net2657;
 wire net2658;
 wire net2659;
 wire net2660;
 wire net2661;
 wire net2662;
 wire net2663;
 wire net2664;
 wire net2665;
 wire net2666;
 wire net2667;
 wire net2668;
 wire net2669;
 wire net2670;
 wire net2671;
 wire net2672;
 wire net2673;
 wire net2674;
 wire net2675;
 wire net2676;
 wire net2677;
 wire net2678;
 wire net2679;
 wire net2680;
 wire net2681;
 wire net2682;
 wire net2683;
 wire net2684;
 wire net2685;
 wire net2686;
 wire net2687;
 wire net2688;
 wire net2689;
 wire net2690;
 wire net2691;
 wire net2692;
 wire net2693;
 wire net2694;
 wire net2695;
 wire net2696;
 wire net2697;
 wire net2698;
 wire net2699;
 wire net2700;
 wire net2701;
 wire net2702;
 wire net2703;
 wire net2704;
 wire net2705;
 wire net2706;
 wire net2707;
 wire net2708;
 wire net2709;
 wire net2710;
 wire net2711;
 wire net2712;
 wire net2713;
 wire net2714;
 wire net2715;
 wire net2716;
 wire net2717;
 wire net2718;
 wire net2719;
 wire net2720;
 wire net2721;
 wire net2722;
 wire net2723;
 wire net2724;
 wire net2725;
 wire net2726;
 wire net2727;
 wire net2728;
 wire net2729;
 wire net2730;
 wire net2731;
 wire net2732;
 wire net2733;
 wire net2734;
 wire net2735;
 wire net2736;
 wire net2737;
 wire net2738;
 wire net2739;
 wire net2740;
 wire net2741;
 wire net2742;
 wire net2743;
 wire net2744;
 wire net2745;
 wire net2746;
 wire net2747;
 wire net2748;
 wire net2749;
 wire net2750;
 wire net2751;
 wire net2752;
 wire net2753;
 wire net2754;
 wire net2755;
 wire net2756;
 wire net2757;
 wire net2758;
 wire net2759;
 wire net2760;
 wire net2761;
 wire net2762;
 wire net2763;
 wire net2764;
 wire net2765;
 wire net2766;
 wire net2767;
 wire net2768;
 wire net2769;
 wire net2770;
 wire net2771;
 wire net2772;
 wire net2773;
 wire net2774;
 wire net2775;
 wire net2776;
 wire net2777;
 wire net2778;
 wire net2779;
 wire net2780;
 wire net2781;
 wire net2782;
 wire net2783;
 wire net2784;
 wire net2785;
 wire net2786;
 wire net2787;
 wire net2788;
 wire net2789;
 wire net2790;
 wire net2791;
 wire net2792;
 wire net2793;
 wire net2794;
 wire net2795;
 wire net2796;
 wire net2797;
 wire net2798;
 wire net2799;
 wire net2800;
 wire net2801;
 wire net2802;
 wire net2803;
 wire net2804;
 wire net2805;
 wire net2806;
 wire net2807;
 wire net2808;
 wire net2809;
 wire net2810;
 wire net2811;
 wire net2812;
 wire net2813;
 wire net2814;
 wire net2815;
 wire net2816;
 wire net2817;
 wire net2818;
 wire net2819;
 wire net2820;
 wire net2821;
 wire net2822;
 wire net2823;
 wire net2824;
 wire net2825;
 wire net2826;
 wire net2827;
 wire net2828;
 wire net2829;
 wire net2830;
 wire net2831;
 wire net2832;
 wire net2833;
 wire net2834;
 wire net2835;
 wire net2836;
 wire net2837;
 wire net2838;
 wire net2839;
 wire net2840;
 wire net2841;
 wire net2842;
 wire net2843;
 wire net2844;
 wire net2845;
 wire net2846;
 wire net2847;
 wire net2848;
 wire net2849;
 wire net2850;
 wire net2851;
 wire net2852;
 wire net2853;
 wire net2854;
 wire net2855;
 wire net2856;
 wire net2857;
 wire net2858;
 wire net2859;
 wire net2860;
 wire net2861;
 wire net2862;
 wire net2863;
 wire net2864;
 wire net2865;
 wire net2866;
 wire net2867;
 wire net2868;
 wire net2869;
 wire net2870;
 wire net2871;
 wire net2872;
 wire net2873;
 wire net2874;
 wire net2875;
 wire net2876;
 wire net2877;
 wire net2878;
 wire net2879;
 wire net2880;
 wire net2881;
 wire net2882;
 wire net2883;
 wire net2884;
 wire net2885;
 wire net2886;
 wire net2887;
 wire net2888;
 wire net2889;
 wire net2890;
 wire net2891;
 wire net2892;
 wire net2893;
 wire net2894;
 wire net2895;
 wire net2896;
 wire net2897;
 wire net2898;
 wire net2899;
 wire net2900;
 wire net2901;
 wire net2902;
 wire net2903;
 wire net2904;
 wire net2905;
 wire net2906;
 wire net2907;
 wire net2908;
 wire net2909;
 wire net2910;
 wire net2911;
 wire net2912;
 wire net2913;
 wire net2914;
 wire net2915;
 wire net2916;
 wire net2917;
 wire net2918;
 wire net2919;
 wire net2920;
 wire net2921;
 wire net2922;
 wire net2923;
 wire net2924;
 wire net2925;
 wire net2926;
 wire net2927;
 wire net2928;
 wire net2929;
 wire net2930;
 wire net2931;
 wire net2932;
 wire net2933;
 wire net2934;
 wire net2935;
 wire net2936;
 wire net2937;
 wire net2938;
 wire net2939;
 wire net2940;
 wire net2941;
 wire net2942;
 wire net2943;
 wire net2944;
 wire net2945;
 wire net2946;
 wire net2947;
 wire net2948;
 wire net2949;
 wire net2950;
 wire net2951;
 wire net2952;
 wire net2953;
 wire net2954;
 wire net2955;
 wire net2956;
 wire net2957;
 wire net2958;
 wire net2959;
 wire net2960;
 wire net2961;
 wire net2962;
 wire net2963;
 wire net2964;
 wire net2965;
 wire net2966;
 wire net2967;
 wire net2968;
 wire net2969;
 wire net2970;
 wire net2971;
 wire net2972;
 wire net2973;
 wire net2974;
 wire net2975;
 wire net2976;
 wire net2977;
 wire net2978;
 wire net2979;
 wire net2980;
 wire net2981;
 wire net2982;
 wire net2983;
 wire net2984;
 wire net2985;
 wire net2986;
 wire net2987;
 wire net2988;
 wire net2989;
 wire net2990;
 wire net2991;
 wire net2992;
 wire net2993;
 wire net2994;
 wire net2995;
 wire net2996;
 wire net2997;
 wire net2998;
 wire net2999;
 wire net3000;
 wire net3001;
 wire net3002;
 wire net3003;
 wire net3004;
 wire net3005;
 wire net3006;
 wire net3007;
 wire net3008;
 wire net3009;
 wire net3010;
 wire net3011;
 wire net3012;
 wire net3013;
 wire net3014;
 wire net3015;
 wire net3016;
 wire net3017;
 wire net3018;
 wire net3019;
 wire net3020;
 wire net3021;
 wire net3022;
 wire net3023;
 wire net3024;
 wire net3025;
 wire net3026;
 wire net3027;
 wire net3028;
 wire net3029;
 wire net3030;
 wire net3031;
 wire net3032;
 wire net3033;
 wire net3034;
 wire net3035;
 wire net3036;
 wire net3037;
 wire net3038;
 wire net3039;
 wire net3040;
 wire net3041;
 wire net3042;
 wire net3043;
 wire net3044;
 wire net3045;
 wire net3046;
 wire net3047;
 wire net3048;
 wire net3049;
 wire net3050;
 wire net3051;
 wire net3052;
 wire net3053;
 wire net3054;
 wire net3055;
 wire net3056;
 wire net3057;
 wire net3058;
 wire net3059;
 wire net3060;
 wire net3061;
 wire net3062;
 wire net3063;
 wire net3064;
 wire net3065;
 wire net3066;
 wire net3067;
 wire net3068;
 wire net3069;
 wire net3070;
 wire net3071;
 wire net3072;
 wire net3073;
 wire net3074;
 wire net3075;
 wire net3076;
 wire net3077;
 wire net3078;
 wire net3079;
 wire net3080;
 wire net3081;
 wire net3082;
 wire net3083;
 wire net3084;
 wire net3085;
 wire net3086;
 wire net3087;
 wire net3088;
 wire net3089;
 wire net3090;
 wire net3091;
 wire net3092;
 wire net3093;
 wire net3094;
 wire net3095;
 wire net3096;
 wire net3097;
 wire net3098;
 wire net3099;
 wire net3100;
 wire net3101;
 wire net3102;
 wire net3103;
 wire net3104;
 wire net3105;
 wire net3106;
 wire net3107;
 wire net3108;
 wire net3109;
 wire net3110;
 wire net3111;
 wire net3112;
 wire net3113;
 wire net3114;
 wire net3115;
 wire net3116;
 wire net3117;
 wire net3118;
 wire net3119;
 wire net3120;
 wire net3121;
 wire net3122;
 wire net3123;
 wire net3124;
 wire net3125;
 wire net3126;
 wire net3127;
 wire net3128;
 wire net3129;
 wire net3130;
 wire net3131;
 wire net3132;
 wire net3133;
 wire net3134;
 wire net3135;
 wire net3136;
 wire net3137;
 wire net3138;
 wire net3139;
 wire net3140;
 wire net3141;
 wire net3142;
 wire net3143;
 wire net3144;
 wire net3145;
 wire net3146;
 wire net3147;
 wire net3148;
 wire net3149;
 wire net3150;
 wire net3151;
 wire net3152;
 wire net3153;
 wire net3154;
 wire net3155;
 wire net3156;
 wire net3157;
 wire net3158;
 wire net3159;
 wire net3160;
 wire net3161;
 wire net3162;
 wire net3163;
 wire net3164;
 wire net3165;
 wire net3166;
 wire net3167;
 wire net3168;
 wire net3169;
 wire net3170;
 wire net3171;
 wire net3172;
 wire net3173;
 wire net3174;
 wire net3175;
 wire net3176;
 wire net3177;
 wire net3178;
 wire net3179;
 wire net3180;
 wire net3181;
 wire net3182;
 wire net3183;
 wire net3184;
 wire net3185;
 wire net3186;
 wire net3187;
 wire net3188;
 wire net3189;
 wire net3190;
 wire net3191;
 wire net3192;
 wire net3193;
 wire net3194;
 wire net3195;
 wire net3196;
 wire net3197;
 wire net3198;
 wire net3199;
 wire net3200;
 wire net3201;
 wire net3202;
 wire net3203;
 wire net3204;
 wire net3205;
 wire net3206;
 wire net3207;
 wire net3208;
 wire net3209;
 wire net3210;
 wire net3211;
 wire net3212;
 wire net3213;
 wire net3214;
 wire net3215;
 wire net3216;
 wire net3217;
 wire net3218;
 wire net3219;
 wire net3220;
 wire net3221;
 wire net3222;
 wire net3223;
 wire net3224;
 wire net3225;
 wire net3226;
 wire net3227;
 wire net3228;
 wire net3229;
 wire net3230;
 wire net3231;
 wire net3232;
 wire net3233;
 wire net3234;
 wire net3235;
 wire net3236;
 wire net3237;
 wire net3238;
 wire net3239;
 wire net3240;
 wire net3241;
 wire net3242;
 wire net3243;
 wire net3244;
 wire net3245;
 wire net3246;
 wire net3247;
 wire net3248;
 wire net3249;
 wire net3250;
 wire net3251;
 wire net3252;
 wire net3253;
 wire net3254;
 wire net3255;
 wire net3256;
 wire net3257;
 wire net3258;
 wire net3259;
 wire net3260;
 wire net3261;
 wire net3262;
 wire net3263;
 wire net3264;
 wire net3265;
 wire net3266;
 wire net3267;
 wire net3268;
 wire net3269;
 wire net3270;
 wire net3271;
 wire net3272;
 wire net3273;
 wire net3274;
 wire net3275;
 wire net3276;
 wire net3277;
 wire net3278;
 wire net3279;
 wire net3280;
 wire net3281;
 wire net3282;
 wire net3283;
 wire net3284;
 wire net3285;
 wire net3286;
 wire net3287;
 wire net3288;
 wire net3289;
 wire net3290;
 wire net3291;
 wire net3292;
 wire net3293;
 wire net3294;
 wire net3295;
 wire net3296;
 wire net3297;
 wire net3298;
 wire net3299;
 wire net3300;
 wire net3301;
 wire net3302;
 wire net3303;
 wire net3304;
 wire net3305;
 wire net3306;
 wire net3307;
 wire net3308;
 wire net3309;
 wire net3310;
 wire net3311;
 wire net3312;
 wire net3313;
 wire net3314;
 wire net3315;
 wire net3316;
 wire net3317;
 wire net3318;
 wire net3319;
 wire net3320;
 wire net3321;
 wire net3322;
 wire net3323;
 wire net3324;
 wire net3325;
 wire net3326;
 wire net3327;
 wire net3328;
 wire net3329;
 wire net3330;
 wire net3331;
 wire net3332;
 wire net3333;
 wire net3334;
 wire net3335;
 wire net3336;
 wire net3337;
 wire net3338;
 wire net3339;
 wire net3340;
 wire net3341;
 wire net3342;
 wire net3343;
 wire net3344;
 wire net3345;
 wire net3346;
 wire net3347;
 wire net3348;
 wire net3349;
 wire net3350;
 wire net3351;
 wire net3352;
 wire net3353;
 wire net3354;
 wire net3355;
 wire net3356;
 wire net3357;
 wire net3358;
 wire net3359;
 wire net3360;
 wire net3361;
 wire net3362;
 wire net3363;
 wire net3364;
 wire net3365;
 wire net3366;
 wire net3367;
 wire net3368;
 wire net3369;
 wire net3370;
 wire net3371;
 wire net3372;
 wire net3373;
 wire net3374;
 wire net3375;
 wire net3376;
 wire net3377;
 wire net3378;
 wire net3379;
 wire net3380;
 wire net3381;
 wire net3382;
 wire net3383;
 wire net3384;
 wire net3385;
 wire net3386;
 wire net3387;
 wire net3388;
 wire net3389;
 wire net3390;
 wire net3391;
 wire net3392;
 wire net3393;
 wire net3394;
 wire net3395;
 wire net3396;
 wire net3397;
 wire net3398;
 wire net3399;
 wire net3400;
 wire net3401;
 wire net3402;
 wire net3403;
 wire net3404;
 wire net3405;
 wire net3406;
 wire net3407;
 wire net3408;
 wire net3409;
 wire net3410;
 wire net3411;
 wire net3412;
 wire net3413;
 wire net3414;
 wire net3415;
 wire net3416;
 wire net3417;
 wire net3418;
 wire net3419;
 wire net3420;
 wire net3421;
 wire net3422;
 wire net3423;
 wire net3424;
 wire net3425;
 wire net3426;
 wire net3427;
 wire net3428;
 wire net3429;
 wire net3430;
 wire net3431;
 wire net3432;
 wire net3433;
 wire net3434;
 wire net3435;
 wire net3436;
 wire net3437;
 wire net3438;
 wire net3439;
 wire net3440;
 wire net3441;
 wire net3442;
 wire net3443;
 wire net3444;
 wire net3445;
 wire net3446;
 wire net3447;
 wire net3448;
 wire net3449;
 wire net3450;
 wire net3451;
 wire net3452;
 wire net3453;
 wire net3454;
 wire net3455;
 wire net3456;
 wire net3457;
 wire net3458;
 wire net3459;
 wire net3460;
 wire net3461;
 wire net3462;
 wire net3463;
 wire net3464;
 wire net3465;
 wire net3466;
 wire net3467;
 wire net3468;
 wire net3469;
 wire net3470;
 wire net3471;
 wire net3472;
 wire net3473;
 wire net3474;
 wire net3475;
 wire net3476;
 wire net3477;
 wire net3478;
 wire net3479;
 wire net3480;
 wire net3481;
 wire net3482;
 wire net3483;
 wire net3484;
 wire net3485;
 wire net3486;
 wire net3487;
 wire net3488;
 wire net3489;
 wire net3490;
 wire net3491;
 wire net3492;
 wire net3493;
 wire net3494;
 wire net3495;
 wire net3496;
 wire net3497;
 wire net3498;
 wire net3499;
 wire net3500;
 wire net3501;
 wire net3502;
 wire net3503;
 wire net3504;
 wire net3505;
 wire net3506;
 wire net3507;
 wire net3508;
 wire net3509;
 wire net3510;
 wire net3511;
 wire net3512;
 wire net3513;
 wire net3514;
 wire net3515;
 wire net3516;
 wire net3517;
 wire net3518;
 wire net3519;
 wire net3520;
 wire net3521;
 wire net3522;
 wire net3523;
 wire net3524;
 wire net3525;
 wire net3526;
 wire net3527;
 wire net3528;
 wire net3529;
 wire net3530;
 wire net3531;
 wire net3532;
 wire net3533;
 wire net3534;
 wire net3535;
 wire net3536;
 wire net3537;
 wire net3538;
 wire net3539;
 wire net3540;
 wire net3541;
 wire net3542;
 wire net3543;
 wire net3544;
 wire net3545;
 wire net3546;
 wire net3547;
 wire net3548;
 wire net3549;
 wire net3550;
 wire net3551;
 wire net3552;
 wire net3553;
 wire net3554;
 wire net3555;
 wire net3556;
 wire net3557;
 wire net3558;
 wire net3559;
 wire net3560;
 wire net3561;
 wire net3562;
 wire net3563;
 wire net3564;
 wire net3565;
 wire net3566;
 wire net3567;
 wire net3568;
 wire net3569;
 wire net3570;
 wire net3571;
 wire net3572;
 wire net3573;
 wire net3574;
 wire net3575;
 wire net3576;
 wire net3577;
 wire net3578;
 wire net3579;
 wire net3580;
 wire net3581;
 wire net3582;
 wire net3583;
 wire net3584;
 wire net3585;
 wire net3586;
 wire net3587;
 wire net3588;
 wire net3589;
 wire net3590;
 wire net3591;
 wire net3592;
 wire net3593;
 wire net3594;
 wire net3595;
 wire net3596;
 wire net3597;
 wire net3598;
 wire net3599;
 wire net3600;
 wire net3601;
 wire net3602;
 wire net3603;
 wire net3604;
 wire net3605;
 wire net3606;
 wire net3607;
 wire net3608;
 wire net3609;
 wire net3610;
 wire net3611;
 wire net3612;
 wire net3613;
 wire net3614;
 wire net3615;
 wire net3616;
 wire net3617;
 wire net3618;
 wire net3619;
 wire net3620;
 wire net3621;
 wire net3622;
 wire net3623;
 wire net3624;
 wire net3625;
 wire net3626;
 wire net3627;
 wire net3628;
 wire net3629;
 wire net3630;
 wire net3631;
 wire net3632;
 wire net3633;
 wire net3634;
 wire net3635;
 wire net3636;
 wire net3637;
 wire net3638;
 wire net3639;
 wire net3640;
 wire net3641;
 wire net3642;
 wire net3643;
 wire net3644;
 wire net3645;
 wire net3646;
 wire net3647;
 wire net3648;
 wire net3649;
 wire net3650;
 wire net3651;
 wire net3652;
 wire net3653;
 wire net3654;
 wire net3655;
 wire net3656;
 wire net3657;
 wire net3658;
 wire net3659;
 wire net3660;
 wire net3661;
 wire net3662;
 wire net3663;
 wire net3664;
 wire net3665;
 wire net3666;
 wire net3667;
 wire net3668;
 wire net3669;
 wire net3670;
 wire net3671;
 wire net3672;
 wire net3673;
 wire net3674;
 wire net3675;
 wire net3676;
 wire net3677;
 wire net3678;
 wire net3679;
 wire net3680;
 wire net3681;
 wire net3682;
 wire net3683;
 wire net3684;
 wire net3685;
 wire net3686;
 wire net3687;
 wire net3688;
 wire net3689;
 wire net3690;
 wire net3691;
 wire net3692;
 wire net3693;
 wire net3694;
 wire net3695;
 wire net3696;
 wire net3697;
 wire net3698;
 wire net3699;
 wire net3700;
 wire net3701;
 wire net3702;
 wire net3703;
 wire net3704;
 wire net3705;
 wire net3706;
 wire net3707;
 wire net3708;
 wire net3709;
 wire net3710;
 wire net3711;
 wire net3712;
 wire net3713;
 wire net3714;
 wire net3715;
 wire net3716;
 wire net3717;
 wire net3718;
 wire net3719;
 wire net3720;
 wire net3721;
 wire net3722;
 wire net3723;
 wire net3724;
 wire net3725;
 wire net3726;
 wire net3727;
 wire net3728;
 wire net3729;
 wire net3730;
 wire net3731;
 wire net3732;
 wire net3733;
 wire net3734;
 wire net3735;
 wire net3736;
 wire net3737;
 wire net3738;
 wire net3739;
 wire net3740;
 wire net3741;
 wire net3742;
 wire net3743;
 wire net3744;
 wire net3745;
 wire net3746;
 wire net3747;
 wire net3748;
 wire net3749;
 wire net3750;
 wire net3751;
 wire net3752;
 wire net3753;
 wire net3754;
 wire net3755;
 wire net3756;
 wire net3757;
 wire net3758;
 wire net3759;
 wire net3760;
 wire net3761;
 wire net3762;
 wire net3763;
 wire net3764;
 wire net3765;
 wire net3766;
 wire net3767;
 wire net3768;
 wire net3769;
 wire net3770;
 wire net3771;
 wire net3772;
 wire net3773;
 wire net3774;
 wire net3775;
 wire net3776;
 wire net3777;
 wire net3778;
 wire net3779;
 wire net3780;
 wire net3781;
 wire net3782;
 wire net3783;
 wire net3784;
 wire net3785;
 wire net3786;
 wire net3787;
 wire net3788;
 wire net3789;
 wire net3790;
 wire net3791;
 wire net3792;
 wire net3793;
 wire net3794;
 wire net3795;
 wire net3796;
 wire net3797;
 wire net3798;
 wire net3799;
 wire net3800;
 wire net3801;
 wire net3802;
 wire net3803;
 wire net3804;
 wire net3805;
 wire net3806;
 wire net3807;
 wire net3808;
 wire net3809;
 wire net3810;
 wire net3811;
 wire net3812;
 wire net3813;
 wire net3814;
 wire net3815;
 wire net3816;
 wire net3817;
 wire net3818;
 wire [0:0] \cpu.cpu.alu.add_cy_r ;
 wire [0:0] \cpu.cpu.alu.i_rs1 ;
 wire [0:0] \cpu.cpu.bufreg.c_r ;
 wire [0:0] \cpu.cpu.csr_imm ;
 wire [0:0] \cpu.cpu.ctrl.pc ;
 wire [0:0] \cpu.cpu.ctrl.pc_plus_4_cy_r_w ;
 wire [0:0] \cpu.cpu.ctrl.pc_plus_offset_cy_r_w ;
 wire [0:0] \cpu.cpu.o_wdata0 ;

 sg13g2_inv_1 _05283_ (.Y(_01333_),
    .A(net3476));
 sg13g2_inv_4 _05284_ (.A(net2599),
    .Y(_01334_));
 sg13g2_inv_1 _05285_ (.Y(_01335_),
    .A(net3720));
 sg13g2_inv_1 _05286_ (.Y(_01336_),
    .A(net3284));
 sg13g2_inv_1 _05287_ (.Y(_01337_),
    .A(net3273));
 sg13g2_inv_1 _05288_ (.Y(_01338_),
    .A(net3391));
 sg13g2_inv_1 _05289_ (.Y(_01339_),
    .A(net3361));
 sg13g2_inv_1 _05290_ (.Y(_01340_),
    .A(net3717));
 sg13g2_inv_1 _05291_ (.Y(_01341_),
    .A(\cpu.cpu.bufreg.data[0] ));
 sg13g2_inv_2 _05292_ (.Y(_01342_),
    .A(net3660));
 sg13g2_inv_1 _05293_ (.Y(_01343_),
    .A(net3725));
 sg13g2_inv_2 _05294_ (.Y(_01344_),
    .A(net3704));
 sg13g2_inv_2 _05295_ (.Y(_01345_),
    .A(net2577));
 sg13g2_inv_2 _05296_ (.Y(_01346_),
    .A(\cpu.cpu.bufreg.i_right_shift_op ));
 sg13g2_inv_1 _05297_ (.Y(_01347_),
    .A(net3757));
 sg13g2_inv_1 _05298_ (.Y(_01348_),
    .A(net3752));
 sg13g2_inv_1 _05299_ (.Y(_01349_),
    .A(net3674));
 sg13g2_inv_1 _05300_ (.Y(_01350_),
    .A(net3734));
 sg13g2_inv_1 _05301_ (.Y(_01351_),
    .A(net3739));
 sg13g2_inv_1 _05302_ (.Y(_01352_),
    .A(net3742));
 sg13g2_inv_2 _05303_ (.Y(_01353_),
    .A(net3728));
 sg13g2_inv_1 _05304_ (.Y(_01354_),
    .A(net3594));
 sg13g2_inv_2 _05305_ (.Y(_01355_),
    .A(net3392));
 sg13g2_inv_2 _05306_ (.Y(_01356_),
    .A(net3724));
 sg13g2_inv_1 _05307_ (.Y(_01357_),
    .A(net3626));
 sg13g2_inv_2 _05308_ (.Y(_01358_),
    .A(net3713));
 sg13g2_inv_1 _05309_ (.Y(_01359_),
    .A(net3707));
 sg13g2_inv_1 _05310_ (.Y(_01360_),
    .A(net3680));
 sg13g2_inv_1 _05311_ (.Y(_01361_),
    .A(net3584));
 sg13g2_inv_1 _05312_ (.Y(_01362_),
    .A(\cpu.cpu.immdec.gen_immdec_w_eq_1.imm24_20[0] ));
 sg13g2_inv_1 _05313_ (.Y(_01363_),
    .A(net3606));
 sg13g2_inv_1 _05314_ (.Y(_01364_),
    .A(net3616));
 sg13g2_inv_1 _05315_ (.Y(_01365_),
    .A(net3582));
 sg13g2_inv_1 _05316_ (.Y(_01366_),
    .A(net3615));
 sg13g2_inv_1 _05317_ (.Y(_01367_),
    .A(\cpu.cpu.immdec.gen_immdec_w_eq_1.imm11_7[3] ));
 sg13g2_inv_1 _05318_ (.Y(_01368_),
    .A(\cpu.cpu.immdec.gen_immdec_w_eq_1.imm19_12_20[8] ));
 sg13g2_inv_1 _05319_ (.Y(_01369_),
    .A(net3440));
 sg13g2_inv_1 _05320_ (.Y(_01370_),
    .A(net3762));
 sg13g2_buf_8 clkbuf_regs_0_clk (.A(clk),
    .X(clk_regs));
 sg13g2_nor2_1 _05322_ (.A(\ram_spi_if.state_reg[1] ),
    .B(\ram_spi_if.state_reg[2] ),
    .Y(_01371_));
 sg13g2_nand2_1 _05323_ (.Y(_01372_),
    .A(_01343_),
    .B(_01344_));
 sg13g2_nor2_2 _05324_ (.A(net2594),
    .B(_01372_),
    .Y(_01373_));
 sg13g2_inv_1 _05325_ (.Y(_01374_),
    .A(_01373_));
 sg13g2_a21o_1 _05326_ (.A2(_01372_),
    .A1(net2594),
    .B1(net2595),
    .X(_01375_));
 sg13g2_nor2_2 _05327_ (.A(_01373_),
    .B(_01375_),
    .Y(_01376_));
 sg13g2_or2_1 _05328_ (.X(_01377_),
    .B(_01375_),
    .A(_01373_));
 sg13g2_nor2_2 _05329_ (.A(\cpu.cpu.bufreg.data[0] ),
    .B(\cpu.cpu.bufreg.data[1] ),
    .Y(_01378_));
 sg13g2_nand3b_1 _05330_ (.B(net3704),
    .C(net3725),
    .Y(_01379_),
    .A_N(net2594));
 sg13g2_nor2_1 _05331_ (.A(net2595),
    .B(_01379_),
    .Y(_01380_));
 sg13g2_nand2_1 _05332_ (.Y(_01381_),
    .A(net2571),
    .B(_01380_));
 sg13g2_o21ai_1 _05333_ (.B1(_01376_),
    .Y(_01382_),
    .A1(_01378_),
    .A2(_01381_));
 sg13g2_nor2_1 _05334_ (.A(net2570),
    .B(\cpu.cpu.bne_or_bge ),
    .Y(_01383_));
 sg13g2_nor2b_1 _05335_ (.A(\cpu.cpu.bufreg.data[0] ),
    .B_N(\cpu.cpu.bufreg.data[1] ),
    .Y(_01384_));
 sg13g2_and2_1 _05336_ (.A(_01383_),
    .B(_01384_),
    .X(_01385_));
 sg13g2_nor3_1 _05337_ (.A(_01341_),
    .B(\cpu.cpu.bufreg.data[1] ),
    .C(net2571),
    .Y(_01386_));
 sg13g2_nor2b_2 _05338_ (.A(net2570),
    .B_N(\cpu.cpu.bne_or_bge ),
    .Y(_01387_));
 sg13g2_a21oi_1 _05339_ (.A1(_01378_),
    .A2(_01387_),
    .Y(_01388_),
    .B1(_01386_));
 sg13g2_o21ai_1 _05340_ (.B1(_01388_),
    .Y(_01389_),
    .A1(\cpu.arbiter.i_wb_mem_rdt[31] ),
    .A2(_01385_));
 sg13g2_a21oi_1 _05341_ (.A1(_01353_),
    .A2(_01385_),
    .Y(_01390_),
    .B1(_01389_));
 sg13g2_nor2b_1 _05342_ (.A(_01388_),
    .B_N(\cpu.arbiter.i_wb_mem_rdt[15] ),
    .Y(_01391_));
 sg13g2_a21oi_1 _05343_ (.A1(_01378_),
    .A2(_01383_),
    .Y(_01392_),
    .B1(_01391_));
 sg13g2_nand2b_1 _05344_ (.Y(_01393_),
    .B(_01392_),
    .A_N(_01390_));
 sg13g2_nand3b_1 _05345_ (.B(_01378_),
    .C(_01383_),
    .Y(_01394_),
    .A_N(\cpu.arbiter.i_wb_mem_rdt[7] ));
 sg13g2_nand3_1 _05346_ (.B(_01393_),
    .C(_01394_),
    .A(_01380_),
    .Y(_01395_));
 sg13g2_nor3_2 _05347_ (.A(net3756),
    .B(net2594),
    .C(_01344_),
    .Y(_01396_));
 sg13g2_nor2b_1 _05348_ (.A(net2596),
    .B_N(_01396_),
    .Y(_01397_));
 sg13g2_nor3_1 _05349_ (.A(_01343_),
    .B(net2594),
    .C(net3704),
    .Y(_01398_));
 sg13g2_nand2b_1 _05350_ (.Y(_01399_),
    .B(_01398_),
    .A_N(net2596));
 sg13g2_inv_1 _05351_ (.Y(_01400_),
    .A(_01399_));
 sg13g2_a221oi_1 _05352_ (.B2(\cpu.arbiter.i_wb_mem_rdt[7] ),
    .C1(_01382_),
    .B1(_01400_),
    .A1(\cpu.arbiter.i_wb_mem_rdt[15] ),
    .Y(_01401_),
    .A2(_01397_));
 sg13g2_a22oi_1 _05353_ (.Y(_00619_),
    .B1(_01395_),
    .B2(_01401_),
    .A2(_01382_),
    .A1(_01333_));
 sg13g2_nor3_1 _05354_ (.A(\cpu.rf_ram_if.rcnt[3] ),
    .B(\cpu.rf_ram_if.rcnt[2] ),
    .C(net3767),
    .Y(_01402_));
 sg13g2_nand2_1 _05355_ (.Y(_01403_),
    .A(\cpu.rf_ram_if.rcnt[0] ),
    .B(_01402_));
 sg13g2_or2_1 _05356_ (.X(_01404_),
    .B(_01403_),
    .A(\cpu.rf_ram_if.rcnt[1] ));
 sg13g2_inv_2 _05357_ (.Y(\cpu.rf_ram_if.rtrig0 ),
    .A(net2377));
 sg13g2_nand3_1 _05358_ (.B(net2594),
    .C(_01371_),
    .A(net2595),
    .Y(_01405_));
 sg13g2_inv_1 _05359_ (.Y(_01406_),
    .A(_01405_));
 sg13g2_nor2_1 _05360_ (.A(net2596),
    .B(_01374_),
    .Y(_01407_));
 sg13g2_o21ai_1 _05361_ (.B1(_01405_),
    .Y(\ram_spi_if.spi_cs_n ),
    .A1(net2595),
    .A2(_01374_));
 sg13g2_nor2_1 _05362_ (.A(net1417),
    .B(_01377_),
    .Y(_00065_));
 sg13g2_xnor2_1 _05363_ (.Y(_01408_),
    .A(net3691),
    .B(net1417));
 sg13g2_nor2_1 _05364_ (.A(_01377_),
    .B(_01408_),
    .Y(_00066_));
 sg13g2_and3_2 _05365_ (.X(_01409_),
    .A(net3341),
    .B(net3691),
    .C(net1417));
 sg13g2_a21oi_1 _05366_ (.A1(\ram_spi_if.cycle_counter[1] ),
    .A2(net1417),
    .Y(_01410_),
    .B1(net3341));
 sg13g2_nor3_1 _05367_ (.A(_01377_),
    .B(_01409_),
    .C(net3342),
    .Y(_00067_));
 sg13g2_o21ai_1 _05368_ (.B1(_01376_),
    .Y(_01411_),
    .A1(net3496),
    .A2(_01409_));
 sg13g2_a21oi_1 _05369_ (.A1(net3496),
    .A2(_01409_),
    .Y(_00068_),
    .B1(_01411_));
 sg13g2_nand3_1 _05370_ (.B(net3496),
    .C(_01409_),
    .A(net3461),
    .Y(_01412_));
 sg13g2_nand2_1 _05371_ (.Y(_01413_),
    .A(_01376_),
    .B(_01412_));
 sg13g2_a21oi_1 _05372_ (.A1(\ram_spi_if.cycle_counter[3] ),
    .A2(_01409_),
    .Y(_01414_),
    .B1(net3461));
 sg13g2_nor2_1 _05373_ (.A(_01413_),
    .B(net3462),
    .Y(_00069_));
 sg13g2_nor2_2 _05374_ (.A(\ram_spi_if.cycle_counter[5] ),
    .B(_01377_),
    .Y(_01415_));
 sg13g2_nand2_1 _05375_ (.Y(_01416_),
    .A(_01340_),
    .B(_01376_));
 sg13g2_a22oi_1 _05376_ (.Y(_00070_),
    .B1(_01413_),
    .B2(_01416_),
    .A2(_01412_),
    .A1(_01340_));
 sg13g2_mux2_1 _05377_ (.A0(net3646),
    .A1(\cpu.i_rf_rdata[1] ),
    .S(net2584),
    .X(_00031_));
 sg13g2_mux2_1 _05378_ (.A0(net3673),
    .A1(net3574),
    .S(net2585),
    .X(_00042_));
 sg13g2_mux2_1 _05379_ (.A0(net3538),
    .A1(\cpu.i_rf_rdata[3] ),
    .S(net2586),
    .X(_00053_));
 sg13g2_mux2_1 _05380_ (.A0(net3357),
    .A1(\cpu.i_rf_rdata[4] ),
    .S(net2586),
    .X(_00054_));
 sg13g2_mux2_1 _05381_ (.A0(net3408),
    .A1(\cpu.i_rf_rdata[5] ),
    .S(net2586),
    .X(_00055_));
 sg13g2_mux2_1 _05382_ (.A0(net3365),
    .A1(\cpu.i_rf_rdata[6] ),
    .S(net2586),
    .X(_00056_));
 sg13g2_mux2_1 _05383_ (.A0(net3444),
    .A1(\cpu.i_rf_rdata[7] ),
    .S(net2586),
    .X(_00057_));
 sg13g2_mux2_1 _05384_ (.A0(net3482),
    .A1(\cpu.i_rf_rdata[8] ),
    .S(net2585),
    .X(_00058_));
 sg13g2_mux2_1 _05385_ (.A0(net3470),
    .A1(\cpu.i_rf_rdata[9] ),
    .S(net2585),
    .X(_00059_));
 sg13g2_mux2_1 _05386_ (.A0(net3355),
    .A1(\cpu.i_rf_rdata[10] ),
    .S(net2585),
    .X(_00060_));
 sg13g2_mux2_1 _05387_ (.A0(net3378),
    .A1(\cpu.i_rf_rdata[11] ),
    .S(net2585),
    .X(_00032_));
 sg13g2_mux2_1 _05388_ (.A0(net3430),
    .A1(\cpu.i_rf_rdata[12] ),
    .S(net2585),
    .X(_00033_));
 sg13g2_mux2_1 _05389_ (.A0(net3351),
    .A1(\cpu.i_rf_rdata[13] ),
    .S(net2585),
    .X(_00034_));
 sg13g2_mux2_1 _05390_ (.A0(net3523),
    .A1(\cpu.i_rf_rdata[14] ),
    .S(net2585),
    .X(_00035_));
 sg13g2_mux2_1 _05391_ (.A0(net3396),
    .A1(\cpu.i_rf_rdata[15] ),
    .S(net2584),
    .X(_00036_));
 sg13g2_mux2_1 _05392_ (.A0(net3353),
    .A1(\cpu.i_rf_rdata[16] ),
    .S(net2584),
    .X(_00037_));
 sg13g2_mux2_1 _05393_ (.A0(net3369),
    .A1(\cpu.i_rf_rdata[17] ),
    .S(net2584),
    .X(_00038_));
 sg13g2_mux2_1 _05394_ (.A0(net3338),
    .A1(\cpu.i_rf_rdata[18] ),
    .S(net2584),
    .X(_00039_));
 sg13g2_mux2_1 _05395_ (.A0(net3512),
    .A1(\cpu.i_rf_rdata[19] ),
    .S(net2584),
    .X(_00040_));
 sg13g2_mux2_1 _05396_ (.A0(\cpu.rf_ram_if.rdata1[20] ),
    .A1(net3502),
    .S(net2584),
    .X(_00041_));
 sg13g2_mux2_1 _05397_ (.A0(net3304),
    .A1(\cpu.i_rf_rdata[21] ),
    .S(net2584),
    .X(_00043_));
 sg13g2_mux2_1 _05398_ (.A0(net3401),
    .A1(\cpu.i_rf_rdata[22] ),
    .S(net2587),
    .X(_00044_));
 sg13g2_mux2_1 _05399_ (.A0(net3604),
    .A1(\cpu.i_rf_rdata[23] ),
    .S(net2583),
    .X(_00045_));
 sg13g2_mux2_1 _05400_ (.A0(net3371),
    .A1(\cpu.i_rf_rdata[24] ),
    .S(net2583),
    .X(_00046_));
 sg13g2_mux2_1 _05401_ (.A0(net3405),
    .A1(\cpu.i_rf_rdata[25] ),
    .S(net2583),
    .X(_00047_));
 sg13g2_mux2_1 _05402_ (.A0(net3446),
    .A1(\cpu.i_rf_rdata[26] ),
    .S(net2581),
    .X(_00048_));
 sg13g2_mux2_1 _05403_ (.A0(net3468),
    .A1(\cpu.i_rf_rdata[27] ),
    .S(net2582),
    .X(_00049_));
 sg13g2_mux2_1 _05404_ (.A0(net3424),
    .A1(\cpu.i_rf_rdata[28] ),
    .S(net2582),
    .X(_00050_));
 sg13g2_mux2_1 _05405_ (.A0(net3412),
    .A1(\cpu.i_rf_rdata[29] ),
    .S(net2581),
    .X(_00051_));
 sg13g2_mux2_1 _05406_ (.A0(net3414),
    .A1(\cpu.i_rf_rdata[30] ),
    .S(net2581),
    .X(_00052_));
 sg13g2_mux2_1 _05407_ (.A0(\cpu.rf_ram_if.rdata0[1] ),
    .A1(net3644),
    .S(\cpu.rf_ram_if.rtrig0 ),
    .X(_00000_));
 sg13g2_mux2_1 _05408_ (.A0(\cpu.i_rf_rdata[1] ),
    .A1(net3656),
    .S(net2380),
    .X(_00011_));
 sg13g2_mux2_1 _05409_ (.A0(net3574),
    .A1(\cpu.rf_ram_if.rdata0[3] ),
    .S(net2382),
    .X(_00022_));
 sg13g2_mux2_1 _05410_ (.A0(\cpu.i_rf_rdata[3] ),
    .A1(net3498),
    .S(net2382),
    .X(_00024_));
 sg13g2_mux2_1 _05411_ (.A0(\cpu.i_rf_rdata[4] ),
    .A1(net3359),
    .S(net2381),
    .X(_00025_));
 sg13g2_mux2_1 _05412_ (.A0(\cpu.i_rf_rdata[5] ),
    .A1(net3375),
    .S(net2382),
    .X(_00026_));
 sg13g2_mux2_1 _05413_ (.A0(\cpu.i_rf_rdata[6] ),
    .A1(net3327),
    .S(net2382),
    .X(_00027_));
 sg13g2_mux2_1 _05414_ (.A0(\cpu.i_rf_rdata[7] ),
    .A1(net3504),
    .S(net2382),
    .X(_00028_));
 sg13g2_mux2_1 _05415_ (.A0(\cpu.i_rf_rdata[8] ),
    .A1(net3452),
    .S(net2381),
    .X(_00029_));
 sg13g2_mux2_1 _05416_ (.A0(\cpu.i_rf_rdata[9] ),
    .A1(net3422),
    .S(net2381),
    .X(_00030_));
 sg13g2_mux2_1 _05417_ (.A0(\cpu.i_rf_rdata[10] ),
    .A1(net3394),
    .S(net2381),
    .X(_00001_));
 sg13g2_mux2_1 _05418_ (.A0(\cpu.i_rf_rdata[11] ),
    .A1(net3448),
    .S(net2381),
    .X(_00002_));
 sg13g2_mux2_1 _05419_ (.A0(\cpu.i_rf_rdata[12] ),
    .A1(net3416),
    .S(net2381),
    .X(_00003_));
 sg13g2_mux2_1 _05420_ (.A0(\cpu.i_rf_rdata[13] ),
    .A1(net3330),
    .S(net2381),
    .X(_00004_));
 sg13g2_mux2_1 _05421_ (.A0(\cpu.i_rf_rdata[14] ),
    .A1(net3530),
    .S(net2381),
    .X(_00005_));
 sg13g2_mux2_1 _05422_ (.A0(\cpu.i_rf_rdata[15] ),
    .A1(net3466),
    .S(net2380),
    .X(_00006_));
 sg13g2_mux2_1 _05423_ (.A0(\cpu.i_rf_rdata[16] ),
    .A1(net3384),
    .S(net2380),
    .X(_00007_));
 sg13g2_mux2_1 _05424_ (.A0(\cpu.i_rf_rdata[17] ),
    .A1(net3347),
    .S(net2380),
    .X(_00008_));
 sg13g2_mux2_1 _05425_ (.A0(\cpu.i_rf_rdata[18] ),
    .A1(net3349),
    .S(net2380),
    .X(_00009_));
 sg13g2_mux2_1 _05426_ (.A0(\cpu.i_rf_rdata[19] ),
    .A1(net3525),
    .S(net2380),
    .X(_00010_));
 sg13g2_mux2_1 _05427_ (.A0(\cpu.i_rf_rdata[20] ),
    .A1(net1404),
    .S(net2380),
    .X(_00012_));
 sg13g2_mux2_1 _05428_ (.A0(\cpu.i_rf_rdata[21] ),
    .A1(net3760),
    .S(net2380),
    .X(_00013_));
 sg13g2_mux2_1 _05429_ (.A0(\cpu.i_rf_rdata[22] ),
    .A1(net3427),
    .S(net2383),
    .X(_00014_));
 sg13g2_mux2_1 _05430_ (.A0(\cpu.i_rf_rdata[23] ),
    .A1(net3572),
    .S(net2379),
    .X(_00015_));
 sg13g2_mux2_1 _05431_ (.A0(\cpu.i_rf_rdata[24] ),
    .A1(net3332),
    .S(net2379),
    .X(_00016_));
 sg13g2_mux2_1 _05432_ (.A0(\cpu.i_rf_rdata[25] ),
    .A1(net3410),
    .S(net2379),
    .X(_00017_));
 sg13g2_mux2_1 _05433_ (.A0(\cpu.i_rf_rdata[26] ),
    .A1(net3459),
    .S(net2378),
    .X(_00018_));
 sg13g2_mux2_1 _05434_ (.A0(\cpu.i_rf_rdata[27] ),
    .A1(net3442),
    .S(net2378),
    .X(_00019_));
 sg13g2_mux2_1 _05435_ (.A0(\cpu.i_rf_rdata[28] ),
    .A1(net3345),
    .S(net2378),
    .X(_00020_));
 sg13g2_mux2_1 _05436_ (.A0(\cpu.i_rf_rdata[29] ),
    .A1(net3389),
    .S(net2377),
    .X(_00021_));
 sg13g2_mux2_1 _05437_ (.A0(\cpu.i_rf_rdata[30] ),
    .A1(net3403),
    .S(net2377),
    .X(_00023_));
 sg13g2_nor4_1 _05438_ (.A(net3364),
    .B(net3439),
    .C(net3492),
    .D(net3334),
    .Y(_01417_));
 sg13g2_or4_1 _05439_ (.A(\cpu.cpu.state.cnt_r[1] ),
    .B(\cpu.cpu.state.cnt_r[0] ),
    .C(\cpu.cpu.state.cnt_r[3] ),
    .D(\cpu.cpu.state.cnt_r[2] ),
    .X(_01418_));
 sg13g2_and2_1 _05440_ (.A(net2575),
    .B(\cpu.cpu.bufreg.i_sh_signed ),
    .X(_01419_));
 sg13g2_nor4_1 _05441_ (.A(net2569),
    .B(net3660),
    .C(net2574),
    .D(_01419_),
    .Y(_01420_));
 sg13g2_and2_1 _05442_ (.A(\cpu.cpu.alu.i_rs1 [0]),
    .B(net3764),
    .X(_01421_));
 sg13g2_xor2_1 _05443_ (.B(net3764),
    .A(\cpu.cpu.alu.i_rs1 [0]),
    .X(_01422_));
 sg13g2_nand2b_2 _05444_ (.Y(_01423_),
    .B(net2575),
    .A_N(net2579));
 sg13g2_nor3_1 _05445_ (.A(net2578),
    .B(net2579),
    .C(\cpu.cpu.decode.opcode[1] ),
    .Y(_01424_));
 sg13g2_nand3_1 _05446_ (.B(\cpu.cpu.state.o_cnt[2] ),
    .C(net3697),
    .A(net3492),
    .Y(_01425_));
 sg13g2_nand3_1 _05447_ (.B(\cpu.cpu.state.o_cnt[2] ),
    .C(\cpu.cpu.bufreg2.i_bytecnt[0] ),
    .A(\cpu.cpu.bufreg2.i_bytecnt[1] ),
    .Y(_01426_));
 sg13g2_nor2_2 _05448_ (.A(_01347_),
    .B(_01425_),
    .Y(_01427_));
 sg13g2_or2_1 _05449_ (.X(_01428_),
    .B(_01425_),
    .A(_01347_));
 sg13g2_a21oi_1 _05450_ (.A1(net2575),
    .A2(_01424_),
    .Y(_01429_),
    .B1(\cpu.cpu.immdec.gen_immdec_w_eq_1.imm24_20[0] ));
 sg13g2_nor4_1 _05451_ (.A(net2578),
    .B(\cpu.cpu.immdec.gen_immdec_w_eq_1.imm11_7[0] ),
    .C(\cpu.cpu.decode.opcode[1] ),
    .D(_01423_),
    .Y(_01430_));
 sg13g2_nand3_1 _05452_ (.B(net2577),
    .C(net2568),
    .A(net2573),
    .Y(_01431_));
 sg13g2_nand2_2 _05453_ (.Y(_01432_),
    .A(\cpu.cpu.immdec.gen_immdec_w_eq_1.imm31 ),
    .B(_01431_));
 sg13g2_nor3_2 _05454_ (.A(_01427_),
    .B(_01429_),
    .C(_01430_),
    .Y(_01433_));
 sg13g2_nor2_2 _05455_ (.A(_01428_),
    .B(_01432_),
    .Y(_01434_));
 sg13g2_nor3_1 _05456_ (.A(net2575),
    .B(_01433_),
    .C(_01434_),
    .Y(_01435_));
 sg13g2_or3_1 _05457_ (.A(net2575),
    .B(_01433_),
    .C(_01434_),
    .X(_01436_));
 sg13g2_nand2b_1 _05458_ (.Y(_01437_),
    .B(\cpu.rf_ram_if.rdata1[0] ),
    .A_N(net2581));
 sg13g2_nand2_1 _05459_ (.Y(_01438_),
    .A(net2582),
    .B(\cpu.i_rf_rdata[0] ));
 sg13g2_and3_1 _05460_ (.X(_01439_),
    .A(net2575),
    .B(_01437_),
    .C(_01438_));
 sg13g2_nand3_1 _05461_ (.B(_01437_),
    .C(_01438_),
    .A(net2576),
    .Y(_01440_));
 sg13g2_nor2_1 _05462_ (.A(_01435_),
    .B(_01439_),
    .Y(_01441_));
 sg13g2_nand3b_1 _05463_ (.B(_01436_),
    .C(_01440_),
    .Y(_01442_),
    .A_N(_01420_));
 sg13g2_o21ai_1 _05464_ (.B1(_01420_),
    .Y(_01443_),
    .A1(_01435_),
    .A2(_01439_));
 sg13g2_and2_1 _05465_ (.A(_01442_),
    .B(_01443_),
    .X(_01444_));
 sg13g2_and3_1 _05466_ (.X(_01445_),
    .A(_01422_),
    .B(_01442_),
    .C(_01443_));
 sg13g2_nor3_1 _05467_ (.A(net2566),
    .B(net3765),
    .C(_01445_),
    .Y(_01446_));
 sg13g2_a21oi_1 _05468_ (.A1(net2566),
    .A2(_01420_),
    .Y(_00061_),
    .B1(_01446_));
 sg13g2_nor2_1 _05469_ (.A(\ram_spi_if.cycle_counter[5] ),
    .B(\ram_spi_if.cycle_counter[4] ),
    .Y(_01447_));
 sg13g2_nor4_1 _05470_ (.A(\ram_spi_if.cycle_counter[3] ),
    .B(\ram_spi_if.cycle_counter[2] ),
    .C(\ram_spi_if.cycle_counter[1] ),
    .D(\ram_spi_if.cycle_counter[0] ),
    .Y(_01448_));
 sg13g2_nand2_1 _05471_ (.Y(_01449_),
    .A(clknet_1_0__leaf_clk),
    .B(_01376_));
 sg13g2_a21oi_1 _05472_ (.A1(_01447_),
    .A2(_01448_),
    .Y(\ram_spi_if.spi_clk ),
    .B1(_01449_));
 sg13g2_nor2_1 _05473_ (.A(net2574),
    .B(net2580),
    .Y(_01450_));
 sg13g2_nor2b_1 _05474_ (.A(net2568),
    .B_N(net2569),
    .Y(_01451_));
 sg13g2_o21ai_1 _05475_ (.B1(_01450_),
    .Y(_01452_),
    .A1(_01387_),
    .A2(_01451_));
 sg13g2_nand2b_1 _05476_ (.Y(_01453_),
    .B(net2577),
    .A_N(net2579));
 sg13g2_nor2_1 _05477_ (.A(net2572),
    .B(_01453_),
    .Y(_01454_));
 sg13g2_a21oi_2 _05478_ (.B1(net3720),
    .Y(_01455_),
    .A2(_01452_),
    .A1(net2577));
 sg13g2_a21oi_1 _05479_ (.A1(net2572),
    .A2(_01345_),
    .Y(_01456_),
    .B1(_01455_));
 sg13g2_nor2_1 _05480_ (.A(net2567),
    .B(_01456_),
    .Y(_01457_));
 sg13g2_nand2b_2 _05481_ (.Y(_01458_),
    .B(net2577),
    .A_N(net2570));
 sg13g2_a221oi_1 _05482_ (.B2(net2577),
    .C1(\cpu.cpu.state.init_done ),
    .B1(_01452_),
    .A1(net2568),
    .Y(_01459_),
    .A2(_01427_));
 sg13g2_nor2_1 _05483_ (.A(_01458_),
    .B(_01459_),
    .Y(_01460_));
 sg13g2_o21ai_1 _05484_ (.B1(net3450),
    .Y(_01461_),
    .A1(_01458_),
    .A2(_01459_));
 sg13g2_or2_1 _05485_ (.X(_01462_),
    .B(\cpu.arbiter.i_wb_cpu_dbus_dat[25] ),
    .A(\cpu.arbiter.i_wb_cpu_dbus_dat[24] ));
 sg13g2_nor4_1 _05486_ (.A(\cpu.arbiter.i_wb_cpu_dbus_dat[26] ),
    .B(\cpu.arbiter.i_wb_cpu_dbus_dat[27] ),
    .C(\cpu.arbiter.i_wb_cpu_dbus_dat[24] ),
    .D(\cpu.arbiter.i_wb_cpu_dbus_dat[25] ),
    .Y(_01463_));
 sg13g2_nand2_1 _05487_ (.Y(_01464_),
    .A(_01351_),
    .B(_01463_));
 sg13g2_xnor2_1 _05488_ (.Y(_01465_),
    .A(_01352_),
    .B(_01464_));
 sg13g2_or3_1 _05489_ (.A(_01458_),
    .B(_01459_),
    .C(_01465_),
    .X(_01466_));
 sg13g2_nand2_1 _05490_ (.Y(_01467_),
    .A(_01461_),
    .B(_01466_));
 sg13g2_nand3_1 _05491_ (.B(_01461_),
    .C(_01466_),
    .A(_01346_),
    .Y(_01468_));
 sg13g2_nor2_1 _05492_ (.A(_01335_),
    .B(_01458_),
    .Y(_01469_));
 sg13g2_a21oi_2 _05493_ (.B1(_01457_),
    .Y(_01470_),
    .A2(_01469_),
    .A1(_01468_));
 sg13g2_inv_1 _05494_ (.Y(_01471_),
    .A(net2330));
 sg13g2_nand2_1 _05495_ (.Y(_01472_),
    .A(net2574),
    .B(\cpu.cpu.decode.opcode[1] ));
 sg13g2_nor2b_1 _05496_ (.A(net2579),
    .B_N(net2573),
    .Y(_01473_));
 sg13g2_nand2b_1 _05497_ (.Y(_01474_),
    .B(net2572),
    .A_N(net2579));
 sg13g2_nand3_1 _05498_ (.B(_01472_),
    .C(_01474_),
    .A(\cpu.cpu.alu.i_rs1 [0]),
    .Y(_01475_));
 sg13g2_nand4_1 _05499_ (.B(net3600),
    .C(_01472_),
    .A(\cpu.cpu.alu.i_rs1 [0]),
    .Y(_01476_),
    .D(_01474_));
 sg13g2_nor3_1 _05500_ (.A(\cpu.cpu.bufreg2.i_bytecnt[1] ),
    .B(\cpu.cpu.state.o_cnt[2] ),
    .C(\cpu.cpu.bufreg2.i_bytecnt[0] ),
    .Y(_01477_));
 sg13g2_and2_1 _05501_ (.A(\cpu.cpu.state.cnt_r[0] ),
    .B(_01477_),
    .X(_01478_));
 sg13g2_xnor2_1 _05502_ (.Y(_01479_),
    .A(net2580),
    .B(\cpu.cpu.decode.opcode[1] ));
 sg13g2_and3_1 _05503_ (.X(_01480_),
    .A(net2574),
    .B(_01478_),
    .C(_01479_));
 sg13g2_o21ai_1 _05504_ (.B1(_01345_),
    .Y(_01481_),
    .A1(_01433_),
    .A2(_01434_));
 sg13g2_xor2_1 _05505_ (.B(_01475_),
    .A(net3600),
    .X(_01482_));
 sg13g2_or3_1 _05506_ (.A(_01480_),
    .B(_01481_),
    .C(_01482_),
    .X(_01483_));
 sg13g2_a21oi_1 _05507_ (.A1(net3601),
    .A2(_01483_),
    .Y(_00062_),
    .B1(net2330));
 sg13g2_nor2_2 _05508_ (.A(net2566),
    .B(net2376),
    .Y(_01484_));
 sg13g2_or2_1 _05509_ (.X(_01485_),
    .B(net2376),
    .A(net2567));
 sg13g2_nand3_1 _05510_ (.B(net2578),
    .C(\cpu.cpu.decode.co_ebreak ),
    .A(net2573),
    .Y(_01486_));
 sg13g2_nor2_1 _05511_ (.A(net2573),
    .B(net2575),
    .Y(_01487_));
 sg13g2_o21ai_1 _05512_ (.B1(_01486_),
    .Y(_01488_),
    .A1(net2572),
    .A2(net2575));
 sg13g2_a21o_1 _05513_ (.A2(\cpu.cpu.decode.opcode[1] ),
    .A1(net2580),
    .B1(_01488_),
    .X(_01489_));
 sg13g2_o21ai_1 _05514_ (.B1(\cpu.cpu.ctrl.pc [0]),
    .Y(_01490_),
    .A1(_01424_),
    .A2(_01489_));
 sg13g2_xnor2_1 _05515_ (.Y(_01491_),
    .A(_01370_),
    .B(_01490_));
 sg13g2_nand2b_1 _05516_ (.Y(_01492_),
    .B(net2579),
    .A_N(net2574));
 sg13g2_or2_1 _05517_ (.X(_01493_),
    .B(_01492_),
    .A(_01345_));
 sg13g2_nand3b_1 _05518_ (.B(_01493_),
    .C(\cpu.cpu.bufreg.data[0] ),
    .Y(_01494_),
    .A_N(net2330));
 sg13g2_a21oi_1 _05519_ (.A1(\cpu.cpu.state.o_cnt[2] ),
    .A2(\cpu.cpu.bufreg2.i_bytecnt[0] ),
    .Y(_01495_),
    .B1(\cpu.cpu.bufreg2.i_bytecnt[1] ));
 sg13g2_nor2_1 _05520_ (.A(_01493_),
    .B(_01495_),
    .Y(_01496_));
 sg13g2_o21ai_1 _05521_ (.B1(_01496_),
    .Y(_01497_),
    .A1(_01433_),
    .A2(_01434_));
 sg13g2_a21o_1 _05522_ (.A2(_01497_),
    .A1(_01494_),
    .B1(_01491_),
    .X(_01498_));
 sg13g2_o21ai_1 _05523_ (.B1(_01498_),
    .Y(_01499_),
    .A1(_01370_),
    .A2(_01490_));
 sg13g2_and2_1 _05524_ (.A(_01484_),
    .B(net3763),
    .X(_00064_));
 sg13g2_nand2_1 _05525_ (.Y(_01500_),
    .A(net3432),
    .B(\cpu.cpu.ctrl.pc [0]));
 sg13g2_xor2_1 _05526_ (.B(\cpu.cpu.ctrl.pc [0]),
    .A(net3432),
    .X(_01501_));
 sg13g2_nand3_1 _05527_ (.B(_01477_),
    .C(_01501_),
    .A(net3334),
    .Y(_01502_));
 sg13g2_a21oi_1 _05528_ (.A1(net3433),
    .A2(_01502_),
    .Y(_00063_),
    .B1(_01485_));
 sg13g2_nand3_1 _05529_ (.B(_01494_),
    .C(_01497_),
    .A(_01491_),
    .Y(_01503_));
 sg13g2_nand3b_1 _05530_ (.B(_01498_),
    .C(_01503_),
    .Y(_01504_),
    .A_N(_01478_));
 sg13g2_nand3_1 _05531_ (.B(_01451_),
    .C(_01478_),
    .A(\cpu.cpu.alu.cmp_r ),
    .Y(_01505_));
 sg13g2_o21ai_1 _05532_ (.B1(_01505_),
    .Y(_01506_),
    .A1(_01341_),
    .A2(net2330));
 sg13g2_xnor2_1 _05533_ (.Y(_01507_),
    .A(_01422_),
    .B(_01444_));
 sg13g2_nor4_1 _05534_ (.A(net2569),
    .B(\cpu.cpu.bne_or_bge ),
    .C(net2568),
    .D(_01507_),
    .Y(_01508_));
 sg13g2_nand3_1 _05535_ (.B(_01436_),
    .C(_01440_),
    .A(\cpu.cpu.alu.i_rs1 [0]),
    .Y(_01509_));
 sg13g2_a21o_1 _05536_ (.A2(_01440_),
    .A1(_01436_),
    .B1(\cpu.cpu.alu.i_rs1 [0]),
    .X(_01510_));
 sg13g2_nand3_1 _05537_ (.B(_01509_),
    .C(_01510_),
    .A(_01342_),
    .Y(_01511_));
 sg13g2_nand3_1 _05538_ (.B(\cpu.cpu.alu.i_rs1 [0]),
    .C(_01441_),
    .A(net2569),
    .Y(_01512_));
 sg13g2_a21oi_1 _05539_ (.A1(_01511_),
    .A2(_01512_),
    .Y(_01513_),
    .B1(_01346_));
 sg13g2_or3_1 _05540_ (.A(_01506_),
    .B(_01508_),
    .C(_01513_),
    .X(_01514_));
 sg13g2_a21oi_1 _05541_ (.A1(_01342_),
    .A2(\cpu.cpu.bufreg2.i_bytecnt[0] ),
    .Y(_01515_),
    .B1(\cpu.cpu.bufreg2.i_bytecnt[1] ));
 sg13g2_nor2_1 _05542_ (.A(net2569),
    .B(_01515_),
    .Y(_01516_));
 sg13g2_nand2_1 _05543_ (.Y(_01517_),
    .A(net2993),
    .B(_01516_));
 sg13g2_mux4_1 _05544_ (.S0(\cpu.cpu.bufreg.data[0] ),
    .A0(\cpu.arbiter.i_wb_cpu_dbus_dat[0] ),
    .A1(\cpu.arbiter.i_wb_cpu_dbus_dat[8] ),
    .A2(\cpu.arbiter.i_wb_cpu_dbus_dat[16] ),
    .A3(\cpu.arbiter.i_wb_cpu_dbus_dat[24] ),
    .S1(\cpu.cpu.bufreg.data[1] ),
    .X(_01518_));
 sg13g2_o21ai_1 _05545_ (.B1(_01518_),
    .Y(_01519_),
    .A1(net2570),
    .A2(_01515_));
 sg13g2_a21o_1 _05546_ (.A2(_01477_),
    .A1(\cpu.cpu.state.cnt_r[2] ),
    .B1(_01501_),
    .X(_01520_));
 sg13g2_and2_1 _05547_ (.A(_01502_),
    .B(_01520_),
    .X(_01521_));
 sg13g2_o21ai_1 _05548_ (.B1(_01519_),
    .Y(_01522_),
    .A1(net2568),
    .A2(_01517_));
 sg13g2_inv_1 _05549_ (.Y(_01523_),
    .A(_01522_));
 sg13g2_nand3_1 _05550_ (.B(net2580),
    .C(_01521_),
    .A(net2572),
    .Y(_01524_));
 sg13g2_o21ai_1 _05551_ (.B1(_01524_),
    .Y(_01525_),
    .A1(net2580),
    .A2(_01523_));
 sg13g2_a22oi_1 _05552_ (.Y(_01526_),
    .B1(_01525_),
    .B2(_01453_),
    .A2(_01514_),
    .A1(_01454_));
 sg13g2_o21ai_1 _05553_ (.B1(_01526_),
    .Y(\cpu.cpu.o_wdata0 [0]),
    .A1(_01493_),
    .A2(_01504_));
 sg13g2_nand2_2 _05554_ (.Y(_01527_),
    .A(net2581),
    .B(\cpu.rf_ram_if.wen0_r ));
 sg13g2_nor2_2 _05555_ (.A(net2588),
    .B(_01527_),
    .Y(_01528_));
 sg13g2_nand2_1 _05556_ (.Y(_01529_),
    .A(\cpu.cpu.immdec.gen_immdec_w_eq_1.imm11_7[2] ),
    .B(_01528_));
 sg13g2_a22oi_1 _05557_ (.Y(_01530_),
    .B1(_01366_),
    .B2(net2377),
    .A2(\cpu.rf_ram_if.wen0_r ),
    .A1(net2581));
 sg13g2_o21ai_1 _05558_ (.B1(_01530_),
    .Y(_01531_),
    .A1(\cpu.cpu.immdec.gen_immdec_w_eq_1.imm24_20[2] ),
    .A2(net2377));
 sg13g2_and2_1 _05559_ (.A(_01529_),
    .B(_01531_),
    .X(_01532_));
 sg13g2_nand2_2 _05560_ (.Y(_01533_),
    .A(_01529_),
    .B(_01531_));
 sg13g2_mux2_1 _05561_ (.A0(\cpu.cpu.immdec.gen_immdec_w_eq_1.imm19_12_20[7] ),
    .A1(\cpu.cpu.immdec.gen_immdec_w_eq_1.imm24_20[3] ),
    .S(\cpu.rf_ram_if.rtrig0 ),
    .X(_01534_));
 sg13g2_a22oi_1 _05562_ (.Y(_01535_),
    .B1(_01534_),
    .B2(_01527_),
    .A2(_01528_),
    .A1(\cpu.cpu.immdec.gen_immdec_w_eq_1.imm11_7[3] ));
 sg13g2_o21ai_1 _05563_ (.B1(_01527_),
    .Y(_01536_),
    .A1(\cpu.cpu.immdec.gen_immdec_w_eq_1.imm24_20[4] ),
    .A2(net2377));
 sg13g2_a21oi_1 _05564_ (.A1(_01368_),
    .A2(net2377),
    .Y(_01537_),
    .B1(_01536_));
 sg13g2_a21oi_2 _05565_ (.B1(_01537_),
    .Y(_01538_),
    .A2(_01528_),
    .A1(\cpu.cpu.immdec.gen_immdec_w_eq_1.imm11_7[4] ));
 sg13g2_nand3_1 _05566_ (.B(_01535_),
    .C(_01538_),
    .A(_01532_),
    .Y(_01539_));
 sg13g2_nand2b_1 _05567_ (.Y(_01540_),
    .B(net2377),
    .A_N(\cpu.cpu.csr_imm [0]));
 sg13g2_a22oi_1 _05568_ (.Y(_01541_),
    .B1(\cpu.rf_ram_if.rtrig0 ),
    .B2(_01362_),
    .A2(\cpu.rf_ram_if.wen0_r ),
    .A1(net2582));
 sg13g2_a22oi_1 _05569_ (.Y(_01542_),
    .B1(_01540_),
    .B2(_01541_),
    .A2(_01528_),
    .A1(\cpu.cpu.immdec.gen_immdec_w_eq_1.imm11_7[0] ));
 sg13g2_o21ai_1 _05570_ (.B1(_01527_),
    .Y(_01543_),
    .A1(\cpu.cpu.immdec.gen_immdec_w_eq_1.imm24_20[1] ),
    .A2(net2378));
 sg13g2_a21oi_1 _05571_ (.A1(_01364_),
    .A2(net2378),
    .Y(_01544_),
    .B1(_01543_));
 sg13g2_a21oi_2 _05572_ (.B1(_01544_),
    .Y(_01545_),
    .A2(_01528_),
    .A1(\cpu.cpu.immdec.gen_immdec_w_eq_1.imm11_7[1] ));
 sg13g2_nor2_1 _05573_ (.A(_01542_),
    .B(_01545_),
    .Y(_01546_));
 sg13g2_nor3_2 _05574_ (.A(_01527_),
    .B(_01542_),
    .C(_01545_),
    .Y(_01547_));
 sg13g2_nand2b_2 _05575_ (.Y(_01548_),
    .B(_01547_),
    .A_N(net2307));
 sg13g2_nand2b_1 _05576_ (.Y(_01549_),
    .B(\cpu.rf_ram_if.wdata0_r[0] ),
    .A_N(net2593));
 sg13g2_nand2_1 _05577_ (.Y(_01550_),
    .A(net3032),
    .B(net2107));
 sg13g2_o21ai_1 _05578_ (.B1(_01550_),
    .Y(_00620_),
    .A1(net2107),
    .A2(net2560));
 sg13g2_nand2b_1 _05579_ (.Y(_01551_),
    .B(net1410),
    .A_N(net2588));
 sg13g2_nand2_1 _05580_ (.Y(_01552_),
    .A(net3121),
    .B(net2116));
 sg13g2_o21ai_1 _05581_ (.B1(_01552_),
    .Y(_00621_),
    .A1(net2110),
    .A2(net2557));
 sg13g2_nand2b_2 _05582_ (.Y(_01553_),
    .B(net1412),
    .A_N(net2591));
 sg13g2_nand2_1 _05583_ (.Y(_01554_),
    .A(net1730),
    .B(net2115));
 sg13g2_o21ai_1 _05584_ (.B1(_01554_),
    .Y(_00622_),
    .A1(net2116),
    .A2(net2554));
 sg13g2_nand2b_1 _05585_ (.Y(_01555_),
    .B(net1387),
    .A_N(net2590));
 sg13g2_nand2_1 _05586_ (.Y(_01556_),
    .A(net3211),
    .B(net2114));
 sg13g2_o21ai_1 _05587_ (.B1(_01556_),
    .Y(_00623_),
    .A1(net2115),
    .A2(net2544));
 sg13g2_nand2b_2 _05588_ (.Y(_01557_),
    .B(net1400),
    .A_N(net2591));
 sg13g2_nand2_1 _05589_ (.Y(_01558_),
    .A(net3036),
    .B(net2114));
 sg13g2_o21ai_1 _05590_ (.B1(_01558_),
    .Y(_00624_),
    .A1(net2115),
    .A2(net2538));
 sg13g2_nand2b_2 _05591_ (.Y(_01559_),
    .B(net1393),
    .A_N(net2591));
 sg13g2_nand2_1 _05592_ (.Y(_01560_),
    .A(net2667),
    .B(net2115));
 sg13g2_o21ai_1 _05593_ (.B1(_01560_),
    .Y(_00625_),
    .A1(net2115),
    .A2(net2534));
 sg13g2_nand2b_1 _05594_ (.Y(_01561_),
    .B(net1408),
    .A_N(net2591));
 sg13g2_nand2_1 _05595_ (.Y(_01562_),
    .A(net1719),
    .B(net2114));
 sg13g2_o21ai_1 _05596_ (.B1(_01562_),
    .Y(_00626_),
    .A1(net2114),
    .A2(net2528));
 sg13g2_nand2b_2 _05597_ (.Y(_01563_),
    .B(net1397),
    .A_N(net2590));
 sg13g2_nand2_1 _05598_ (.Y(_01564_),
    .A(net1502),
    .B(net2114));
 sg13g2_o21ai_1 _05599_ (.B1(_01564_),
    .Y(_00627_),
    .A1(net2114),
    .A2(net2523));
 sg13g2_nand2b_2 _05600_ (.Y(_01565_),
    .B(net1402),
    .A_N(net2590));
 sg13g2_nand2_1 _05601_ (.Y(_01566_),
    .A(net2949),
    .B(net2111));
 sg13g2_o21ai_1 _05602_ (.B1(_01566_),
    .Y(_00628_),
    .A1(net2111),
    .A2(net2518));
 sg13g2_nand2b_1 _05603_ (.Y(_01567_),
    .B(net1409),
    .A_N(net2590));
 sg13g2_nand2_1 _05604_ (.Y(_01568_),
    .A(net2850),
    .B(net2111));
 sg13g2_o21ai_1 _05605_ (.B1(_01568_),
    .Y(_00629_),
    .A1(net2111),
    .A2(net2513));
 sg13g2_nand2b_2 _05606_ (.Y(_01569_),
    .B(net1392),
    .A_N(net2590));
 sg13g2_nand2_1 _05607_ (.Y(_01570_),
    .A(net1468),
    .B(net2112));
 sg13g2_o21ai_1 _05608_ (.B1(_01570_),
    .Y(_00630_),
    .A1(net2112),
    .A2(net2507));
 sg13g2_nand2b_1 _05609_ (.Y(_01571_),
    .B(net1381),
    .A_N(net2590));
 sg13g2_nand2_1 _05610_ (.Y(_01572_),
    .A(net2744),
    .B(net2111));
 sg13g2_o21ai_1 _05611_ (.B1(_01572_),
    .Y(_00631_),
    .A1(net2111),
    .A2(net2502));
 sg13g2_nand2b_2 _05612_ (.Y(_01573_),
    .B(net1401),
    .A_N(net2590));
 sg13g2_nand2_1 _05613_ (.Y(_01574_),
    .A(net3165),
    .B(net2111));
 sg13g2_o21ai_1 _05614_ (.B1(_01574_),
    .Y(_00632_),
    .A1(net2111),
    .A2(net2496));
 sg13g2_nand2b_1 _05615_ (.Y(_01575_),
    .B(net1396),
    .A_N(net2590));
 sg13g2_nand2_1 _05616_ (.Y(_01576_),
    .A(net1564),
    .B(net2112));
 sg13g2_o21ai_1 _05617_ (.B1(_01576_),
    .Y(_00633_),
    .A1(net2112),
    .A2(net2492));
 sg13g2_nand2b_1 _05618_ (.Y(_01577_),
    .B(net1389),
    .A_N(net2589));
 sg13g2_nand2_1 _05619_ (.Y(_01578_),
    .A(net3015),
    .B(net2108));
 sg13g2_o21ai_1 _05620_ (.B1(_01578_),
    .Y(_00634_),
    .A1(net2108),
    .A2(net2486));
 sg13g2_nand2b_1 _05621_ (.Y(_01579_),
    .B(net1385),
    .A_N(net2589));
 sg13g2_nand2_1 _05622_ (.Y(_01580_),
    .A(net2868),
    .B(net2113));
 sg13g2_o21ai_1 _05623_ (.B1(_01580_),
    .Y(_00635_),
    .A1(net2113),
    .A2(net2481));
 sg13g2_nand2b_2 _05624_ (.Y(_01581_),
    .B(net1394),
    .A_N(net2589));
 sg13g2_nand2_1 _05625_ (.Y(_01582_),
    .A(net1565),
    .B(net2114));
 sg13g2_o21ai_1 _05626_ (.B1(_01582_),
    .Y(_00636_),
    .A1(net2114),
    .A2(net2478));
 sg13g2_nand2b_2 _05627_ (.Y(_01583_),
    .B(net1398),
    .A_N(net2589));
 sg13g2_nand2_1 _05628_ (.Y(_01584_),
    .A(net3298),
    .B(net2113));
 sg13g2_o21ai_1 _05629_ (.B1(_01584_),
    .Y(_00637_),
    .A1(net2113),
    .A2(net2470));
 sg13g2_nand2b_1 _05630_ (.Y(_01585_),
    .B(net1388),
    .A_N(net2589));
 sg13g2_nand2_1 _05631_ (.Y(_01586_),
    .A(net1655),
    .B(net2113));
 sg13g2_o21ai_1 _05632_ (.B1(_01586_),
    .Y(_00638_),
    .A1(net2113),
    .A2(net2465));
 sg13g2_nand2b_2 _05633_ (.Y(_01587_),
    .B(net1390),
    .A_N(net2589));
 sg13g2_nand2_1 _05634_ (.Y(_01588_),
    .A(net3158),
    .B(net2108));
 sg13g2_o21ai_1 _05635_ (.B1(_01588_),
    .Y(_00639_),
    .A1(net2108),
    .A2(net2463));
 sg13g2_nand2b_2 _05636_ (.Y(_01589_),
    .B(net1413),
    .A_N(net2589));
 sg13g2_nand2_1 _05637_ (.Y(_01590_),
    .A(net1683),
    .B(net2108));
 sg13g2_o21ai_1 _05638_ (.B1(_01590_),
    .Y(_00640_),
    .A1(net2108),
    .A2(net2455));
 sg13g2_nand2b_2 _05639_ (.Y(_01591_),
    .B(net1403),
    .A_N(net2592));
 sg13g2_nand2_1 _05640_ (.Y(_01592_),
    .A(net1614),
    .B(net2109));
 sg13g2_o21ai_1 _05641_ (.B1(_01592_),
    .Y(_00641_),
    .A1(net2109),
    .A2(net2450));
 sg13g2_nand2b_1 _05642_ (.Y(_01593_),
    .B(net1383),
    .A_N(net2592));
 sg13g2_nand2_1 _05643_ (.Y(_01594_),
    .A(net3123),
    .B(net2116));
 sg13g2_o21ai_1 _05644_ (.B1(_01594_),
    .Y(_00642_),
    .A1(net2116),
    .A2(net2445));
 sg13g2_nand2b_2 _05645_ (.Y(_01595_),
    .B(net1399),
    .A_N(net2593));
 sg13g2_nand2_1 _05646_ (.Y(_01596_),
    .A(net3037),
    .B(net2108));
 sg13g2_o21ai_1 _05647_ (.B1(_01596_),
    .Y(_00643_),
    .A1(net2108),
    .A2(net2439));
 sg13g2_nand2b_2 _05648_ (.Y(_01597_),
    .B(net1391),
    .A_N(net2589));
 sg13g2_nand2_1 _05649_ (.Y(_01598_),
    .A(net2857),
    .B(net2116));
 sg13g2_o21ai_1 _05650_ (.B1(_01598_),
    .Y(_00644_),
    .A1(net2116),
    .A2(net2436));
 sg13g2_nand2b_1 _05651_ (.Y(_01599_),
    .B(net1407),
    .A_N(net2593));
 sg13g2_nand2_1 _05652_ (.Y(_01600_),
    .A(net1627),
    .B(net2109));
 sg13g2_o21ai_1 _05653_ (.B1(_01600_),
    .Y(_00645_),
    .A1(net2109),
    .A2(net2429));
 sg13g2_nand2b_2 _05654_ (.Y(_01601_),
    .B(net1411),
    .A_N(net2588));
 sg13g2_nand2_1 _05655_ (.Y(_01602_),
    .A(net3090),
    .B(net2110));
 sg13g2_o21ai_1 _05656_ (.B1(_01602_),
    .Y(_00646_),
    .A1(net2110),
    .A2(net2425));
 sg13g2_nand2b_1 _05657_ (.Y(_01603_),
    .B(net1382),
    .A_N(net2588));
 sg13g2_nand2_1 _05658_ (.Y(_01604_),
    .A(net2910),
    .B(net2109));
 sg13g2_o21ai_1 _05659_ (.B1(_01604_),
    .Y(_00647_),
    .A1(net2109),
    .A2(net2418));
 sg13g2_nand2b_1 _05660_ (.Y(_01605_),
    .B(net1406),
    .A_N(net2588));
 sg13g2_nand2_1 _05661_ (.Y(_01606_),
    .A(net2617),
    .B(net2109));
 sg13g2_o21ai_1 _05662_ (.B1(_01606_),
    .Y(_00648_),
    .A1(net2109),
    .A2(net2413));
 sg13g2_nand2b_2 _05663_ (.Y(_01607_),
    .B(net1395),
    .A_N(net2588));
 sg13g2_nand2_1 _05664_ (.Y(_01608_),
    .A(net3265),
    .B(net2107));
 sg13g2_o21ai_1 _05665_ (.B1(_01608_),
    .Y(_00649_),
    .A1(net2107),
    .A2(net2410));
 sg13g2_nand2b_1 _05666_ (.Y(_01609_),
    .B(net1386),
    .A_N(net2588));
 sg13g2_nand2_1 _05667_ (.Y(_01610_),
    .A(net3039),
    .B(net2107));
 sg13g2_o21ai_1 _05668_ (.B1(_01610_),
    .Y(_00650_),
    .A1(net2107),
    .A2(net2403));
 sg13g2_nand2b_1 _05669_ (.Y(_01611_),
    .B(net1384),
    .A_N(net2588));
 sg13g2_nand2_1 _05670_ (.Y(_01612_),
    .A(net3164),
    .B(net2107));
 sg13g2_o21ai_1 _05671_ (.B1(_01612_),
    .Y(_00651_),
    .A1(net2107),
    .A2(net2397));
 sg13g2_and3_2 _05672_ (.X(_01613_),
    .A(net2325),
    .B(_01535_),
    .C(_01538_));
 sg13g2_nand3_1 _05673_ (.B(_01535_),
    .C(_01538_),
    .A(net2325),
    .Y(_01614_));
 sg13g2_and2_1 _05674_ (.A(_01542_),
    .B(_01545_),
    .X(_01615_));
 sg13g2_nor2b_2 _05675_ (.A(_01527_),
    .B_N(net2221),
    .Y(_01616_));
 sg13g2_nand2_1 _05676_ (.Y(_01617_),
    .A(_01613_),
    .B(_01616_));
 sg13g2_nand2_1 _05677_ (.Y(_01618_),
    .A(net1446),
    .B(net2056));
 sg13g2_o21ai_1 _05678_ (.B1(_01618_),
    .Y(_00652_),
    .A1(net2562),
    .A2(net2056));
 sg13g2_nand2_1 _05679_ (.Y(_01619_),
    .A(net2707),
    .B(net2058));
 sg13g2_o21ai_1 _05680_ (.B1(_01619_),
    .Y(_00653_),
    .A1(net2555),
    .A2(net2058));
 sg13g2_nand2_1 _05681_ (.Y(_01620_),
    .A(net3266),
    .B(net2062));
 sg13g2_o21ai_1 _05682_ (.B1(_01620_),
    .Y(_00654_),
    .A1(net2550),
    .A2(net2062));
 sg13g2_nand2_1 _05683_ (.Y(_01621_),
    .A(net1634),
    .B(net2061));
 sg13g2_o21ai_1 _05684_ (.B1(_01621_),
    .Y(_00655_),
    .A1(net2545),
    .A2(net2061));
 sg13g2_nand2_1 _05685_ (.Y(_01622_),
    .A(net1428),
    .B(net2061));
 sg13g2_o21ai_1 _05686_ (.B1(_01622_),
    .Y(_00656_),
    .A1(net2541),
    .A2(net2061));
 sg13g2_nand2_1 _05687_ (.Y(_01623_),
    .A(net1651),
    .B(net2061));
 sg13g2_o21ai_1 _05688_ (.B1(_01623_),
    .Y(_00657_),
    .A1(net2537),
    .A2(net2061));
 sg13g2_nand2_1 _05689_ (.Y(_01624_),
    .A(net3169),
    .B(net2063));
 sg13g2_o21ai_1 _05690_ (.B1(_01624_),
    .Y(_00658_),
    .A1(net2531),
    .A2(net2063));
 sg13g2_nand2_1 _05691_ (.Y(_01625_),
    .A(net3146),
    .B(net2061));
 sg13g2_o21ai_1 _05692_ (.B1(_01625_),
    .Y(_00659_),
    .A1(net2524),
    .A2(net2061));
 sg13g2_nand2_1 _05693_ (.Y(_01626_),
    .A(net2953),
    .B(net2060));
 sg13g2_o21ai_1 _05694_ (.B1(_01626_),
    .Y(_00660_),
    .A1(net2520),
    .A2(net2060));
 sg13g2_nand2_1 _05695_ (.Y(_01627_),
    .A(net2816),
    .B(net2060));
 sg13g2_o21ai_1 _05696_ (.B1(_01627_),
    .Y(_00661_),
    .A1(net2516),
    .A2(net2060));
 sg13g2_nand2_1 _05697_ (.Y(_01628_),
    .A(net2942),
    .B(net2060));
 sg13g2_o21ai_1 _05698_ (.B1(_01628_),
    .Y(_00662_),
    .A1(net2508),
    .A2(net2060));
 sg13g2_nand2_1 _05699_ (.Y(_01629_),
    .A(net3044),
    .B(net2059));
 sg13g2_o21ai_1 _05700_ (.B1(_01629_),
    .Y(_00663_),
    .A1(net2503),
    .A2(net2059));
 sg13g2_nand2_1 _05701_ (.Y(_01630_),
    .A(net3308),
    .B(net2060));
 sg13g2_o21ai_1 _05702_ (.B1(_01630_),
    .Y(_00664_),
    .A1(net2497),
    .A2(net2060));
 sg13g2_nand2_1 _05703_ (.Y(_01631_),
    .A(net3240),
    .B(net2059));
 sg13g2_o21ai_1 _05704_ (.B1(_01631_),
    .Y(_00665_),
    .A1(net2491),
    .A2(net2059));
 sg13g2_nand2_1 _05705_ (.Y(_01632_),
    .A(net2618),
    .B(net2056));
 sg13g2_o21ai_1 _05706_ (.B1(_01632_),
    .Y(_00666_),
    .A1(net2488),
    .A2(net2064));
 sg13g2_nand2_1 _05707_ (.Y(_01633_),
    .A(net2631),
    .B(net2059));
 sg13g2_o21ai_1 _05708_ (.B1(_01633_),
    .Y(_00667_),
    .A1(net2483),
    .A2(net2059));
 sg13g2_nand2_1 _05709_ (.Y(_01634_),
    .A(net1429),
    .B(net2062));
 sg13g2_o21ai_1 _05710_ (.B1(_01634_),
    .Y(_00668_),
    .A1(net2480),
    .A2(net2062));
 sg13g2_nand2_1 _05711_ (.Y(_01635_),
    .A(net2895),
    .B(net2056));
 sg13g2_o21ai_1 _05712_ (.B1(_01635_),
    .Y(_00669_),
    .A1(net2471),
    .A2(net2056));
 sg13g2_nand2_1 _05713_ (.Y(_01636_),
    .A(net1648),
    .B(net2059));
 sg13g2_o21ai_1 _05714_ (.B1(_01636_),
    .Y(_00670_),
    .A1(net2467),
    .A2(net2059));
 sg13g2_nand2_1 _05715_ (.Y(_01637_),
    .A(net1450),
    .B(net2055));
 sg13g2_o21ai_1 _05716_ (.B1(_01637_),
    .Y(_00671_),
    .A1(net2461),
    .A2(net2055));
 sg13g2_nand2_1 _05717_ (.Y(_01638_),
    .A(net2692),
    .B(net2056));
 sg13g2_o21ai_1 _05718_ (.B1(_01638_),
    .Y(_00672_),
    .A1(net2459),
    .A2(net2056));
 sg13g2_nand2_1 _05719_ (.Y(_01639_),
    .A(net2847),
    .B(net2058));
 sg13g2_o21ai_1 _05720_ (.B1(_01639_),
    .Y(_00673_),
    .A1(net2453),
    .A2(net2058));
 sg13g2_nand2_1 _05721_ (.Y(_01640_),
    .A(net3238),
    .B(net2062));
 sg13g2_o21ai_1 _05722_ (.B1(_01640_),
    .Y(_00674_),
    .A1(net2447),
    .A2(net2062));
 sg13g2_nand2_1 _05723_ (.Y(_01641_),
    .A(net3113),
    .B(net2057));
 sg13g2_o21ai_1 _05724_ (.B1(_01641_),
    .Y(_00675_),
    .A1(net2440),
    .A2(net2057));
 sg13g2_nand2_1 _05725_ (.Y(_01642_),
    .A(net2724),
    .B(net2062));
 sg13g2_o21ai_1 _05726_ (.B1(_01642_),
    .Y(_00676_),
    .A1(net2434),
    .A2(net2062));
 sg13g2_nand2_1 _05727_ (.Y(_01643_),
    .A(net1465),
    .B(net2057));
 sg13g2_o21ai_1 _05728_ (.B1(_01643_),
    .Y(_00677_),
    .A1(net2428),
    .A2(net2057));
 sg13g2_nand2_1 _05729_ (.Y(_01644_),
    .A(net1623),
    .B(net2058));
 sg13g2_o21ai_1 _05730_ (.B1(_01644_),
    .Y(_00678_),
    .A1(net2423),
    .A2(net2057));
 sg13g2_nand2_1 _05731_ (.Y(_01645_),
    .A(net3280),
    .B(net2057));
 sg13g2_o21ai_1 _05732_ (.B1(_01645_),
    .Y(_00679_),
    .A1(net2419),
    .A2(net2058));
 sg13g2_nand2_1 _05733_ (.Y(_01646_),
    .A(net2614),
    .B(net2057));
 sg13g2_o21ai_1 _05734_ (.B1(_01646_),
    .Y(_00680_),
    .A1(net2415),
    .A2(net2057));
 sg13g2_nand2_1 _05735_ (.Y(_01647_),
    .A(net2957),
    .B(net2055));
 sg13g2_o21ai_1 _05736_ (.B1(_01647_),
    .Y(_00681_),
    .A1(net2412),
    .A2(net2055));
 sg13g2_nand2_1 _05737_ (.Y(_01648_),
    .A(net2660),
    .B(net2055));
 sg13g2_o21ai_1 _05738_ (.B1(_01648_),
    .Y(_00682_),
    .A1(net2404),
    .A2(net2055));
 sg13g2_nand2_1 _05739_ (.Y(_01649_),
    .A(net2732),
    .B(net2055));
 sg13g2_o21ai_1 _05740_ (.B1(_01649_),
    .Y(_00683_),
    .A1(net2399),
    .A2(net2055));
 sg13g2_nor2_1 _05741_ (.A(\ram_spi_if.cycle_counter[3] ),
    .B(_01399_),
    .Y(_01650_));
 sg13g2_nand2_1 _05742_ (.Y(_01651_),
    .A(\cpu.cpu.state.init_done ),
    .B(net2567));
 sg13g2_nor3_1 _05743_ (.A(net2572),
    .B(net2577),
    .C(_01651_),
    .Y(_01652_));
 sg13g2_nor2_2 _05744_ (.A(\cpu.arbiter.i_wb_cpu_dbus_adr[31] ),
    .B(\cpu.arbiter.i_wb_cpu_dbus_adr[30] ),
    .Y(_01653_));
 sg13g2_or2_1 _05745_ (.X(_01654_),
    .B(\cpu.arbiter.i_wb_cpu_dbus_adr[30] ),
    .A(\cpu.arbiter.i_wb_cpu_dbus_adr[31] ));
 sg13g2_and2_1 _05746_ (.A(net2598),
    .B(\cpu.cpu.state.ibus_cyc ),
    .X(_01655_));
 sg13g2_nand2_2 _05747_ (.Y(_01656_),
    .A(net2598),
    .B(\cpu.cpu.state.ibus_cyc ));
 sg13g2_a21oi_1 _05748_ (.A1(_01652_),
    .A2(net2396),
    .Y(_01657_),
    .B1(net2393));
 sg13g2_nand3b_1 _05749_ (.B(net2594),
    .C(_01371_),
    .Y(_01658_),
    .A_N(net2595));
 sg13g2_and2_1 _05750_ (.A(\ram_spi_if.cycle_counter[5] ),
    .B(net2571),
    .X(_01659_));
 sg13g2_o21ai_1 _05751_ (.B1(\ram_spi_if.cycle_counter[3] ),
    .Y(_01660_),
    .A1(\cpu.cpu.bufreg.data[0] ),
    .A2(_01342_));
 sg13g2_a21oi_1 _05752_ (.A1(_01447_),
    .A2(_01660_),
    .Y(_01661_),
    .B1(net2571));
 sg13g2_a21oi_1 _05753_ (.A1(_01378_),
    .A2(_01659_),
    .Y(_01662_),
    .B1(_01661_));
 sg13g2_o21ai_1 _05754_ (.B1(_01447_),
    .Y(_01663_),
    .A1(_01397_),
    .A2(_01650_));
 sg13g2_o21ai_1 _05755_ (.B1(_01663_),
    .Y(_01664_),
    .A1(net3717),
    .A2(_01658_));
 sg13g2_a221oi_1 _05756_ (.B2(_01380_),
    .C1(_01664_),
    .B1(_01662_),
    .A1(_01407_),
    .Y(_01665_),
    .A2(_01657_));
 sg13g2_nor2b_1 _05757_ (.A(_01375_),
    .B_N(_01665_),
    .Y(_00684_));
 sg13g2_nand2_1 _05758_ (.Y(_01666_),
    .A(net2576),
    .B(net2391));
 sg13g2_a22oi_1 _05759_ (.Y(_01667_),
    .B1(_01396_),
    .B2(_01666_),
    .A2(_01373_),
    .A1(net2596));
 sg13g2_nand2b_2 _05760_ (.Y(_01668_),
    .B(net2595),
    .A_N(net2594));
 sg13g2_nor3_2 _05761_ (.A(net3725),
    .B(_01344_),
    .C(_01668_),
    .Y(_01669_));
 sg13g2_nand2_2 _05762_ (.Y(_01670_),
    .A(net2596),
    .B(_01396_));
 sg13g2_nand3_1 _05763_ (.B(_01667_),
    .C(_01670_),
    .A(_01399_),
    .Y(_01671_));
 sg13g2_nand2_1 _05764_ (.Y(_01672_),
    .A(_01665_),
    .B(_01671_));
 sg13g2_o21ai_1 _05765_ (.B1(_01672_),
    .Y(_00685_),
    .A1(_01343_),
    .A2(_01665_));
 sg13g2_nand2_2 _05766_ (.Y(_01673_),
    .A(net2595),
    .B(_01398_));
 sg13g2_a21oi_1 _05767_ (.A1(net2595),
    .A2(_01398_),
    .Y(_01674_),
    .B1(_01396_));
 sg13g2_nor2_1 _05768_ (.A(net3704),
    .B(_01665_),
    .Y(_01675_));
 sg13g2_a21oi_1 _05769_ (.A1(_01665_),
    .A2(_01674_),
    .Y(_00686_),
    .B1(net3705));
 sg13g2_nand2_1 _05770_ (.Y(_01676_),
    .A(_01379_),
    .B(_01658_));
 sg13g2_mux2_1 _05771_ (.A0(net3726),
    .A1(_01676_),
    .S(_01665_),
    .X(_00687_));
 sg13g2_nand2b_2 _05772_ (.Y(_01677_),
    .B(_01538_),
    .A_N(_01535_));
 sg13g2_nor2_2 _05773_ (.A(_01532_),
    .B(_01677_),
    .Y(_01678_));
 sg13g2_nand2b_1 _05774_ (.Y(_01679_),
    .B(net2325),
    .A_N(_01677_));
 sg13g2_nand2_2 _05775_ (.Y(_01680_),
    .A(_01547_),
    .B(_01678_));
 sg13g2_nand2_1 _05776_ (.Y(_01681_),
    .A(net3156),
    .B(net2046));
 sg13g2_o21ai_1 _05777_ (.B1(_01681_),
    .Y(_00688_),
    .A1(net2564),
    .A2(net2046));
 sg13g2_nand2_1 _05778_ (.Y(_01682_),
    .A(net3225),
    .B(net2048));
 sg13g2_o21ai_1 _05779_ (.B1(_01682_),
    .Y(_00689_),
    .A1(net2557),
    .A2(net2048));
 sg13g2_nand2_1 _05780_ (.Y(_01683_),
    .A(net3230),
    .B(net2052));
 sg13g2_o21ai_1 _05781_ (.B1(_01683_),
    .Y(_00690_),
    .A1(net2553),
    .A2(net2053));
 sg13g2_nand2_1 _05782_ (.Y(_01684_),
    .A(net2778),
    .B(net2053));
 sg13g2_o21ai_1 _05783_ (.B1(_01684_),
    .Y(_00691_),
    .A1(net2547),
    .A2(net2053));
 sg13g2_nand2_1 _05784_ (.Y(_01685_),
    .A(net2999),
    .B(net2052));
 sg13g2_o21ai_1 _05785_ (.B1(_01685_),
    .Y(_00692_),
    .A1(net2539),
    .A2(net2053));
 sg13g2_nand2_1 _05786_ (.Y(_01686_),
    .A(net1597),
    .B(net2053));
 sg13g2_o21ai_1 _05787_ (.B1(_01686_),
    .Y(_00693_),
    .A1(net2535),
    .A2(net2053));
 sg13g2_nand2_1 _05788_ (.Y(_01687_),
    .A(net3221),
    .B(net2054));
 sg13g2_o21ai_1 _05789_ (.B1(_01687_),
    .Y(_00694_),
    .A1(net2530),
    .A2(net2054));
 sg13g2_nand2_1 _05790_ (.Y(_01688_),
    .A(net2686),
    .B(net2053));
 sg13g2_o21ai_1 _05791_ (.B1(_01688_),
    .Y(_00695_),
    .A1(net2526),
    .A2(net2054));
 sg13g2_nand2_1 _05792_ (.Y(_01689_),
    .A(net3099),
    .B(net2051));
 sg13g2_o21ai_1 _05793_ (.B1(_01689_),
    .Y(_00696_),
    .A1(net2522),
    .A2(net2051));
 sg13g2_nand2_1 _05794_ (.Y(_01690_),
    .A(net2718),
    .B(net2051));
 sg13g2_o21ai_1 _05795_ (.B1(_01690_),
    .Y(_00697_),
    .A1(net2515),
    .A2(net2051));
 sg13g2_nand2_1 _05796_ (.Y(_01691_),
    .A(net1633),
    .B(net2050));
 sg13g2_o21ai_1 _05797_ (.B1(_01691_),
    .Y(_00698_),
    .A1(net2510),
    .A2(net2050));
 sg13g2_nand2_1 _05798_ (.Y(_01692_),
    .A(net3047),
    .B(net2050));
 sg13g2_o21ai_1 _05799_ (.B1(_01692_),
    .Y(_00699_),
    .A1(net2505),
    .A2(net2050));
 sg13g2_nand2_1 _05800_ (.Y(_01693_),
    .A(net1475),
    .B(net2051));
 sg13g2_o21ai_1 _05801_ (.B1(_01693_),
    .Y(_00700_),
    .A1(net2500),
    .A2(net2051));
 sg13g2_nand2_1 _05802_ (.Y(_01694_),
    .A(net3070),
    .B(net2052));
 sg13g2_o21ai_1 _05803_ (.B1(_01694_),
    .Y(_00701_),
    .A1(net2495),
    .A2(net2052));
 sg13g2_nand2_1 _05804_ (.Y(_01695_),
    .A(net2944),
    .B(net2049));
 sg13g2_o21ai_1 _05805_ (.B1(_01695_),
    .Y(_00702_),
    .A1(net2490),
    .A2(net2049));
 sg13g2_nand2_1 _05806_ (.Y(_01696_),
    .A(net3182),
    .B(net2046));
 sg13g2_o21ai_1 _05807_ (.B1(_01696_),
    .Y(_00703_),
    .A1(net2481),
    .A2(net2046));
 sg13g2_nand2_1 _05808_ (.Y(_01697_),
    .A(net2661),
    .B(net2050));
 sg13g2_o21ai_1 _05809_ (.B1(_01697_),
    .Y(_00704_),
    .A1(net2475),
    .A2(net2050));
 sg13g2_nand2_1 _05810_ (.Y(_01698_),
    .A(net1460),
    .B(net2046));
 sg13g2_o21ai_1 _05811_ (.B1(_01698_),
    .Y(_00705_),
    .A1(net2474),
    .A2(net2046));
 sg13g2_nand2_1 _05812_ (.Y(_01699_),
    .A(net3125),
    .B(net2050));
 sg13g2_o21ai_1 _05813_ (.B1(_01699_),
    .Y(_00706_),
    .A1(net2467),
    .A2(net2050));
 sg13g2_nand2_1 _05814_ (.Y(_01700_),
    .A(net2928),
    .B(net2045));
 sg13g2_o21ai_1 _05815_ (.B1(_01700_),
    .Y(_00707_),
    .A1(net2461),
    .A2(net2045));
 sg13g2_nand2_1 _05816_ (.Y(_01701_),
    .A(net3154),
    .B(net2046));
 sg13g2_o21ai_1 _05817_ (.B1(_01701_),
    .Y(_00708_),
    .A1(net2456),
    .A2(net2049));
 sg13g2_nand2_1 _05818_ (.Y(_01702_),
    .A(net3278),
    .B(net2048));
 sg13g2_o21ai_1 _05819_ (.B1(_01702_),
    .Y(_00709_),
    .A1(net2454),
    .A2(net2048));
 sg13g2_nand2_1 _05820_ (.Y(_01703_),
    .A(net1710),
    .B(net2052));
 sg13g2_o21ai_1 _05821_ (.B1(_01703_),
    .Y(_00710_),
    .A1(net2448),
    .A2(net2052));
 sg13g2_nand2_1 _05822_ (.Y(_01704_),
    .A(net2725),
    .B(net2047));
 sg13g2_o21ai_1 _05823_ (.B1(_01704_),
    .Y(_00711_),
    .A1(net2442),
    .A2(net2047));
 sg13g2_nand2_1 _05824_ (.Y(_01705_),
    .A(net3249),
    .B(net2052));
 sg13g2_o21ai_1 _05825_ (.B1(_01705_),
    .Y(_00712_),
    .A1(net2437),
    .A2(net2052));
 sg13g2_nand2_1 _05826_ (.Y(_01706_),
    .A(net3023),
    .B(net2047));
 sg13g2_o21ai_1 _05827_ (.B1(_01706_),
    .Y(_00713_),
    .A1(net2431),
    .A2(net2047));
 sg13g2_nand2_1 _05828_ (.Y(_01707_),
    .A(net2668),
    .B(net2047));
 sg13g2_o21ai_1 _05829_ (.B1(_01707_),
    .Y(_00714_),
    .A1(net2426),
    .A2(net2047));
 sg13g2_nand2_1 _05830_ (.Y(_01708_),
    .A(net3089),
    .B(net2048));
 sg13g2_o21ai_1 _05831_ (.B1(_01708_),
    .Y(_00715_),
    .A1(net2420),
    .A2(net2048));
 sg13g2_nand2_1 _05832_ (.Y(_01709_),
    .A(net3007),
    .B(net2047));
 sg13g2_o21ai_1 _05833_ (.B1(_01709_),
    .Y(_00716_),
    .A1(net2417),
    .A2(net2047));
 sg13g2_nand2_1 _05834_ (.Y(_01710_),
    .A(net2907),
    .B(net2045));
 sg13g2_o21ai_1 _05835_ (.B1(_01710_),
    .Y(_00717_),
    .A1(net2411),
    .A2(net2045));
 sg13g2_nand2_1 _05836_ (.Y(_01711_),
    .A(net2793),
    .B(net2045));
 sg13g2_o21ai_1 _05837_ (.B1(_01711_),
    .Y(_00718_),
    .A1(net2406),
    .A2(net2045));
 sg13g2_nand2_1 _05838_ (.Y(_01712_),
    .A(net2990),
    .B(net2045));
 sg13g2_o21ai_1 _05839_ (.B1(_01712_),
    .Y(_00719_),
    .A1(net2400),
    .A2(net2045));
 sg13g2_nor2_1 _05840_ (.A(_01533_),
    .B(_01677_),
    .Y(_01713_));
 sg13g2_or2_1 _05841_ (.X(_01714_),
    .B(_01677_),
    .A(net2325));
 sg13g2_nor2b_1 _05842_ (.A(_01542_),
    .B_N(_01545_),
    .Y(_01715_));
 sg13g2_nor2b_2 _05843_ (.A(_01527_),
    .B_N(net2186),
    .Y(_01716_));
 sg13g2_nand2_1 _05844_ (.Y(_01717_),
    .A(_01713_),
    .B(_01716_));
 sg13g2_nand2_1 _05845_ (.Y(_01718_),
    .A(net2918),
    .B(net2034));
 sg13g2_o21ai_1 _05846_ (.B1(_01718_),
    .Y(_00720_),
    .A1(net2564),
    .A2(net2034));
 sg13g2_nand2_1 _05847_ (.Y(_01719_),
    .A(net1547),
    .B(net2037));
 sg13g2_o21ai_1 _05848_ (.B1(_01719_),
    .Y(_00721_),
    .A1(net2556),
    .A2(net2037));
 sg13g2_nand2_1 _05849_ (.Y(_01720_),
    .A(net3049),
    .B(net2043));
 sg13g2_o21ai_1 _05850_ (.B1(_01720_),
    .Y(_00722_),
    .A1(net2550),
    .A2(net2043));
 sg13g2_nand2_1 _05851_ (.Y(_01721_),
    .A(net2934),
    .B(net2041));
 sg13g2_o21ai_1 _05852_ (.B1(_01721_),
    .Y(_00723_),
    .A1(net2544),
    .A2(net2041));
 sg13g2_nand2_1 _05853_ (.Y(_01722_),
    .A(net2739),
    .B(net2041));
 sg13g2_o21ai_1 _05854_ (.B1(_01722_),
    .Y(_00724_),
    .A1(net2540),
    .A2(net2041));
 sg13g2_nand2_1 _05855_ (.Y(_01723_),
    .A(net1546),
    .B(net2041));
 sg13g2_o21ai_1 _05856_ (.B1(_01723_),
    .Y(_00725_),
    .A1(net2533),
    .A2(net2041));
 sg13g2_nand2_1 _05857_ (.Y(_01724_),
    .A(net1529),
    .B(net2043));
 sg13g2_o21ai_1 _05858_ (.B1(_01724_),
    .Y(_00726_),
    .A1(net2528),
    .A2(net2042));
 sg13g2_nand2_1 _05859_ (.Y(_01725_),
    .A(net2819),
    .B(net2042));
 sg13g2_o21ai_1 _05860_ (.B1(_01725_),
    .Y(_00727_),
    .A1(net2523),
    .A2(net2042));
 sg13g2_nand2_1 _05861_ (.Y(_01726_),
    .A(net2881),
    .B(net2042));
 sg13g2_o21ai_1 _05862_ (.B1(_01726_),
    .Y(_00728_),
    .A1(net2518),
    .A2(net2042));
 sg13g2_nand2_1 _05863_ (.Y(_01727_),
    .A(net1498),
    .B(net2040));
 sg13g2_o21ai_1 _05864_ (.B1(_01727_),
    .Y(_00729_),
    .A1(net2512),
    .A2(net2040));
 sg13g2_nand2_1 _05865_ (.Y(_01728_),
    .A(net2848),
    .B(net2039));
 sg13g2_o21ai_1 _05866_ (.B1(_01728_),
    .Y(_00730_),
    .A1(net2507),
    .A2(net2039));
 sg13g2_nand2_1 _05867_ (.Y(_01729_),
    .A(net3276),
    .B(net2040));
 sg13g2_o21ai_1 _05868_ (.B1(_01729_),
    .Y(_00731_),
    .A1(net2504),
    .A2(net2040));
 sg13g2_nand2_1 _05869_ (.Y(_01730_),
    .A(net3168),
    .B(net2040));
 sg13g2_o21ai_1 _05870_ (.B1(_01730_),
    .Y(_00732_),
    .A1(net2498),
    .A2(net2040));
 sg13g2_nand2_1 _05871_ (.Y(_01731_),
    .A(net1641),
    .B(net2042));
 sg13g2_o21ai_1 _05872_ (.B1(_01731_),
    .Y(_00733_),
    .A1(net2494),
    .A2(net2042));
 sg13g2_nand2_1 _05873_ (.Y(_01732_),
    .A(net3136),
    .B(net2035));
 sg13g2_o21ai_1 _05874_ (.B1(_01732_),
    .Y(_00734_),
    .A1(net2487),
    .A2(net2035));
 sg13g2_nand2_1 _05875_ (.Y(_01733_),
    .A(net2706),
    .B(net2039));
 sg13g2_o21ai_1 _05876_ (.B1(_01733_),
    .Y(_00735_),
    .A1(net2484),
    .A2(net2039));
 sg13g2_nand2_1 _05877_ (.Y(_01734_),
    .A(net3134),
    .B(net2041));
 sg13g2_o21ai_1 _05878_ (.B1(_01734_),
    .Y(_00736_),
    .A1(net2478),
    .A2(net2041));
 sg13g2_nand2_1 _05879_ (.Y(_01735_),
    .A(net3236),
    .B(net2039));
 sg13g2_o21ai_1 _05880_ (.B1(_01735_),
    .Y(_00737_),
    .A1(net2470),
    .A2(net2039));
 sg13g2_nand2_1 _05881_ (.Y(_01736_),
    .A(net1489),
    .B(net2039));
 sg13g2_o21ai_1 _05882_ (.B1(_01736_),
    .Y(_00738_),
    .A1(net2465),
    .A2(net2039));
 sg13g2_nand2_1 _05883_ (.Y(_01737_),
    .A(net3062),
    .B(net2035));
 sg13g2_o21ai_1 _05884_ (.B1(_01737_),
    .Y(_00739_),
    .A1(net2462),
    .A2(net2035));
 sg13g2_nand2_1 _05885_ (.Y(_01738_),
    .A(net1592),
    .B(net2035));
 sg13g2_o21ai_1 _05886_ (.B1(_01738_),
    .Y(_00740_),
    .A1(net2455),
    .A2(net2035));
 sg13g2_nand2_1 _05887_ (.Y(_01739_),
    .A(net3167),
    .B(net2037));
 sg13g2_o21ai_1 _05888_ (.B1(_01739_),
    .Y(_00741_),
    .A1(net2450),
    .A2(net2037));
 sg13g2_nand2_1 _05889_ (.Y(_01740_),
    .A(net2886),
    .B(net2043));
 sg13g2_o21ai_1 _05890_ (.B1(_01740_),
    .Y(_00742_),
    .A1(net2446),
    .A2(net2043));
 sg13g2_nand2_1 _05891_ (.Y(_01741_),
    .A(net1743),
    .B(net2037));
 sg13g2_o21ai_1 _05892_ (.B1(_01741_),
    .Y(_00743_),
    .A1(net2439),
    .A2(net2037));
 sg13g2_nand2_1 _05893_ (.Y(_01742_),
    .A(net1548),
    .B(net2043));
 sg13g2_o21ai_1 _05894_ (.B1(_01742_),
    .Y(_00744_),
    .A1(net2434),
    .A2(net2043));
 sg13g2_nand2_1 _05895_ (.Y(_01743_),
    .A(net3208),
    .B(net2036));
 sg13g2_o21ai_1 _05896_ (.B1(_01743_),
    .Y(_00745_),
    .A1(net2428),
    .A2(net2036));
 sg13g2_nand2_1 _05897_ (.Y(_01744_),
    .A(net1599),
    .B(net2036));
 sg13g2_o21ai_1 _05898_ (.B1(_01744_),
    .Y(_00746_),
    .A1(net2423),
    .A2(net2036));
 sg13g2_nand2_1 _05899_ (.Y(_01745_),
    .A(net3214),
    .B(net2036));
 sg13g2_o21ai_1 _05900_ (.B1(_01745_),
    .Y(_00747_),
    .A1(net2418),
    .A2(net2036));
 sg13g2_nand2_1 _05901_ (.Y(_01746_),
    .A(net1523),
    .B(net2036));
 sg13g2_o21ai_1 _05902_ (.B1(_01746_),
    .Y(_00748_),
    .A1(net2413),
    .A2(net2036));
 sg13g2_nand2_1 _05903_ (.Y(_01747_),
    .A(net3288),
    .B(net2034));
 sg13g2_o21ai_1 _05904_ (.B1(_01747_),
    .Y(_00749_),
    .A1(net2409),
    .A2(net2034));
 sg13g2_nand2_1 _05905_ (.Y(_01748_),
    .A(net2702),
    .B(net2034));
 sg13g2_o21ai_1 _05906_ (.B1(_01748_),
    .Y(_00750_),
    .A1(net2403),
    .A2(net2034));
 sg13g2_nand2_1 _05907_ (.Y(_01749_),
    .A(net1509),
    .B(net2034));
 sg13g2_o21ai_1 _05908_ (.B1(_01749_),
    .Y(_00751_),
    .A1(net2397),
    .A2(net2034));
 sg13g2_nor2b_1 _05909_ (.A(_01545_),
    .B_N(_01542_),
    .Y(_01750_));
 sg13g2_nor2b_2 _05910_ (.A(_01527_),
    .B_N(net2142),
    .Y(_01751_));
 sg13g2_nand2_2 _05911_ (.Y(_01752_),
    .A(_01678_),
    .B(_01751_));
 sg13g2_nand2_1 _05912_ (.Y(_01753_),
    .A(net2898),
    .B(net2024));
 sg13g2_o21ai_1 _05913_ (.B1(_01753_),
    .Y(_00752_),
    .A1(net2564),
    .A2(net2024));
 sg13g2_nand2_1 _05914_ (.Y(_01754_),
    .A(net1461),
    .B(net2026));
 sg13g2_o21ai_1 _05915_ (.B1(_01754_),
    .Y(_00753_),
    .A1(net2557),
    .A2(net2026));
 sg13g2_nand2_1 _05916_ (.Y(_01755_),
    .A(net2749),
    .B(net2031));
 sg13g2_o21ai_1 _05917_ (.B1(_01755_),
    .Y(_00754_),
    .A1(net2553),
    .A2(net2032));
 sg13g2_nand2_1 _05918_ (.Y(_01756_),
    .A(net1644),
    .B(net2032));
 sg13g2_o21ai_1 _05919_ (.B1(_01756_),
    .Y(_00755_),
    .A1(net2546),
    .A2(net2032));
 sg13g2_nand2_1 _05920_ (.Y(_01757_),
    .A(net2627),
    .B(net2031));
 sg13g2_o21ai_1 _05921_ (.B1(_01757_),
    .Y(_00756_),
    .A1(net2539),
    .A2(net2032));
 sg13g2_nand2_1 _05922_ (.Y(_01758_),
    .A(net1658),
    .B(net2032));
 sg13g2_o21ai_1 _05923_ (.B1(_01758_),
    .Y(_00757_),
    .A1(net2535),
    .A2(net2032));
 sg13g2_nand2_1 _05924_ (.Y(_01759_),
    .A(net2696),
    .B(net2033));
 sg13g2_o21ai_1 _05925_ (.B1(_01759_),
    .Y(_00758_),
    .A1(net2532),
    .A2(net2033));
 sg13g2_nand2_1 _05926_ (.Y(_01760_),
    .A(net3274),
    .B(net2032));
 sg13g2_o21ai_1 _05927_ (.B1(_01760_),
    .Y(_00759_),
    .A1(net2526),
    .A2(net2033));
 sg13g2_nand2_1 _05928_ (.Y(_01761_),
    .A(net2955),
    .B(net2030));
 sg13g2_o21ai_1 _05929_ (.B1(_01761_),
    .Y(_00760_),
    .A1(net2522),
    .A2(net2030));
 sg13g2_nand2_1 _05930_ (.Y(_01762_),
    .A(net1422),
    .B(net2030));
 sg13g2_o21ai_1 _05931_ (.B1(_01762_),
    .Y(_00761_),
    .A1(net2515),
    .A2(net2030));
 sg13g2_nand2_1 _05932_ (.Y(_01763_),
    .A(net2714),
    .B(net2029));
 sg13g2_o21ai_1 _05933_ (.B1(_01763_),
    .Y(_00762_),
    .A1(net2510),
    .A2(net2029));
 sg13g2_nand2_1 _05934_ (.Y(_01764_),
    .A(net1645),
    .B(net2029));
 sg13g2_o21ai_1 _05935_ (.B1(_01764_),
    .Y(_00763_),
    .A1(net2505),
    .A2(net2029));
 sg13g2_nand2_1 _05936_ (.Y(_01765_),
    .A(net2833),
    .B(net2030));
 sg13g2_o21ai_1 _05937_ (.B1(_01765_),
    .Y(_00764_),
    .A1(net2500),
    .A2(net2030));
 sg13g2_nand2_1 _05938_ (.Y(_01766_),
    .A(net1650),
    .B(net2031));
 sg13g2_o21ai_1 _05939_ (.B1(_01766_),
    .Y(_00765_),
    .A1(net2494),
    .A2(net2031));
 sg13g2_nand2_1 _05940_ (.Y(_01767_),
    .A(net1747),
    .B(net2028));
 sg13g2_o21ai_1 _05941_ (.B1(_01767_),
    .Y(_00766_),
    .A1(net2487),
    .A2(net2028));
 sg13g2_nand2_1 _05942_ (.Y(_01768_),
    .A(net1588),
    .B(net2025));
 sg13g2_o21ai_1 _05943_ (.B1(_01768_),
    .Y(_00767_),
    .A1(net2481),
    .A2(net2025));
 sg13g2_nand2_1 _05944_ (.Y(_01769_),
    .A(net2814),
    .B(net2029));
 sg13g2_o21ai_1 _05945_ (.B1(_01769_),
    .Y(_00768_),
    .A1(net2475),
    .A2(net2029));
 sg13g2_nand2_1 _05946_ (.Y(_01770_),
    .A(net3179),
    .B(net2025));
 sg13g2_o21ai_1 _05947_ (.B1(_01770_),
    .Y(_00769_),
    .A1(net2473),
    .A2(net2025));
 sg13g2_nand2_1 _05948_ (.Y(_01771_),
    .A(net1745),
    .B(net2029));
 sg13g2_o21ai_1 _05949_ (.B1(_01771_),
    .Y(_00770_),
    .A1(net2467),
    .A2(net2029));
 sg13g2_nand2_1 _05950_ (.Y(_01772_),
    .A(net1471),
    .B(net2023));
 sg13g2_o21ai_1 _05951_ (.B1(_01772_),
    .Y(_00771_),
    .A1(net2461),
    .A2(net2023));
 sg13g2_nand2_1 _05952_ (.Y(_01773_),
    .A(net1554),
    .B(net2025));
 sg13g2_o21ai_1 _05953_ (.B1(_01773_),
    .Y(_00772_),
    .A1(net2455),
    .A2(net2025));
 sg13g2_nand2_1 _05954_ (.Y(_01774_),
    .A(net2633),
    .B(net2027));
 sg13g2_o21ai_1 _05955_ (.B1(_01774_),
    .Y(_00773_),
    .A1(net2453),
    .A2(net2027));
 sg13g2_nand2_1 _05956_ (.Y(_01775_),
    .A(net1476),
    .B(net2031));
 sg13g2_o21ai_1 _05957_ (.B1(_01775_),
    .Y(_00774_),
    .A1(net2448),
    .A2(net2031));
 sg13g2_nand2_1 _05958_ (.Y(_01776_),
    .A(net3247),
    .B(net2024));
 sg13g2_o21ai_1 _05959_ (.B1(_01776_),
    .Y(_00775_),
    .A1(net2441),
    .A2(net2024));
 sg13g2_nand2_1 _05960_ (.Y(_01777_),
    .A(net1722),
    .B(net2031));
 sg13g2_o21ai_1 _05961_ (.B1(_01777_),
    .Y(_00776_),
    .A1(net2436),
    .A2(net2031));
 sg13g2_nand2_1 _05962_ (.Y(_01778_),
    .A(net2872),
    .B(net2027));
 sg13g2_o21ai_1 _05963_ (.B1(_01778_),
    .Y(_00777_),
    .A1(net2431),
    .A2(net2027));
 sg13g2_nand2_1 _05964_ (.Y(_01779_),
    .A(net3086),
    .B(net2026));
 sg13g2_o21ai_1 _05965_ (.B1(_01779_),
    .Y(_00778_),
    .A1(net2427),
    .A2(net2026));
 sg13g2_nand2_1 _05966_ (.Y(_01780_),
    .A(net2731),
    .B(net2026));
 sg13g2_o21ai_1 _05967_ (.B1(_01780_),
    .Y(_00779_),
    .A1(net2420),
    .A2(net2026));
 sg13g2_nand2_1 _05968_ (.Y(_01781_),
    .A(net1521),
    .B(net2026));
 sg13g2_o21ai_1 _05969_ (.B1(_01781_),
    .Y(_00780_),
    .A1(net2417),
    .A2(net2026));
 sg13g2_nand2_1 _05970_ (.Y(_01782_),
    .A(net1581),
    .B(net2023));
 sg13g2_o21ai_1 _05971_ (.B1(_01782_),
    .Y(_00781_),
    .A1(net2409),
    .A2(net2023));
 sg13g2_nand2_1 _05972_ (.Y(_01783_),
    .A(net2882),
    .B(net2023));
 sg13g2_o21ai_1 _05973_ (.B1(_01783_),
    .Y(_00782_),
    .A1(net2405),
    .A2(net2023));
 sg13g2_nand2_1 _05974_ (.Y(_01784_),
    .A(net2639),
    .B(net2023));
 sg13g2_o21ai_1 _05975_ (.B1(_01784_),
    .Y(_00783_),
    .A1(net2398),
    .A2(net2023));
 sg13g2_and2_1 _05976_ (.A(_01652_),
    .B(net2395),
    .X(_01785_));
 sg13g2_nand2_2 _05977_ (.Y(_01786_),
    .A(net2576),
    .B(_01785_));
 sg13g2_o21ai_1 _05978_ (.B1(net2602),
    .Y(_01787_),
    .A1(net3612),
    .A2(_01786_));
 sg13g2_a21oi_1 _05979_ (.A1(_01339_),
    .A2(_01786_),
    .Y(_00784_),
    .B1(_01787_));
 sg13g2_o21ai_1 _05980_ (.B1(net2602),
    .Y(_01788_),
    .A1(net3652),
    .A2(_01786_));
 sg13g2_a21oi_1 _05981_ (.A1(_01338_),
    .A2(_01786_),
    .Y(_00785_),
    .B1(_01788_));
 sg13g2_o21ai_1 _05982_ (.B1(net1),
    .Y(_01789_),
    .A1(net3576),
    .A2(_01786_));
 sg13g2_a21oi_1 _05983_ (.A1(_01337_),
    .A2(_01786_),
    .Y(_00786_),
    .B1(_01789_));
 sg13g2_o21ai_1 _05984_ (.B1(net2599),
    .Y(_01790_),
    .A1(net3621),
    .A2(_01786_));
 sg13g2_a21oi_1 _05985_ (.A1(_01336_),
    .A2(_01786_),
    .Y(_00787_),
    .B1(_01790_));
 sg13g2_nand2_1 _05986_ (.Y(_01791_),
    .A(_01547_),
    .B(_01613_));
 sg13g2_nand2_1 _05987_ (.Y(_01792_),
    .A(net2913),
    .B(net2088));
 sg13g2_o21ai_1 _05988_ (.B1(_01792_),
    .Y(_00788_),
    .A1(net2562),
    .A2(net2088));
 sg13g2_nand2_1 _05989_ (.Y(_01793_),
    .A(net3163),
    .B(net2090));
 sg13g2_o21ai_1 _05990_ (.B1(_01793_),
    .Y(_00789_),
    .A1(net2555),
    .A2(net2090));
 sg13g2_nand2_1 _05991_ (.Y(_01794_),
    .A(net2651),
    .B(net2094));
 sg13g2_o21ai_1 _05992_ (.B1(_01794_),
    .Y(_00790_),
    .A1(net2550),
    .A2(net2094));
 sg13g2_nand2_1 _05993_ (.Y(_01795_),
    .A(net2893),
    .B(net2093));
 sg13g2_o21ai_1 _05994_ (.B1(_01795_),
    .Y(_00791_),
    .A1(net2545),
    .A2(net2093));
 sg13g2_nand2_1 _05995_ (.Y(_01796_),
    .A(net2672),
    .B(net2093));
 sg13g2_o21ai_1 _05996_ (.B1(_01796_),
    .Y(_00792_),
    .A1(net2541),
    .A2(net2093));
 sg13g2_nand2_1 _05997_ (.Y(_01797_),
    .A(net2781),
    .B(net2093));
 sg13g2_o21ai_1 _05998_ (.B1(_01797_),
    .Y(_00793_),
    .A1(net2537),
    .A2(net2093));
 sg13g2_nand2_1 _05999_ (.Y(_01798_),
    .A(net1513),
    .B(net2095));
 sg13g2_o21ai_1 _06000_ (.B1(_01798_),
    .Y(_00794_),
    .A1(net2531),
    .A2(net2095));
 sg13g2_nand2_1 _06001_ (.Y(_01799_),
    .A(net2982),
    .B(net2093));
 sg13g2_o21ai_1 _06002_ (.B1(_01799_),
    .Y(_00795_),
    .A1(net2524),
    .A2(net2093));
 sg13g2_nand2_1 _06003_ (.Y(_01800_),
    .A(net3073),
    .B(net2092));
 sg13g2_o21ai_1 _06004_ (.B1(_01800_),
    .Y(_00796_),
    .A1(net2520),
    .A2(net2092));
 sg13g2_nand2_1 _06005_ (.Y(_01801_),
    .A(net1702),
    .B(net2092));
 sg13g2_o21ai_1 _06006_ (.B1(_01801_),
    .Y(_00797_),
    .A1(net2516),
    .A2(net2092));
 sg13g2_nand2_1 _06007_ (.Y(_01802_),
    .A(net1716),
    .B(net2092));
 sg13g2_o21ai_1 _06008_ (.B1(_01802_),
    .Y(_00798_),
    .A1(net2508),
    .A2(net2092));
 sg13g2_nand2_1 _06009_ (.Y(_01803_),
    .A(net2858),
    .B(net2091));
 sg13g2_o21ai_1 _06010_ (.B1(_01803_),
    .Y(_00799_),
    .A1(net2503),
    .A2(net2091));
 sg13g2_nand2_1 _06011_ (.Y(_01804_),
    .A(net3377),
    .B(net2092));
 sg13g2_o21ai_1 _06012_ (.B1(_01804_),
    .Y(_00800_),
    .A1(net2497),
    .A2(net2092));
 sg13g2_nand2_1 _06013_ (.Y(_01805_),
    .A(net3018),
    .B(net2091));
 sg13g2_o21ai_1 _06014_ (.B1(_01805_),
    .Y(_00801_),
    .A1(net2491),
    .A2(net2091));
 sg13g2_nand2_1 _06015_ (.Y(_01806_),
    .A(net1578),
    .B(net2088));
 sg13g2_o21ai_1 _06016_ (.B1(_01806_),
    .Y(_00802_),
    .A1(net2488),
    .A2(net2096));
 sg13g2_nand2_1 _06017_ (.Y(_01807_),
    .A(net1445),
    .B(net2091));
 sg13g2_o21ai_1 _06018_ (.B1(_01807_),
    .Y(_00803_),
    .A1(net2484),
    .A2(net2091));
 sg13g2_nand2_1 _06019_ (.Y(_01808_),
    .A(net2799),
    .B(net2094));
 sg13g2_o21ai_1 _06020_ (.B1(_01808_),
    .Y(_00804_),
    .A1(net2480),
    .A2(net2094));
 sg13g2_nand2_1 _06021_ (.Y(_01809_),
    .A(net1605),
    .B(net2088));
 sg13g2_o21ai_1 _06022_ (.B1(_01809_),
    .Y(_00805_),
    .A1(net2470),
    .A2(net2088));
 sg13g2_nand2_1 _06023_ (.Y(_01810_),
    .A(net2608),
    .B(net2091));
 sg13g2_o21ai_1 _06024_ (.B1(_01810_),
    .Y(_00806_),
    .A1(net2467),
    .A2(net2091));
 sg13g2_nand2_1 _06025_ (.Y(_01811_),
    .A(net2626),
    .B(net2087));
 sg13g2_o21ai_1 _06026_ (.B1(_01811_),
    .Y(_00807_),
    .A1(net2461),
    .A2(net2087));
 sg13g2_nand2_1 _06027_ (.Y(_01812_),
    .A(net2609),
    .B(net2088));
 sg13g2_o21ai_1 _06028_ (.B1(_01812_),
    .Y(_00808_),
    .A1(net2459),
    .A2(net2088));
 sg13g2_nand2_1 _06029_ (.Y(_01813_),
    .A(net2623),
    .B(net2090));
 sg13g2_o21ai_1 _06030_ (.B1(_01813_),
    .Y(_00809_),
    .A1(net2450),
    .A2(net2090));
 sg13g2_nand2_1 _06031_ (.Y(_01814_),
    .A(net1629),
    .B(net2094));
 sg13g2_o21ai_1 _06032_ (.B1(_01814_),
    .Y(_00810_),
    .A1(net2447),
    .A2(net2094));
 sg13g2_nand2_1 _06033_ (.Y(_01815_),
    .A(net1669),
    .B(net2089));
 sg13g2_o21ai_1 _06034_ (.B1(_01815_),
    .Y(_00811_),
    .A1(net2440),
    .A2(net2089));
 sg13g2_nand2_1 _06035_ (.Y(_01816_),
    .A(net1695),
    .B(net2094));
 sg13g2_o21ai_1 _06036_ (.B1(_01816_),
    .Y(_00812_),
    .A1(net2434),
    .A2(net2094));
 sg13g2_nand2_1 _06037_ (.Y(_01817_),
    .A(net2669),
    .B(net2089));
 sg13g2_o21ai_1 _06038_ (.B1(_01817_),
    .Y(_00813_),
    .A1(net2428),
    .A2(net2089));
 sg13g2_nand2_1 _06039_ (.Y(_01818_),
    .A(net3020),
    .B(net2090));
 sg13g2_o21ai_1 _06040_ (.B1(_01818_),
    .Y(_00814_),
    .A1(net2423),
    .A2(net2089));
 sg13g2_nand2_1 _06041_ (.Y(_01819_),
    .A(net3014),
    .B(net2089));
 sg13g2_o21ai_1 _06042_ (.B1(_01819_),
    .Y(_00815_),
    .A1(net2418),
    .A2(net2090));
 sg13g2_nand2_1 _06043_ (.Y(_01820_),
    .A(net2842),
    .B(net2089));
 sg13g2_o21ai_1 _06044_ (.B1(_01820_),
    .Y(_00816_),
    .A1(net2415),
    .A2(net2089));
 sg13g2_nand2_1 _06045_ (.Y(_01821_),
    .A(net2709),
    .B(net2087));
 sg13g2_o21ai_1 _06046_ (.B1(_01821_),
    .Y(_00817_),
    .A1(net2412),
    .A2(net2087));
 sg13g2_nand2_1 _06047_ (.Y(_01822_),
    .A(net3004),
    .B(net2087));
 sg13g2_o21ai_1 _06048_ (.B1(_01822_),
    .Y(_00818_),
    .A1(net2402),
    .A2(net2087));
 sg13g2_nand2_1 _06049_ (.Y(_01823_),
    .A(net3253),
    .B(net2087));
 sg13g2_o21ai_1 _06050_ (.B1(_01823_),
    .Y(_00819_),
    .A1(net2400),
    .A2(net2087));
 sg13g2_or2_1 _06051_ (.X(_01824_),
    .B(_01538_),
    .A(_01535_));
 sg13g2_nor2_2 _06052_ (.A(net2325),
    .B(_01824_),
    .Y(_01825_));
 sg13g2_or2_1 _06053_ (.X(_01826_),
    .B(_01824_),
    .A(net2325));
 sg13g2_nand2_1 _06054_ (.Y(_01827_),
    .A(_01751_),
    .B(_01825_));
 sg13g2_nand2_1 _06055_ (.Y(_01828_),
    .A(net1707),
    .B(net2012));
 sg13g2_o21ai_1 _06056_ (.B1(_01828_),
    .Y(_00820_),
    .A1(net2561),
    .A2(net2012));
 sg13g2_nand2_1 _06057_ (.Y(_01829_),
    .A(net1542),
    .B(net2015));
 sg13g2_o21ai_1 _06058_ (.B1(_01829_),
    .Y(_00821_),
    .A1(net2557),
    .A2(net2015));
 sg13g2_nand2_1 _06059_ (.Y(_01830_),
    .A(net2700),
    .B(net2020));
 sg13g2_o21ai_1 _06060_ (.B1(_01830_),
    .Y(_00822_),
    .A1(net2552),
    .A2(net2020));
 sg13g2_nand2_1 _06061_ (.Y(_01831_),
    .A(net1686),
    .B(net2021));
 sg13g2_o21ai_1 _06062_ (.B1(_01831_),
    .Y(_00823_),
    .A1(net2548),
    .A2(net2021));
 sg13g2_nand2_1 _06063_ (.Y(_01832_),
    .A(net1494),
    .B(net2020));
 sg13g2_o21ai_1 _06064_ (.B1(_01832_),
    .Y(_00824_),
    .A1(net2543),
    .A2(net2020));
 sg13g2_nand2_1 _06065_ (.Y(_01833_),
    .A(net3329),
    .B(net2021));
 sg13g2_o21ai_1 _06066_ (.B1(_01833_),
    .Y(_00825_),
    .A1(net2534),
    .A2(net2021));
 sg13g2_nand2_1 _06067_ (.Y(_01834_),
    .A(net2693),
    .B(net2021));
 sg13g2_o21ai_1 _06068_ (.B1(_01834_),
    .Y(_00826_),
    .A1(net2528),
    .A2(net2021));
 sg13g2_nand2_1 _06069_ (.Y(_01835_),
    .A(net1621),
    .B(net2018));
 sg13g2_o21ai_1 _06070_ (.B1(_01835_),
    .Y(_00827_),
    .A1(net2525),
    .A2(net2018));
 sg13g2_nand2_1 _06071_ (.Y(_01836_),
    .A(net3061),
    .B(net2018));
 sg13g2_o21ai_1 _06072_ (.B1(_01836_),
    .Y(_00828_),
    .A1(net2519),
    .A2(net2018));
 sg13g2_nand2_1 _06073_ (.Y(_01837_),
    .A(net2960),
    .B(net2017));
 sg13g2_o21ai_1 _06074_ (.B1(_01837_),
    .Y(_00829_),
    .A1(net2512),
    .A2(net2017));
 sg13g2_nand2_1 _06075_ (.Y(_01838_),
    .A(net2973),
    .B(net2017));
 sg13g2_o21ai_1 _06076_ (.B1(_01838_),
    .Y(_00830_),
    .A1(net2508),
    .A2(net2017));
 sg13g2_nand2_1 _06077_ (.Y(_01839_),
    .A(net3267),
    .B(net2017));
 sg13g2_o21ai_1 _06078_ (.B1(_01839_),
    .Y(_00831_),
    .A1(net2504),
    .A2(net2017));
 sg13g2_nand2_1 _06079_ (.Y(_01840_),
    .A(net1528),
    .B(net2017));
 sg13g2_o21ai_1 _06080_ (.B1(_01840_),
    .Y(_00832_),
    .A1(net2499),
    .A2(net2017));
 sg13g2_nand2_1 _06081_ (.Y(_01841_),
    .A(net1703),
    .B(net2018));
 sg13g2_o21ai_1 _06082_ (.B1(_01841_),
    .Y(_00833_),
    .A1(net2493),
    .A2(net2018));
 sg13g2_nand2_1 _06083_ (.Y(_01842_),
    .A(net1426),
    .B(net2013));
 sg13g2_o21ai_1 _06084_ (.B1(_01842_),
    .Y(_00834_),
    .A1(net2487),
    .A2(net2013));
 sg13g2_nand2_1 _06085_ (.Y(_01843_),
    .A(net2737),
    .B(net2019));
 sg13g2_o21ai_1 _06086_ (.B1(_01843_),
    .Y(_00835_),
    .A1(net2481),
    .A2(net2019));
 sg13g2_nand2_1 _06087_ (.Y(_01844_),
    .A(net3050),
    .B(net2019));
 sg13g2_o21ai_1 _06088_ (.B1(_01844_),
    .Y(_00836_),
    .A1(net2476),
    .A2(net2019));
 sg13g2_nand2_1 _06089_ (.Y(_01845_),
    .A(net2726),
    .B(net2013));
 sg13g2_o21ai_1 _06090_ (.B1(_01845_),
    .Y(_00837_),
    .A1(net2473),
    .A2(net2013));
 sg13g2_nand2_1 _06091_ (.Y(_01846_),
    .A(net1500),
    .B(net2019));
 sg13g2_o21ai_1 _06092_ (.B1(_01846_),
    .Y(_00838_),
    .A1(net2465),
    .A2(net2019));
 sg13g2_nand2_1 _06093_ (.Y(_01847_),
    .A(net3000),
    .B(net2013));
 sg13g2_o21ai_1 _06094_ (.B1(_01847_),
    .Y(_00839_),
    .A1(net2463),
    .A2(net2013));
 sg13g2_nand2_1 _06095_ (.Y(_01848_),
    .A(net1663),
    .B(net2013));
 sg13g2_o21ai_1 _06096_ (.B1(_01848_),
    .Y(_00840_),
    .A1(net2458),
    .A2(net2013));
 sg13g2_nand2_1 _06097_ (.Y(_01849_),
    .A(net1568),
    .B(net2015));
 sg13g2_o21ai_1 _06098_ (.B1(_01849_),
    .Y(_00841_),
    .A1(net2454),
    .A2(net2015));
 sg13g2_nand2_1 _06099_ (.Y(_01850_),
    .A(net1643),
    .B(net2020));
 sg13g2_o21ai_1 _06100_ (.B1(_01850_),
    .Y(_00842_),
    .A1(net2446),
    .A2(net2020));
 sg13g2_nand2_1 _06101_ (.Y(_01851_),
    .A(net2912),
    .B(net2014));
 sg13g2_o21ai_1 _06102_ (.B1(_01851_),
    .Y(_00843_),
    .A1(net2441),
    .A2(net2014));
 sg13g2_nand2_1 _06103_ (.Y(_01852_),
    .A(net3176),
    .B(net2020));
 sg13g2_o21ai_1 _06104_ (.B1(_01852_),
    .Y(_00844_),
    .A1(net2436),
    .A2(net2020));
 sg13g2_nand2_1 _06105_ (.Y(_01853_),
    .A(net2974),
    .B(net2014));
 sg13g2_o21ai_1 _06106_ (.B1(_01853_),
    .Y(_00845_),
    .A1(net2429),
    .A2(net2014));
 sg13g2_nand2_1 _06107_ (.Y(_01854_),
    .A(net1596),
    .B(net2015));
 sg13g2_o21ai_1 _06108_ (.B1(_01854_),
    .Y(_00846_),
    .A1(net2427),
    .A2(net2015));
 sg13g2_nand2_1 _06109_ (.Y(_01855_),
    .A(net3016),
    .B(net2014));
 sg13g2_o21ai_1 _06110_ (.B1(_01855_),
    .Y(_00847_),
    .A1(net2421),
    .A2(net2014));
 sg13g2_nand2_1 _06111_ (.Y(_01856_),
    .A(net1628),
    .B(net2014));
 sg13g2_o21ai_1 _06112_ (.B1(_01856_),
    .Y(_00848_),
    .A1(net2414),
    .A2(net2014));
 sg13g2_nand2_1 _06113_ (.Y(_01857_),
    .A(net1632),
    .B(net2012));
 sg13g2_o21ai_1 _06114_ (.B1(_01857_),
    .Y(_00849_),
    .A1(net2408),
    .A2(net2012));
 sg13g2_nand2_1 _06115_ (.Y(_01858_),
    .A(net1507),
    .B(net2012));
 sg13g2_o21ai_1 _06116_ (.B1(_01858_),
    .Y(_00850_),
    .A1(net2405),
    .A2(net2012));
 sg13g2_nand2_1 _06117_ (.Y(_01859_),
    .A(net2698),
    .B(net2012));
 sg13g2_o21ai_1 _06118_ (.B1(_01859_),
    .Y(_00851_),
    .A1(net2398),
    .A2(net2012));
 sg13g2_nand2_1 _06119_ (.Y(_01860_),
    .A(_01613_),
    .B(_01751_));
 sg13g2_nand2_1 _06120_ (.Y(_01861_),
    .A(net2824),
    .B(net2002));
 sg13g2_o21ai_1 _06121_ (.B1(_01861_),
    .Y(_00852_),
    .A1(net2562),
    .A2(net2002));
 sg13g2_nand2_1 _06122_ (.Y(_01862_),
    .A(net3064),
    .B(net2005));
 sg13g2_o21ai_1 _06123_ (.B1(_01862_),
    .Y(_00853_),
    .A1(net2555),
    .A2(net2005));
 sg13g2_nand2_1 _06124_ (.Y(_01863_),
    .A(net3055),
    .B(net2009));
 sg13g2_o21ai_1 _06125_ (.B1(_01863_),
    .Y(_00854_),
    .A1(net2550),
    .A2(net2009));
 sg13g2_nand2_1 _06126_ (.Y(_01864_),
    .A(net2808),
    .B(net2008));
 sg13g2_o21ai_1 _06127_ (.B1(_01864_),
    .Y(_00855_),
    .A1(net2545),
    .A2(net2008));
 sg13g2_nand2_1 _06128_ (.Y(_01865_),
    .A(net2613),
    .B(net2008));
 sg13g2_o21ai_1 _06129_ (.B1(_01865_),
    .Y(_00856_),
    .A1(net2541),
    .A2(net2008));
 sg13g2_nand2_1 _06130_ (.Y(_01866_),
    .A(net2877),
    .B(net2008));
 sg13g2_o21ai_1 _06131_ (.B1(_01866_),
    .Y(_00857_),
    .A1(net2533),
    .A2(net2008));
 sg13g2_nand2_1 _06132_ (.Y(_01867_),
    .A(net2762),
    .B(net2010));
 sg13g2_o21ai_1 _06133_ (.B1(_01867_),
    .Y(_00858_),
    .A1(net2531),
    .A2(net2010));
 sg13g2_nand2_1 _06134_ (.Y(_01868_),
    .A(net3132),
    .B(net2008));
 sg13g2_o21ai_1 _06135_ (.B1(_01868_),
    .Y(_00859_),
    .A1(net2524),
    .A2(net2008));
 sg13g2_nand2_1 _06136_ (.Y(_01869_),
    .A(net2846),
    .B(net2007));
 sg13g2_o21ai_1 _06137_ (.B1(_01869_),
    .Y(_00860_),
    .A1(net2519),
    .A2(net2007));
 sg13g2_nand2_1 _06138_ (.Y(_01870_),
    .A(net2603),
    .B(net2007));
 sg13g2_o21ai_1 _06139_ (.B1(_01870_),
    .Y(_00861_),
    .A1(net2516),
    .A2(net2007));
 sg13g2_nand2_1 _06140_ (.Y(_01871_),
    .A(net2701),
    .B(net2007));
 sg13g2_o21ai_1 _06141_ (.B1(_01871_),
    .Y(_00862_),
    .A1(net2508),
    .A2(net2007));
 sg13g2_nand2_1 _06142_ (.Y(_01872_),
    .A(net2647),
    .B(net2006));
 sg13g2_o21ai_1 _06143_ (.B1(_01872_),
    .Y(_00863_),
    .A1(net2503),
    .A2(net2006));
 sg13g2_nand2_1 _06144_ (.Y(_01873_),
    .A(net3186),
    .B(net2007));
 sg13g2_o21ai_1 _06145_ (.B1(_01873_),
    .Y(_00864_),
    .A1(net2497),
    .A2(net2007));
 sg13g2_nand2_1 _06146_ (.Y(_01874_),
    .A(net1642),
    .B(net2006));
 sg13g2_o21ai_1 _06147_ (.B1(_01874_),
    .Y(_00865_),
    .A1(net2491),
    .A2(net2006));
 sg13g2_nand2_1 _06148_ (.Y(_01875_),
    .A(net1423),
    .B(net2003));
 sg13g2_o21ai_1 _06149_ (.B1(_01875_),
    .Y(_00866_),
    .A1(net2488),
    .A2(net2003));
 sg13g2_nand2_1 _06150_ (.Y(_01876_),
    .A(net1618),
    .B(net2006));
 sg13g2_o21ai_1 _06151_ (.B1(_01876_),
    .Y(_00867_),
    .A1(net2483),
    .A2(net2006));
 sg13g2_nand2_1 _06152_ (.Y(_01877_),
    .A(net3162),
    .B(net2009));
 sg13g2_o21ai_1 _06153_ (.B1(_01877_),
    .Y(_00868_),
    .A1(net2480),
    .A2(net2009));
 sg13g2_nand2_1 _06154_ (.Y(_01878_),
    .A(net2694),
    .B(net2003));
 sg13g2_o21ai_1 _06155_ (.B1(_01878_),
    .Y(_00869_),
    .A1(net2470),
    .A2(net2003));
 sg13g2_nand2_1 _06156_ (.Y(_01879_),
    .A(net1512),
    .B(net2006));
 sg13g2_o21ai_1 _06157_ (.B1(_01879_),
    .Y(_00870_),
    .A1(net2467),
    .A2(net2006));
 sg13g2_nand2_1 _06158_ (.Y(_01880_),
    .A(net2728),
    .B(net2001));
 sg13g2_o21ai_1 _06159_ (.B1(_01880_),
    .Y(_00871_),
    .A1(net2461),
    .A2(net2001));
 sg13g2_nand2_1 _06160_ (.Y(_01881_),
    .A(net3001),
    .B(net2003));
 sg13g2_o21ai_1 _06161_ (.B1(_01881_),
    .Y(_00872_),
    .A1(net2458),
    .A2(net2003));
 sg13g2_nand2_1 _06162_ (.Y(_01882_),
    .A(net2774),
    .B(net2005));
 sg13g2_o21ai_1 _06163_ (.B1(_01882_),
    .Y(_00873_),
    .A1(net2450),
    .A2(net2005));
 sg13g2_nand2_1 _06164_ (.Y(_01883_),
    .A(net1604),
    .B(net2009));
 sg13g2_o21ai_1 _06165_ (.B1(_01883_),
    .Y(_00874_),
    .A1(net2447),
    .A2(net2009));
 sg13g2_nand2_1 _06166_ (.Y(_01884_),
    .A(net2736),
    .B(net2002));
 sg13g2_o21ai_1 _06167_ (.B1(_01884_),
    .Y(_00875_),
    .A1(net2440),
    .A2(net2002));
 sg13g2_nand2_1 _06168_ (.Y(_01885_),
    .A(net3227),
    .B(net2009));
 sg13g2_o21ai_1 _06169_ (.B1(_01885_),
    .Y(_00876_),
    .A1(net2435),
    .A2(net2009));
 sg13g2_nand2_1 _06170_ (.Y(_01886_),
    .A(net1679),
    .B(net2004));
 sg13g2_o21ai_1 _06171_ (.B1(_01886_),
    .Y(_00877_),
    .A1(net2428),
    .A2(net2004));
 sg13g2_nand2_1 _06172_ (.Y(_01887_),
    .A(net1725),
    .B(net2004));
 sg13g2_o21ai_1 _06173_ (.B1(_01887_),
    .Y(_00878_),
    .A1(net2423),
    .A2(net2004));
 sg13g2_nand2_1 _06174_ (.Y(_01888_),
    .A(net2754),
    .B(net2004));
 sg13g2_o21ai_1 _06175_ (.B1(_01888_),
    .Y(_00879_),
    .A1(net2419),
    .A2(net2004));
 sg13g2_nand2_1 _06176_ (.Y(_01889_),
    .A(net1673),
    .B(net2004));
 sg13g2_o21ai_1 _06177_ (.B1(_01889_),
    .Y(_00880_),
    .A1(net2415),
    .A2(net2004));
 sg13g2_nand2_1 _06178_ (.Y(_01890_),
    .A(net3034),
    .B(net2001));
 sg13g2_o21ai_1 _06179_ (.B1(_01890_),
    .Y(_00881_),
    .A1(net2412),
    .A2(net2001));
 sg13g2_nand2_1 _06180_ (.Y(_01891_),
    .A(net2753),
    .B(net2001));
 sg13g2_o21ai_1 _06181_ (.B1(_01891_),
    .Y(_00882_),
    .A1(net2404),
    .A2(net2001));
 sg13g2_nand2_1 _06182_ (.Y(_01892_),
    .A(net2673),
    .B(net2001));
 sg13g2_o21ai_1 _06183_ (.B1(_01892_),
    .Y(_00883_),
    .A1(net2400),
    .A2(net2001));
 sg13g2_nand2_1 _06184_ (.Y(_01893_),
    .A(_01716_),
    .B(_01825_));
 sg13g2_nand2_1 _06185_ (.Y(_01894_),
    .A(net1685),
    .B(net1991));
 sg13g2_o21ai_1 _06186_ (.B1(_01894_),
    .Y(_00884_),
    .A1(net2561),
    .A2(net1991));
 sg13g2_nand2_1 _06187_ (.Y(_01895_),
    .A(net2662),
    .B(net1992));
 sg13g2_o21ai_1 _06188_ (.B1(_01895_),
    .Y(_00885_),
    .A1(net2557),
    .A2(net1992));
 sg13g2_nand2_1 _06189_ (.Y(_01896_),
    .A(net3092),
    .B(net1998));
 sg13g2_o21ai_1 _06190_ (.B1(_01896_),
    .Y(_00886_),
    .A1(net2552),
    .A2(net1998));
 sg13g2_nand2_1 _06191_ (.Y(_01897_),
    .A(net3246),
    .B(net1999));
 sg13g2_o21ai_1 _06192_ (.B1(_01897_),
    .Y(_00887_),
    .A1(net2548),
    .A2(net1999));
 sg13g2_nand2_1 _06193_ (.Y(_01898_),
    .A(net2646),
    .B(net1998));
 sg13g2_o21ai_1 _06194_ (.B1(_01898_),
    .Y(_00888_),
    .A1(net2543),
    .A2(net1998));
 sg13g2_nand2_1 _06195_ (.Y(_01899_),
    .A(net3312),
    .B(net1999));
 sg13g2_o21ai_1 _06196_ (.B1(_01899_),
    .Y(_00889_),
    .A1(net2534),
    .A2(net1999));
 sg13g2_nand2_1 _06197_ (.Y(_01900_),
    .A(net1637),
    .B(net1999));
 sg13g2_o21ai_1 _06198_ (.B1(_01900_),
    .Y(_00890_),
    .A1(net2528),
    .A2(net1999));
 sg13g2_nand2_1 _06199_ (.Y(_01901_),
    .A(net1646),
    .B(net1996));
 sg13g2_o21ai_1 _06200_ (.B1(_01901_),
    .Y(_00891_),
    .A1(net2525),
    .A2(net1996));
 sg13g2_nand2_1 _06201_ (.Y(_01902_),
    .A(net1453),
    .B(net1996));
 sg13g2_o21ai_1 _06202_ (.B1(_01902_),
    .Y(_00892_),
    .A1(net2519),
    .A2(net1996));
 sg13g2_nand2_1 _06203_ (.Y(_01903_),
    .A(net1552),
    .B(net1995));
 sg13g2_o21ai_1 _06204_ (.B1(_01903_),
    .Y(_00893_),
    .A1(net2512),
    .A2(net1995));
 sg13g2_nand2_1 _06205_ (.Y(_01904_),
    .A(net2677),
    .B(net1995));
 sg13g2_o21ai_1 _06206_ (.B1(_01904_),
    .Y(_00894_),
    .A1(net2508),
    .A2(net1995));
 sg13g2_nand2_1 _06207_ (.Y(_01905_),
    .A(net2987),
    .B(net1995));
 sg13g2_o21ai_1 _06208_ (.B1(_01905_),
    .Y(_00895_),
    .A1(net2504),
    .A2(net1995));
 sg13g2_nand2_1 _06209_ (.Y(_01906_),
    .A(net1717),
    .B(net1995));
 sg13g2_o21ai_1 _06210_ (.B1(_01906_),
    .Y(_00896_),
    .A1(net2499),
    .A2(net1995));
 sg13g2_nand2_1 _06211_ (.Y(_01907_),
    .A(net3148),
    .B(net1996));
 sg13g2_o21ai_1 _06212_ (.B1(_01907_),
    .Y(_00897_),
    .A1(net2493),
    .A2(net1996));
 sg13g2_nand2_1 _06213_ (.Y(_01908_),
    .A(net3010),
    .B(net1991));
 sg13g2_o21ai_1 _06214_ (.B1(_01908_),
    .Y(_00898_),
    .A1(net2487),
    .A2(net1991));
 sg13g2_nand2_1 _06215_ (.Y(_01909_),
    .A(net2923),
    .B(net1997));
 sg13g2_o21ai_1 _06216_ (.B1(_01909_),
    .Y(_00899_),
    .A1(net2482),
    .A2(net1997));
 sg13g2_nand2_1 _06217_ (.Y(_01910_),
    .A(net2997),
    .B(net1997));
 sg13g2_o21ai_1 _06218_ (.B1(_01910_),
    .Y(_00900_),
    .A1(net2476),
    .A2(net1997));
 sg13g2_nand2_1 _06219_ (.Y(_01911_),
    .A(net2980),
    .B(net1991));
 sg13g2_o21ai_1 _06220_ (.B1(_01911_),
    .Y(_00901_),
    .A1(net2473),
    .A2(net1991));
 sg13g2_nand2_1 _06221_ (.Y(_01912_),
    .A(net2796),
    .B(net1997));
 sg13g2_o21ai_1 _06222_ (.B1(_01912_),
    .Y(_00902_),
    .A1(net2469),
    .A2(net1997));
 sg13g2_nand2_1 _06223_ (.Y(_01913_),
    .A(net2649),
    .B(net1994));
 sg13g2_o21ai_1 _06224_ (.B1(_01913_),
    .Y(_00903_),
    .A1(net2463),
    .A2(net1994));
 sg13g2_nand2_1 _06225_ (.Y(_01914_),
    .A(net3300),
    .B(net1991));
 sg13g2_o21ai_1 _06226_ (.B1(_01914_),
    .Y(_00904_),
    .A1(net2458),
    .A2(net1994));
 sg13g2_nand2_1 _06227_ (.Y(_01915_),
    .A(net3296),
    .B(net1993));
 sg13g2_o21ai_1 _06228_ (.B1(_01915_),
    .Y(_00905_),
    .A1(net2454),
    .A2(net1993));
 sg13g2_nand2_1 _06229_ (.Y(_01916_),
    .A(net2648),
    .B(net1998));
 sg13g2_o21ai_1 _06230_ (.B1(_01916_),
    .Y(_00906_),
    .A1(net2446),
    .A2(net1998));
 sg13g2_nand2_1 _06231_ (.Y(_01917_),
    .A(net3301),
    .B(net1990));
 sg13g2_o21ai_1 _06232_ (.B1(_01917_),
    .Y(_00907_),
    .A1(net2441),
    .A2(net1990));
 sg13g2_nand2_1 _06233_ (.Y(_01918_),
    .A(net3220),
    .B(net1998));
 sg13g2_o21ai_1 _06234_ (.B1(_01918_),
    .Y(_00908_),
    .A1(net2436),
    .A2(net1998));
 sg13g2_nand2_1 _06235_ (.Y(_01919_),
    .A(net3026),
    .B(net1992));
 sg13g2_o21ai_1 _06236_ (.B1(_01919_),
    .Y(_00909_),
    .A1(net2430),
    .A2(net1992));
 sg13g2_nand2_1 _06237_ (.Y(_01920_),
    .A(net1442),
    .B(net1993));
 sg13g2_o21ai_1 _06238_ (.B1(_01920_),
    .Y(_00910_),
    .A1(net2427),
    .A2(net1993));
 sg13g2_nand2_1 _06239_ (.Y(_01921_),
    .A(net3189),
    .B(net1992));
 sg13g2_o21ai_1 _06240_ (.B1(_01921_),
    .Y(_00911_),
    .A1(net2421),
    .A2(net1992));
 sg13g2_nand2_1 _06241_ (.Y(_01922_),
    .A(net3097),
    .B(net1992));
 sg13g2_o21ai_1 _06242_ (.B1(_01922_),
    .Y(_00912_),
    .A1(net2413),
    .A2(net1992));
 sg13g2_nand2_1 _06243_ (.Y(_01923_),
    .A(net2971),
    .B(net1990));
 sg13g2_o21ai_1 _06244_ (.B1(_01923_),
    .Y(_00913_),
    .A1(net2408),
    .A2(net1990));
 sg13g2_nand2_1 _06245_ (.Y(_01924_),
    .A(net1590),
    .B(net1990));
 sg13g2_o21ai_1 _06246_ (.B1(_01924_),
    .Y(_00914_),
    .A1(net2405),
    .A2(net1990));
 sg13g2_nand2_1 _06247_ (.Y(_01925_),
    .A(net1594),
    .B(net1990));
 sg13g2_o21ai_1 _06248_ (.B1(_01925_),
    .Y(_00915_),
    .A1(net2397),
    .A2(net1990));
 sg13g2_nand2_1 _06249_ (.Y(_01926_),
    .A(_01613_),
    .B(_01716_));
 sg13g2_nand2_1 _06250_ (.Y(_01927_),
    .A(net3142),
    .B(net1980));
 sg13g2_o21ai_1 _06251_ (.B1(_01927_),
    .Y(_00916_),
    .A1(net2562),
    .A2(net1980));
 sg13g2_nand2_1 _06252_ (.Y(_01928_),
    .A(net2785),
    .B(net1983));
 sg13g2_o21ai_1 _06253_ (.B1(_01928_),
    .Y(_00917_),
    .A1(net2555),
    .A2(net1983));
 sg13g2_nand2_1 _06254_ (.Y(_01929_),
    .A(net2929),
    .B(net1987));
 sg13g2_o21ai_1 _06255_ (.B1(_01929_),
    .Y(_00918_),
    .A1(net2550),
    .A2(net1987));
 sg13g2_nand2_1 _06256_ (.Y(_01930_),
    .A(net2659),
    .B(net1986));
 sg13g2_o21ai_1 _06257_ (.B1(_01930_),
    .Y(_00919_),
    .A1(net2545),
    .A2(net1986));
 sg13g2_nand2_1 _06258_ (.Y(_01931_),
    .A(net1480),
    .B(net1986));
 sg13g2_o21ai_1 _06259_ (.B1(_01931_),
    .Y(_00920_),
    .A1(net2543),
    .A2(net1986));
 sg13g2_nand2_1 _06260_ (.Y(_01932_),
    .A(net1515),
    .B(net1986));
 sg13g2_o21ai_1 _06261_ (.B1(_01932_),
    .Y(_00921_),
    .A1(net2533),
    .A2(net1986));
 sg13g2_nand2_1 _06262_ (.Y(_01933_),
    .A(net2717),
    .B(net1988));
 sg13g2_o21ai_1 _06263_ (.B1(_01933_),
    .Y(_00922_),
    .A1(net2531),
    .A2(net1988));
 sg13g2_nand2_1 _06264_ (.Y(_01934_),
    .A(net2965),
    .B(net1986));
 sg13g2_o21ai_1 _06265_ (.B1(_01934_),
    .Y(_00923_),
    .A1(net2524),
    .A2(net1986));
 sg13g2_nand2_1 _06266_ (.Y(_01935_),
    .A(net3069),
    .B(net1985));
 sg13g2_o21ai_1 _06267_ (.B1(_01935_),
    .Y(_00924_),
    .A1(net2519),
    .A2(net1985));
 sg13g2_nand2_1 _06268_ (.Y(_01936_),
    .A(net1638),
    .B(net1985));
 sg13g2_o21ai_1 _06269_ (.B1(_01936_),
    .Y(_00925_),
    .A1(net2516),
    .A2(net1985));
 sg13g2_nand2_1 _06270_ (.Y(_01937_),
    .A(net1560),
    .B(net1985));
 sg13g2_o21ai_1 _06271_ (.B1(_01937_),
    .Y(_00926_),
    .A1(net2508),
    .A2(net1985));
 sg13g2_nand2_1 _06272_ (.Y(_01938_),
    .A(net2927),
    .B(net1984));
 sg13g2_o21ai_1 _06273_ (.B1(_01938_),
    .Y(_00927_),
    .A1(net2503),
    .A2(net1984));
 sg13g2_nand2_1 _06274_ (.Y(_01939_),
    .A(net3318),
    .B(net1985));
 sg13g2_o21ai_1 _06275_ (.B1(_01939_),
    .Y(_00928_),
    .A1(net2497),
    .A2(net1985));
 sg13g2_nand2_1 _06276_ (.Y(_01940_),
    .A(net3213),
    .B(net1984));
 sg13g2_o21ai_1 _06277_ (.B1(_01940_),
    .Y(_00929_),
    .A1(net2491),
    .A2(net1984));
 sg13g2_nand2_1 _06278_ (.Y(_01941_),
    .A(net2820),
    .B(net1981));
 sg13g2_o21ai_1 _06279_ (.B1(_01941_),
    .Y(_00930_),
    .A1(net2488),
    .A2(net1981));
 sg13g2_nand2_1 _06280_ (.Y(_01942_),
    .A(net3135),
    .B(net1984));
 sg13g2_o21ai_1 _06281_ (.B1(_01942_),
    .Y(_00931_),
    .A1(net2485),
    .A2(net1984));
 sg13g2_nand2_1 _06282_ (.Y(_01943_),
    .A(net2690),
    .B(net1987));
 sg13g2_o21ai_1 _06283_ (.B1(_01943_),
    .Y(_00932_),
    .A1(net2480),
    .A2(net1987));
 sg13g2_nand2_1 _06284_ (.Y(_01944_),
    .A(net2723),
    .B(net1981));
 sg13g2_o21ai_1 _06285_ (.B1(_01944_),
    .Y(_00933_),
    .A1(net2470),
    .A2(net1981));
 sg13g2_nand2_1 _06286_ (.Y(_01945_),
    .A(net1708),
    .B(net1984));
 sg13g2_o21ai_1 _06287_ (.B1(_01945_),
    .Y(_00934_),
    .A1(net2468),
    .A2(net1984));
 sg13g2_nand2_1 _06288_ (.Y(_01946_),
    .A(net1744),
    .B(net1979));
 sg13g2_o21ai_1 _06289_ (.B1(_01946_),
    .Y(_00935_),
    .A1(net2461),
    .A2(net1979));
 sg13g2_nand2_1 _06290_ (.Y(_01947_),
    .A(net1616),
    .B(net1981));
 sg13g2_o21ai_1 _06291_ (.B1(_01947_),
    .Y(_00936_),
    .A1(net2459),
    .A2(net1981));
 sg13g2_nand2_1 _06292_ (.Y(_01948_),
    .A(net2951),
    .B(net1983));
 sg13g2_o21ai_1 _06293_ (.B1(_01948_),
    .Y(_00937_),
    .A1(net2452),
    .A2(net1983));
 sg13g2_nand2_1 _06294_ (.Y(_01949_),
    .A(net2821),
    .B(net1987));
 sg13g2_o21ai_1 _06295_ (.B1(_01949_),
    .Y(_00938_),
    .A1(net2447),
    .A2(net1987));
 sg13g2_nand2_1 _06296_ (.Y(_01950_),
    .A(net3006),
    .B(net1980));
 sg13g2_o21ai_1 _06297_ (.B1(_01950_),
    .Y(_00939_),
    .A1(net2440),
    .A2(net1980));
 sg13g2_nand2_1 _06298_ (.Y(_01951_),
    .A(net2838),
    .B(net1987));
 sg13g2_o21ai_1 _06299_ (.B1(_01951_),
    .Y(_00940_),
    .A1(net2435),
    .A2(net1987));
 sg13g2_nand2_1 _06300_ (.Y(_01952_),
    .A(net1674),
    .B(net1982));
 sg13g2_o21ai_1 _06301_ (.B1(_01952_),
    .Y(_00941_),
    .A1(net2433),
    .A2(net1982));
 sg13g2_nand2_1 _06302_ (.Y(_01953_),
    .A(net2804),
    .B(net1982));
 sg13g2_o21ai_1 _06303_ (.B1(_01953_),
    .Y(_00942_),
    .A1(net2423),
    .A2(net1982));
 sg13g2_nand2_1 _06304_ (.Y(_01954_),
    .A(net2900),
    .B(net1982));
 sg13g2_o21ai_1 _06305_ (.B1(_01954_),
    .Y(_00943_),
    .A1(net2419),
    .A2(net1982));
 sg13g2_nand2_1 _06306_ (.Y(_01955_),
    .A(net3100),
    .B(net1982));
 sg13g2_o21ai_1 _06307_ (.B1(_01955_),
    .Y(_00944_),
    .A1(net2415),
    .A2(net1982));
 sg13g2_nand2_1 _06308_ (.Y(_01956_),
    .A(net3114),
    .B(net1979));
 sg13g2_o21ai_1 _06309_ (.B1(_01956_),
    .Y(_00945_),
    .A1(net2412),
    .A2(net1979));
 sg13g2_nand2_1 _06310_ (.Y(_01957_),
    .A(net2938),
    .B(net1979));
 sg13g2_o21ai_1 _06311_ (.B1(_01957_),
    .Y(_00946_),
    .A1(net2402),
    .A2(net1979));
 sg13g2_nand2_1 _06312_ (.Y(_01958_),
    .A(net3041),
    .B(net1979));
 sg13g2_o21ai_1 _06313_ (.B1(_01958_),
    .Y(_00947_),
    .A1(net2400),
    .A2(net1979));
 sg13g2_nand2_1 _06314_ (.Y(_01959_),
    .A(_01616_),
    .B(_01825_));
 sg13g2_nand2_1 _06315_ (.Y(_01960_),
    .A(net2683),
    .B(net1969));
 sg13g2_o21ai_1 _06316_ (.B1(_01960_),
    .Y(_00948_),
    .A1(net2561),
    .A2(net1969));
 sg13g2_nand2_1 _06317_ (.Y(_01961_),
    .A(net2612),
    .B(net1970));
 sg13g2_o21ai_1 _06318_ (.B1(_01961_),
    .Y(_00949_),
    .A1(net2557),
    .A2(net1970));
 sg13g2_nand2_1 _06319_ (.Y(_01962_),
    .A(net3309),
    .B(net1977));
 sg13g2_o21ai_1 _06320_ (.B1(_01962_),
    .Y(_00950_),
    .A1(net2552),
    .A2(net1977));
 sg13g2_nand2_1 _06321_ (.Y(_01963_),
    .A(net2803),
    .B(net1978));
 sg13g2_o21ai_1 _06322_ (.B1(_01963_),
    .Y(_00951_),
    .A1(net2548),
    .A2(net1977));
 sg13g2_nand2_1 _06323_ (.Y(_01964_),
    .A(net2658),
    .B(net1976));
 sg13g2_o21ai_1 _06324_ (.B1(_01964_),
    .Y(_00952_),
    .A1(net2542),
    .A2(net1976));
 sg13g2_nand2_1 _06325_ (.Y(_01965_),
    .A(net2992),
    .B(net1976));
 sg13g2_o21ai_1 _06326_ (.B1(_01965_),
    .Y(_00953_),
    .A1(net2534),
    .A2(net1976));
 sg13g2_nand2_1 _06327_ (.Y(_01966_),
    .A(net2874),
    .B(net1976));
 sg13g2_o21ai_1 _06328_ (.B1(_01966_),
    .Y(_00954_),
    .A1(net2529),
    .A2(net1976));
 sg13g2_nand2_1 _06329_ (.Y(_01967_),
    .A(net2666),
    .B(net1976));
 sg13g2_o21ai_1 _06330_ (.B1(_01967_),
    .Y(_00955_),
    .A1(net2525),
    .A2(net1976));
 sg13g2_nand2_1 _06331_ (.Y(_01968_),
    .A(net2637),
    .B(net1974));
 sg13g2_o21ai_1 _06332_ (.B1(_01968_),
    .Y(_00956_),
    .A1(net2520),
    .A2(net1974));
 sg13g2_nand2_1 _06333_ (.Y(_01969_),
    .A(net3042),
    .B(net1973));
 sg13g2_o21ai_1 _06334_ (.B1(_01969_),
    .Y(_00957_),
    .A1(net2513),
    .A2(net1973));
 sg13g2_nand2_1 _06335_ (.Y(_01970_),
    .A(net3285),
    .B(net1973));
 sg13g2_o21ai_1 _06336_ (.B1(_01970_),
    .Y(_00958_),
    .A1(net2508),
    .A2(net1973));
 sg13g2_nand2_1 _06337_ (.Y(_01971_),
    .A(net1660),
    .B(net1973));
 sg13g2_o21ai_1 _06338_ (.B1(_01971_),
    .Y(_00959_),
    .A1(net2505),
    .A2(net1973));
 sg13g2_nand2_1 _06339_ (.Y(_01972_),
    .A(net2954),
    .B(net1973));
 sg13g2_o21ai_1 _06340_ (.B1(_01972_),
    .Y(_00960_),
    .A1(net2499),
    .A2(net1973));
 sg13g2_nand2_1 _06341_ (.Y(_01973_),
    .A(net3094),
    .B(net1974));
 sg13g2_o21ai_1 _06342_ (.B1(_01973_),
    .Y(_00961_),
    .A1(net2493),
    .A2(net1974));
 sg13g2_nand2_1 _06343_ (.Y(_01974_),
    .A(net2894),
    .B(net1969));
 sg13g2_o21ai_1 _06344_ (.B1(_01974_),
    .Y(_00962_),
    .A1(net2487),
    .A2(net1969));
 sg13g2_nand2_1 _06345_ (.Y(_01975_),
    .A(net3275),
    .B(net1975));
 sg13g2_o21ai_1 _06346_ (.B1(_01975_),
    .Y(_00963_),
    .A1(net2482),
    .A2(net1975));
 sg13g2_nand2_1 _06347_ (.Y(_01976_),
    .A(net2758),
    .B(net1975));
 sg13g2_o21ai_1 _06348_ (.B1(_01976_),
    .Y(_00964_),
    .A1(net2475),
    .A2(net1975));
 sg13g2_nand2_1 _06349_ (.Y(_01977_),
    .A(net3003),
    .B(net1969));
 sg13g2_o21ai_1 _06350_ (.B1(_01977_),
    .Y(_00965_),
    .A1(net2473),
    .A2(net1969));
 sg13g2_nand2_1 _06351_ (.Y(_01978_),
    .A(net1527),
    .B(net1975));
 sg13g2_o21ai_1 _06352_ (.B1(_01978_),
    .Y(_00966_),
    .A1(net2465),
    .A2(net1975));
 sg13g2_nand2_1 _06353_ (.Y(_01979_),
    .A(net1724),
    .B(net1972));
 sg13g2_o21ai_1 _06354_ (.B1(_01979_),
    .Y(_00967_),
    .A1(net2463),
    .A2(net1972));
 sg13g2_nand2_1 _06355_ (.Y(_01980_),
    .A(net3283),
    .B(net1969));
 sg13g2_o21ai_1 _06356_ (.B1(_01980_),
    .Y(_00968_),
    .A1(net2459),
    .A2(net1972));
 sg13g2_nand2_1 _06357_ (.Y(_01981_),
    .A(net1742),
    .B(net1971));
 sg13g2_o21ai_1 _06358_ (.B1(_01981_),
    .Y(_00969_),
    .A1(net2454),
    .A2(net1971));
 sg13g2_nand2_1 _06359_ (.Y(_01982_),
    .A(net3295),
    .B(net1977));
 sg13g2_o21ai_1 _06360_ (.B1(_01982_),
    .Y(_00970_),
    .A1(net2446),
    .A2(net1977));
 sg13g2_nand2_1 _06361_ (.Y(_01983_),
    .A(net1458),
    .B(net1968));
 sg13g2_o21ai_1 _06362_ (.B1(_01983_),
    .Y(_00971_),
    .A1(net2441),
    .A2(net1968));
 sg13g2_nand2_1 _06363_ (.Y(_01984_),
    .A(net3291),
    .B(net1977));
 sg13g2_o21ai_1 _06364_ (.B1(_01984_),
    .Y(_00972_),
    .A1(net2434),
    .A2(net1977));
 sg13g2_nand2_1 _06365_ (.Y(_01985_),
    .A(net3193),
    .B(net1970));
 sg13g2_o21ai_1 _06366_ (.B1(_01985_),
    .Y(_00973_),
    .A1(net2430),
    .A2(net1970));
 sg13g2_nand2_1 _06367_ (.Y(_01986_),
    .A(net3058),
    .B(net1971));
 sg13g2_o21ai_1 _06368_ (.B1(_01986_),
    .Y(_00974_),
    .A1(net2427),
    .A2(net1971));
 sg13g2_nand2_1 _06369_ (.Y(_01987_),
    .A(net3323),
    .B(net1970));
 sg13g2_o21ai_1 _06370_ (.B1(_01987_),
    .Y(_00975_),
    .A1(net2421),
    .A2(net1970));
 sg13g2_nand2_1 _06371_ (.Y(_01988_),
    .A(net2977),
    .B(net1970));
 sg13g2_o21ai_1 _06372_ (.B1(_01988_),
    .Y(_00976_),
    .A1(net2414),
    .A2(net1970));
 sg13g2_nand2_1 _06373_ (.Y(_01989_),
    .A(net2906),
    .B(net1968));
 sg13g2_o21ai_1 _06374_ (.B1(_01989_),
    .Y(_00977_),
    .A1(net2408),
    .A2(net1968));
 sg13g2_nand2_1 _06375_ (.Y(_01990_),
    .A(net1545),
    .B(net1968));
 sg13g2_o21ai_1 _06376_ (.B1(_01990_),
    .Y(_00978_),
    .A1(net2405),
    .A2(net1968));
 sg13g2_nand2_1 _06377_ (.Y(_01991_),
    .A(net3209),
    .B(net1968));
 sg13g2_o21ai_1 _06378_ (.B1(_01991_),
    .Y(_00979_),
    .A1(net2398),
    .A2(net1968));
 sg13g2_nor2_2 _06379_ (.A(_01532_),
    .B(_01824_),
    .Y(_01992_));
 sg13g2_nand2b_1 _06380_ (.Y(_01993_),
    .B(_01533_),
    .A_N(_01824_));
 sg13g2_nand2_2 _06381_ (.Y(_01994_),
    .A(_01751_),
    .B(_01992_));
 sg13g2_nand2_1 _06382_ (.Y(_01995_),
    .A(net3197),
    .B(net1958));
 sg13g2_o21ai_1 _06383_ (.B1(_01995_),
    .Y(_00980_),
    .A1(net2562),
    .A2(net1958));
 sg13g2_nand2_1 _06384_ (.Y(_01996_),
    .A(net3155),
    .B(net1961));
 sg13g2_o21ai_1 _06385_ (.B1(_01996_),
    .Y(_00981_),
    .A1(net2555),
    .A2(net1961));
 sg13g2_nand2_1 _06386_ (.Y(_01997_),
    .A(net1555),
    .B(net1966));
 sg13g2_o21ai_1 _06387_ (.B1(_01997_),
    .Y(_00982_),
    .A1(net2552),
    .A2(net1966));
 sg13g2_nand2_1 _06388_ (.Y(_01998_),
    .A(net1714),
    .B(net1965));
 sg13g2_o21ai_1 _06389_ (.B1(_01998_),
    .Y(_00983_),
    .A1(net2546),
    .A2(net1965));
 sg13g2_nand2_1 _06390_ (.Y(_01999_),
    .A(net2770),
    .B(net1965));
 sg13g2_o21ai_1 _06391_ (.B1(_01999_),
    .Y(_00984_),
    .A1(net2541),
    .A2(net1965));
 sg13g2_nand2_1 _06392_ (.Y(_02000_),
    .A(net2852),
    .B(net1967));
 sg13g2_o21ai_1 _06393_ (.B1(_02000_),
    .Y(_00985_),
    .A1(net2536),
    .A2(net1966));
 sg13g2_nand2_1 _06394_ (.Y(_02001_),
    .A(net1504),
    .B(net1965));
 sg13g2_o21ai_1 _06395_ (.B1(_02001_),
    .Y(_00986_),
    .A1(net2530),
    .A2(net1965));
 sg13g2_nand2_1 _06396_ (.Y(_02002_),
    .A(net2795),
    .B(net1965));
 sg13g2_o21ai_1 _06397_ (.B1(_02002_),
    .Y(_00987_),
    .A1(net2526),
    .A2(net1965));
 sg13g2_nand2_1 _06398_ (.Y(_02003_),
    .A(net1484),
    .B(net1964));
 sg13g2_o21ai_1 _06399_ (.B1(_02003_),
    .Y(_00988_),
    .A1(net2521),
    .A2(net1964));
 sg13g2_nand2_1 _06400_ (.Y(_02004_),
    .A(net1721),
    .B(net1964));
 sg13g2_o21ai_1 _06401_ (.B1(_02004_),
    .Y(_00989_),
    .A1(net2514),
    .A2(net1964));
 sg13g2_nand2_1 _06402_ (.Y(_02005_),
    .A(net2751),
    .B(net1964));
 sg13g2_o21ai_1 _06403_ (.B1(_02005_),
    .Y(_00990_),
    .A1(net2509),
    .A2(net1964));
 sg13g2_nand2_1 _06404_ (.Y(_02006_),
    .A(net2878),
    .B(net1963));
 sg13g2_o21ai_1 _06405_ (.B1(_02006_),
    .Y(_00991_),
    .A1(net2506),
    .A2(net1963));
 sg13g2_nand2_1 _06406_ (.Y(_02007_),
    .A(net3192),
    .B(net1964));
 sg13g2_o21ai_1 _06407_ (.B1(_02007_),
    .Y(_00992_),
    .A1(net2501),
    .A2(net1964));
 sg13g2_nand2_1 _06408_ (.Y(_02008_),
    .A(net2922),
    .B(net1966));
 sg13g2_o21ai_1 _06409_ (.B1(_02008_),
    .Y(_00993_),
    .A1(net2493),
    .A2(net1966));
 sg13g2_nand2_1 _06410_ (.Y(_02009_),
    .A(net2680),
    .B(net1959));
 sg13g2_o21ai_1 _06411_ (.B1(_02009_),
    .Y(_00994_),
    .A1(net2489),
    .A2(net1962));
 sg13g2_nand2_1 _06412_ (.Y(_02010_),
    .A(net1449),
    .B(net1963));
 sg13g2_o21ai_1 _06413_ (.B1(_02010_),
    .Y(_00995_),
    .A1(net2484),
    .A2(net1963));
 sg13g2_nand2_1 _06414_ (.Y(_02011_),
    .A(net1706),
    .B(net1963));
 sg13g2_o21ai_1 _06415_ (.B1(_02011_),
    .Y(_00996_),
    .A1(net2475),
    .A2(net1963));
 sg13g2_nand2_1 _06416_ (.Y(_02012_),
    .A(net1510),
    .B(net1959));
 sg13g2_o21ai_1 _06417_ (.B1(_02012_),
    .Y(_00997_),
    .A1(net2471),
    .A2(net1959));
 sg13g2_nand2_1 _06418_ (.Y(_02013_),
    .A(net2832),
    .B(net1963));
 sg13g2_o21ai_1 _06419_ (.B1(_02013_),
    .Y(_00998_),
    .A1(net2466),
    .A2(net1963));
 sg13g2_nand2_1 _06420_ (.Y(_02014_),
    .A(net1611),
    .B(net1958));
 sg13g2_o21ai_1 _06421_ (.B1(_02014_),
    .Y(_00999_),
    .A1(net2460),
    .A2(net1958));
 sg13g2_nand2_1 _06422_ (.Y(_02015_),
    .A(net2670),
    .B(net1959));
 sg13g2_o21ai_1 _06423_ (.B1(_02015_),
    .Y(_01000_),
    .A1(net2456),
    .A2(net1959));
 sg13g2_nand2_1 _06424_ (.Y(_02016_),
    .A(net3017),
    .B(net1961));
 sg13g2_o21ai_1 _06425_ (.B1(_02016_),
    .Y(_01001_),
    .A1(net2451),
    .A2(net1962));
 sg13g2_nand2_1 _06426_ (.Y(_02017_),
    .A(net3210),
    .B(net1966));
 sg13g2_o21ai_1 _06427_ (.B1(_02017_),
    .Y(_01002_),
    .A1(net2447),
    .A2(net1966));
 sg13g2_nand2_1 _06428_ (.Y(_02018_),
    .A(net1487),
    .B(net1960));
 sg13g2_o21ai_1 _06429_ (.B1(_02018_),
    .Y(_01003_),
    .A1(net2442),
    .A2(net1960));
 sg13g2_nand2_1 _06430_ (.Y(_02019_),
    .A(net2790),
    .B(net1961));
 sg13g2_o21ai_1 _06431_ (.B1(_02019_),
    .Y(_01004_),
    .A1(net2438),
    .A2(net1961));
 sg13g2_nand2_1 _06432_ (.Y(_02020_),
    .A(net1653),
    .B(net1960));
 sg13g2_o21ai_1 _06433_ (.B1(_02020_),
    .Y(_01005_),
    .A1(net2431),
    .A2(net1960));
 sg13g2_nand2_1 _06434_ (.Y(_02021_),
    .A(net1469),
    .B(net1961));
 sg13g2_o21ai_1 _06435_ (.B1(_02021_),
    .Y(_01006_),
    .A1(net2424),
    .A2(net1961));
 sg13g2_nand2_1 _06436_ (.Y(_02022_),
    .A(net2767),
    .B(net1960));
 sg13g2_o21ai_1 _06437_ (.B1(_02022_),
    .Y(_01007_),
    .A1(net2420),
    .A2(net1960));
 sg13g2_nand2_1 _06438_ (.Y(_02023_),
    .A(net2715),
    .B(net1960));
 sg13g2_o21ai_1 _06439_ (.B1(_02023_),
    .Y(_01008_),
    .A1(net2416),
    .A2(net1960));
 sg13g2_nand2_1 _06440_ (.Y(_02024_),
    .A(net3104),
    .B(net1959));
 sg13g2_o21ai_1 _06441_ (.B1(_02024_),
    .Y(_01009_),
    .A1(net2411),
    .A2(net1959));
 sg13g2_nand2_1 _06442_ (.Y(_02025_),
    .A(net3095),
    .B(net1958));
 sg13g2_o21ai_1 _06443_ (.B1(_02025_),
    .Y(_01010_),
    .A1(net2402),
    .A2(net1958));
 sg13g2_nand2_1 _06444_ (.Y(_02026_),
    .A(net1569),
    .B(net1958));
 sg13g2_o21ai_1 _06445_ (.B1(_02026_),
    .Y(_01011_),
    .A1(net2399),
    .A2(net1958));
 sg13g2_nor2b_1 _06446_ (.A(_01387_),
    .B_N(_01378_),
    .Y(_02027_));
 sg13g2_a21o_1 _06447_ (.A2(_01387_),
    .A1(_01384_),
    .B1(_01666_),
    .X(_02028_));
 sg13g2_nor4_1 _06448_ (.A(_01378_),
    .B(_01385_),
    .C(net2372),
    .D(_02028_),
    .Y(_02029_));
 sg13g2_a22oi_1 _06449_ (.Y(_02030_),
    .B1(_02029_),
    .B2(net2571),
    .A2(_01668_),
    .A1(_01416_));
 sg13g2_or2_1 _06450_ (.X(_02031_),
    .B(_01668_),
    .A(_01371_));
 sg13g2_a221oi_1 _06451_ (.B2(_01666_),
    .C1(_02029_),
    .B1(_02031_),
    .A1(\cpu.arbiter.i_wb_cpu_dbus_dat[0] ),
    .Y(_02032_),
    .A2(net2389));
 sg13g2_nor2_1 _06452_ (.A(net2361),
    .B(_02032_),
    .Y(_02033_));
 sg13g2_a21oi_1 _06453_ (.A1(net6),
    .A2(net2361),
    .Y(_02034_),
    .B1(_02033_));
 sg13g2_nor2_1 _06454_ (.A(net3594),
    .B(net2323),
    .Y(_02035_));
 sg13g2_a21oi_1 _06455_ (.A1(net2323),
    .A2(_02034_),
    .Y(_01012_),
    .B1(_02035_));
 sg13g2_or4_1 _06456_ (.A(_01386_),
    .B(net2372),
    .C(_02027_),
    .D(_02028_),
    .X(_02036_));
 sg13g2_a21oi_1 _06457_ (.A1(net3652),
    .A2(net2389),
    .Y(_02037_),
    .B1(_02031_));
 sg13g2_a22oi_1 _06458_ (.Y(_02038_),
    .B1(_02036_),
    .B2(_02037_),
    .A2(net2361),
    .A1(_01354_));
 sg13g2_mux2_1 _06459_ (.A0(net3668),
    .A1(_02038_),
    .S(net2323),
    .X(_01013_));
 sg13g2_a21oi_1 _06460_ (.A1(_01355_),
    .A2(net2391),
    .Y(_02039_),
    .B1(net2372));
 sg13g2_o21ai_1 _06461_ (.B1(_02039_),
    .Y(_02040_),
    .A1(net3544),
    .A2(net2391));
 sg13g2_a22oi_1 _06462_ (.Y(_02041_),
    .B1(net2389),
    .B2(net3576),
    .A2(net2362),
    .A1(\cpu.arbiter.i_wb_mem_rdt[1] ));
 sg13g2_and2_1 _06463_ (.A(_02040_),
    .B(_02041_),
    .X(_02042_));
 sg13g2_nor2_1 _06464_ (.A(net3637),
    .B(net2322),
    .Y(_02043_));
 sg13g2_a21oi_1 _06465_ (.A1(net2322),
    .A2(_02042_),
    .Y(_01014_),
    .B1(_02043_));
 sg13g2_nor2_1 _06466_ (.A(net3534),
    .B(net2391),
    .Y(_02044_));
 sg13g2_nor2_1 _06467_ (.A(net3676),
    .B(net2393),
    .Y(_02045_));
 sg13g2_nor3_1 _06468_ (.A(net2372),
    .B(_02044_),
    .C(_02045_),
    .Y(_02046_));
 sg13g2_a221oi_1 _06469_ (.B2(net3621),
    .C1(_02046_),
    .B1(net2389),
    .A1(net3637),
    .Y(_02047_),
    .A2(net2361));
 sg13g2_nor2_1 _06470_ (.A(net3690),
    .B(net2323),
    .Y(_02048_));
 sg13g2_a21oi_1 _06471_ (.A1(net2323),
    .A2(_02047_),
    .Y(_01015_),
    .B1(_02048_));
 sg13g2_nor2_1 _06472_ (.A(net3630),
    .B(net2391),
    .Y(_02049_));
 sg13g2_nor2_1 _06473_ (.A(net3703),
    .B(net2393),
    .Y(_02050_));
 sg13g2_nor3_1 _06474_ (.A(net2372),
    .B(_02049_),
    .C(_02050_),
    .Y(_02051_));
 sg13g2_a221oi_1 _06475_ (.B2(net3635),
    .C1(_02051_),
    .B1(net2389),
    .A1(net3690),
    .Y(_02052_),
    .A2(net2361));
 sg13g2_nor2_1 _06476_ (.A(net3718),
    .B(net2322),
    .Y(_02053_));
 sg13g2_a21oi_1 _06477_ (.A1(net2322),
    .A2(_02052_),
    .Y(_01016_),
    .B1(_02053_));
 sg13g2_nor2_1 _06478_ (.A(net3634),
    .B(net2391),
    .Y(_02054_));
 sg13g2_nor2_1 _06479_ (.A(net3670),
    .B(_01655_),
    .Y(_02055_));
 sg13g2_nor3_1 _06480_ (.A(net2372),
    .B(_02054_),
    .C(_02055_),
    .Y(_02056_));
 sg13g2_a221oi_1 _06481_ (.B2(\cpu.arbiter.i_wb_cpu_dbus_dat[5] ),
    .C1(_02056_),
    .B1(net2389),
    .A1(\cpu.arbiter.i_wb_mem_rdt[4] ),
    .Y(_02057_),
    .A2(net2361));
 sg13g2_nor2_1 _06482_ (.A(net3678),
    .B(net2322),
    .Y(_02058_));
 sg13g2_a21oi_1 _06483_ (.A1(net2322),
    .A2(_02057_),
    .Y(_01017_),
    .B1(_02058_));
 sg13g2_nor2_1 _06484_ (.A(net3596),
    .B(net2391),
    .Y(_02059_));
 sg13g2_nor2_1 _06485_ (.A(net3654),
    .B(net2393),
    .Y(_02060_));
 sg13g2_nor3_1 _06486_ (.A(net2372),
    .B(_02059_),
    .C(_02060_),
    .Y(_02061_));
 sg13g2_a221oi_1 _06487_ (.B2(net3632),
    .C1(_02061_),
    .B1(net2389),
    .A1(net3678),
    .Y(_02062_),
    .A2(net2361));
 sg13g2_nor2_1 _06488_ (.A(net3683),
    .B(net2323),
    .Y(_02063_));
 sg13g2_a21oi_1 _06489_ (.A1(net2322),
    .A2(_02062_),
    .Y(_01018_),
    .B1(_02063_));
 sg13g2_nor2_1 _06490_ (.A(net3500),
    .B(net2392),
    .Y(_02064_));
 sg13g2_nor2_1 _06491_ (.A(\cpu.arbiter.i_wb_cpu_dbus_adr[7] ),
    .B(net2393),
    .Y(_02065_));
 sg13g2_nor3_1 _06492_ (.A(_01673_),
    .B(_02064_),
    .C(_02065_),
    .Y(_02066_));
 sg13g2_a221oi_1 _06493_ (.B2(net3648),
    .C1(_02066_),
    .B1(_01669_),
    .A1(net3683),
    .Y(_02067_),
    .A2(net2361));
 sg13g2_nor2_1 _06494_ (.A(net3749),
    .B(net2324),
    .Y(_02068_));
 sg13g2_a21oi_1 _06495_ (.A1(net2322),
    .A2(_02067_),
    .Y(_01019_),
    .B1(_02068_));
 sg13g2_nor2_1 _06496_ (.A(net3692),
    .B(net2321),
    .Y(_02069_));
 sg13g2_nor2_1 _06497_ (.A(net3664),
    .B(net2393),
    .Y(_02070_));
 sg13g2_nor2_1 _06498_ (.A(net3527),
    .B(_01656_),
    .Y(_02071_));
 sg13g2_nor3_1 _06499_ (.A(net2372),
    .B(_02070_),
    .C(_02071_),
    .Y(_02072_));
 sg13g2_a221oi_1 _06500_ (.B2(\cpu.arbiter.i_wb_cpu_dbus_dat[8] ),
    .C1(_02072_),
    .B1(net2389),
    .A1(\cpu.arbiter.i_wb_mem_rdt[7] ),
    .Y(_02073_),
    .A2(net2362));
 sg13g2_a21oi_1 _06501_ (.A1(net2321),
    .A2(_02073_),
    .Y(_01020_),
    .B1(_02069_));
 sg13g2_and2_1 _06502_ (.A(net3667),
    .B(net2392),
    .X(_02074_));
 sg13g2_a21oi_1 _06503_ (.A1(net3666),
    .A2(net2394),
    .Y(_02075_),
    .B1(_02074_));
 sg13g2_a22oi_1 _06504_ (.Y(_02076_),
    .B1(net2390),
    .B2(net3552),
    .A2(net2360),
    .A1(net3692));
 sg13g2_o21ai_1 _06505_ (.B1(_02076_),
    .Y(_02077_),
    .A1(net2373),
    .A2(_02075_));
 sg13g2_nand2_1 _06506_ (.Y(_02078_),
    .A(net2321),
    .B(_02077_));
 sg13g2_o21ai_1 _06507_ (.B1(_02078_),
    .Y(_01021_),
    .A1(_01356_),
    .A2(net2321));
 sg13g2_nor2_1 _06508_ (.A(net3626),
    .B(net2320),
    .Y(_02079_));
 sg13g2_nor2_1 _06509_ (.A(\cpu.arbiter.i_wb_cpu_dbus_adr[10] ),
    .B(net2394),
    .Y(_02080_));
 sg13g2_nor2_1 _06510_ (.A(net3569),
    .B(net2392),
    .Y(_02081_));
 sg13g2_nor3_1 _06511_ (.A(net2373),
    .B(_02080_),
    .C(_02081_),
    .Y(_02082_));
 sg13g2_a221oi_1 _06512_ (.B2(net3546),
    .C1(_02082_),
    .B1(net2390),
    .A1(\cpu.arbiter.i_wb_mem_rdt[9] ),
    .Y(_02083_),
    .A2(net2360));
 sg13g2_a21oi_1 _06513_ (.A1(net2320),
    .A2(_02083_),
    .Y(_01022_),
    .B1(_02079_));
 sg13g2_and2_1 _06514_ (.A(net3662),
    .B(net2392),
    .X(_02084_));
 sg13g2_a21oi_1 _06515_ (.A1(net3567),
    .A2(net2394),
    .Y(_02085_),
    .B1(_02084_));
 sg13g2_a22oi_1 _06516_ (.Y(_02086_),
    .B1(net2390),
    .B2(net3610),
    .A2(net2360),
    .A1(net3626));
 sg13g2_o21ai_1 _06517_ (.B1(_02086_),
    .Y(_02087_),
    .A1(net2373),
    .A2(_02085_));
 sg13g2_nand2_1 _06518_ (.Y(_02088_),
    .A(net2319),
    .B(_02087_));
 sg13g2_o21ai_1 _06519_ (.B1(_02088_),
    .Y(_01023_),
    .A1(_01358_),
    .A2(net2319));
 sg13g2_nor2_1 _06520_ (.A(net3542),
    .B(net2392),
    .Y(_02089_));
 sg13g2_nor2_1 _06521_ (.A(net3685),
    .B(net2394),
    .Y(_02090_));
 sg13g2_nor3_1 _06522_ (.A(net2373),
    .B(_02089_),
    .C(_02090_),
    .Y(_02091_));
 sg13g2_a221oi_1 _06523_ (.B2(net3548),
    .C1(_02091_),
    .B1(net2390),
    .A1(net3713),
    .Y(_02092_),
    .A2(net2359));
 sg13g2_nor2_1 _06524_ (.A(net3669),
    .B(net2319),
    .Y(_02093_));
 sg13g2_a21oi_1 _06525_ (.A1(net2319),
    .A2(_02092_),
    .Y(_01024_),
    .B1(_02093_));
 sg13g2_nor2_1 _06526_ (.A(net3490),
    .B(net2392),
    .Y(_02094_));
 sg13g2_nor2_1 _06527_ (.A(\cpu.arbiter.i_wb_cpu_dbus_adr[13] ),
    .B(net2394),
    .Y(_02095_));
 sg13g2_nor3_1 _06528_ (.A(net2373),
    .B(_02094_),
    .C(_02095_),
    .Y(_02096_));
 sg13g2_a221oi_1 _06529_ (.B2(net3617),
    .C1(_02096_),
    .B1(net2390),
    .A1(net3669),
    .Y(_02097_),
    .A2(net2359));
 sg13g2_nor2_1 _06530_ (.A(net3694),
    .B(net2319),
    .Y(_02098_));
 sg13g2_a21oi_1 _06531_ (.A1(net2319),
    .A2(_02097_),
    .Y(_01025_),
    .B1(_02098_));
 sg13g2_nor2_1 _06532_ (.A(net3479),
    .B(net2392),
    .Y(_02099_));
 sg13g2_nor2_1 _06533_ (.A(\cpu.arbiter.i_wb_cpu_dbus_adr[14] ),
    .B(net2394),
    .Y(_02100_));
 sg13g2_nor3_1 _06534_ (.A(net2373),
    .B(_02099_),
    .C(_02100_),
    .Y(_02101_));
 sg13g2_a221oi_1 _06535_ (.B2(\cpu.arbiter.i_wb_cpu_dbus_dat[14] ),
    .C1(_02101_),
    .B1(net2390),
    .A1(\cpu.arbiter.i_wb_mem_rdt[13] ),
    .Y(_02102_),
    .A2(net2359));
 sg13g2_nor2_1 _06536_ (.A(net3628),
    .B(net2319),
    .Y(_02103_));
 sg13g2_a21oi_1 _06537_ (.A1(net2319),
    .A2(_02102_),
    .Y(_01026_),
    .B1(_02103_));
 sg13g2_nor2_1 _06538_ (.A(net3741),
    .B(net2320),
    .Y(_02104_));
 sg13g2_nor2_1 _06539_ (.A(net3684),
    .B(net2394),
    .Y(_02105_));
 sg13g2_nor2_1 _06540_ (.A(net3608),
    .B(net2392),
    .Y(_02106_));
 sg13g2_nor3_1 _06541_ (.A(net2373),
    .B(_02105_),
    .C(_02106_),
    .Y(_02107_));
 sg13g2_a221oi_1 _06542_ (.B2(net3598),
    .C1(_02107_),
    .B1(net2390),
    .A1(net3628),
    .Y(_02108_),
    .A2(net2360));
 sg13g2_a21oi_1 _06543_ (.A1(net2320),
    .A2(_02108_),
    .Y(_01027_),
    .B1(_02104_));
 sg13g2_nand2b_2 _06544_ (.Y(_02109_),
    .B(_01751_),
    .A_N(net2307));
 sg13g2_nand2_1 _06545_ (.Y(_02110_),
    .A(net1572),
    .B(net1947));
 sg13g2_o21ai_1 _06546_ (.B1(_02110_),
    .Y(_01028_),
    .A1(net2560),
    .A2(net1947));
 sg13g2_nand2_1 _06547_ (.Y(_02111_),
    .A(net3303),
    .B(net1949));
 sg13g2_o21ai_1 _06548_ (.B1(_02111_),
    .Y(_01029_),
    .A1(net2556),
    .A2(net1950));
 sg13g2_nand2_1 _06549_ (.Y(_02112_),
    .A(net3185),
    .B(net1957));
 sg13g2_o21ai_1 _06550_ (.B1(_02112_),
    .Y(_01030_),
    .A1(net2554),
    .A2(net1957));
 sg13g2_nand2_1 _06551_ (.Y(_02113_),
    .A(net2681),
    .B(net1955));
 sg13g2_o21ai_1 _06552_ (.B1(_02113_),
    .Y(_01031_),
    .A1(net2544),
    .A2(net1955));
 sg13g2_nand2_1 _06553_ (.Y(_02114_),
    .A(net2836),
    .B(net1956));
 sg13g2_o21ai_1 _06554_ (.B1(_02114_),
    .Y(_01032_),
    .A1(net2538),
    .A2(net1956));
 sg13g2_nand2_1 _06555_ (.Y(_02115_),
    .A(net2610),
    .B(net1956));
 sg13g2_o21ai_1 _06556_ (.B1(_02115_),
    .Y(_01033_),
    .A1(net2533),
    .A2(net1956));
 sg13g2_nand2_1 _06557_ (.Y(_02116_),
    .A(net1661),
    .B(net1955));
 sg13g2_o21ai_1 _06558_ (.B1(_02116_),
    .Y(_01034_),
    .A1(net2529),
    .A2(net1955));
 sg13g2_nand2_1 _06559_ (.Y(_02117_),
    .A(net3293),
    .B(net1955));
 sg13g2_o21ai_1 _06560_ (.B1(_02117_),
    .Y(_01035_),
    .A1(net2523),
    .A2(net1955));
 sg13g2_nand2_1 _06561_ (.Y(_02118_),
    .A(net1612),
    .B(net1952));
 sg13g2_o21ai_1 _06562_ (.B1(_02118_),
    .Y(_01036_),
    .A1(net2518),
    .A2(net1952));
 sg13g2_nand2_1 _06563_ (.Y(_02119_),
    .A(net2629),
    .B(net1952));
 sg13g2_o21ai_1 _06564_ (.B1(_02119_),
    .Y(_01037_),
    .A1(net2513),
    .A2(net1952));
 sg13g2_nand2_1 _06565_ (.Y(_02120_),
    .A(net1501),
    .B(net1953));
 sg13g2_o21ai_1 _06566_ (.B1(_02120_),
    .Y(_01038_),
    .A1(net2507),
    .A2(net1953));
 sg13g2_nand2_1 _06567_ (.Y(_02121_),
    .A(net3250),
    .B(net1952));
 sg13g2_o21ai_1 _06568_ (.B1(_02121_),
    .Y(_01039_),
    .A1(net2502),
    .A2(net1952));
 sg13g2_nand2_1 _06569_ (.Y(_02122_),
    .A(net3160),
    .B(net1952));
 sg13g2_o21ai_1 _06570_ (.B1(_02122_),
    .Y(_01040_),
    .A1(net2496),
    .A2(net1952));
 sg13g2_nand2_1 _06571_ (.Y(_02123_),
    .A(net1516),
    .B(net1953));
 sg13g2_o21ai_1 _06572_ (.B1(_02123_),
    .Y(_01041_),
    .A1(net2492),
    .A2(net1953));
 sg13g2_nand2_1 _06573_ (.Y(_02124_),
    .A(net1419),
    .B(net1948));
 sg13g2_o21ai_1 _06574_ (.B1(_02124_),
    .Y(_01042_),
    .A1(net2486),
    .A2(net1948));
 sg13g2_nand2_1 _06575_ (.Y(_02125_),
    .A(net3059),
    .B(net1954));
 sg13g2_o21ai_1 _06576_ (.B1(_02125_),
    .Y(_01043_),
    .A1(net2481),
    .A2(net1954));
 sg13g2_nand2_1 _06577_ (.Y(_02126_),
    .A(net3190),
    .B(net1955));
 sg13g2_o21ai_1 _06578_ (.B1(_02126_),
    .Y(_01044_),
    .A1(net2479),
    .A2(net1955));
 sg13g2_nand2_1 _06579_ (.Y(_02127_),
    .A(net1491),
    .B(net1954));
 sg13g2_o21ai_1 _06580_ (.B1(_02127_),
    .Y(_01045_),
    .A1(net2470),
    .A2(net1954));
 sg13g2_nand2_1 _06581_ (.Y(_02128_),
    .A(net2897),
    .B(net1954));
 sg13g2_o21ai_1 _06582_ (.B1(_02128_),
    .Y(_01046_),
    .A1(net2465),
    .A2(net1954));
 sg13g2_nand2_1 _06583_ (.Y(_02129_),
    .A(net1434),
    .B(net1948));
 sg13g2_o21ai_1 _06584_ (.B1(_02129_),
    .Y(_01047_),
    .A1(net2464),
    .A2(net1948));
 sg13g2_nand2_1 _06585_ (.Y(_02130_),
    .A(net2606),
    .B(net1948));
 sg13g2_o21ai_1 _06586_ (.B1(_02130_),
    .Y(_01048_),
    .A1(net2455),
    .A2(net1948));
 sg13g2_nand2_1 _06587_ (.Y(_02131_),
    .A(net1689),
    .B(net1949));
 sg13g2_o21ai_1 _06588_ (.B1(_02131_),
    .Y(_01049_),
    .A1(net2451),
    .A2(net1950));
 sg13g2_nand2_1 _06589_ (.Y(_02132_),
    .A(net2915),
    .B(net1957));
 sg13g2_o21ai_1 _06590_ (.B1(_02132_),
    .Y(_01050_),
    .A1(net2445),
    .A2(net1957));
 sg13g2_nand2_1 _06591_ (.Y(_02133_),
    .A(net3229),
    .B(net1948));
 sg13g2_o21ai_1 _06592_ (.B1(_02133_),
    .Y(_01051_),
    .A1(net2439),
    .A2(net1948));
 sg13g2_nand2_1 _06593_ (.Y(_02134_),
    .A(net3057),
    .B(net1957));
 sg13g2_o21ai_1 _06594_ (.B1(_02134_),
    .Y(_01052_),
    .A1(net2436),
    .A2(net1957));
 sg13g2_nand2_1 _06595_ (.Y(_02135_),
    .A(net1464),
    .B(net1949));
 sg13g2_o21ai_1 _06596_ (.B1(_02135_),
    .Y(_01053_),
    .A1(net2429),
    .A2(net1949));
 sg13g2_nand2_1 _06597_ (.Y(_02136_),
    .A(net3205),
    .B(net1950));
 sg13g2_o21ai_1 _06598_ (.B1(_02136_),
    .Y(_01054_),
    .A1(net2425),
    .A2(net1950));
 sg13g2_nand2_1 _06599_ (.Y(_02137_),
    .A(net1496),
    .B(net1949));
 sg13g2_o21ai_1 _06600_ (.B1(_02137_),
    .Y(_01055_),
    .A1(net2418),
    .A2(net1949));
 sg13g2_nand2_1 _06601_ (.Y(_02138_),
    .A(net1671),
    .B(net1949));
 sg13g2_o21ai_1 _06602_ (.B1(_02138_),
    .Y(_01056_),
    .A1(net2413),
    .A2(net1949));
 sg13g2_nand2_1 _06603_ (.Y(_02139_),
    .A(net2869),
    .B(net1947));
 sg13g2_o21ai_1 _06604_ (.B1(_02139_),
    .Y(_01057_),
    .A1(net2410),
    .A2(net1947));
 sg13g2_nand2_1 _06605_ (.Y(_02140_),
    .A(net1723),
    .B(net1947));
 sg13g2_o21ai_1 _06606_ (.B1(_02140_),
    .Y(_01058_),
    .A1(net2403),
    .A2(net1947));
 sg13g2_nand2_1 _06607_ (.Y(_02141_),
    .A(net2703),
    .B(net1947));
 sg13g2_o21ai_1 _06608_ (.B1(_02141_),
    .Y(_01059_),
    .A1(net2397),
    .A2(net1947));
 sg13g2_nand2_2 _06609_ (.Y(_02142_),
    .A(_01616_),
    .B(_01992_));
 sg13g2_nand2_1 _06610_ (.Y(_02143_),
    .A(net2719),
    .B(net1938));
 sg13g2_o21ai_1 _06611_ (.B1(_02143_),
    .Y(_01060_),
    .A1(net2562),
    .A2(net1938));
 sg13g2_nand2_1 _06612_ (.Y(_02144_),
    .A(net1593),
    .B(net1940));
 sg13g2_o21ai_1 _06613_ (.B1(_02144_),
    .Y(_01061_),
    .A1(net2558),
    .A2(net1940));
 sg13g2_nand2_1 _06614_ (.Y(_02145_),
    .A(net1585),
    .B(net1945));
 sg13g2_o21ai_1 _06615_ (.B1(_02145_),
    .Y(_01062_),
    .A1(net2552),
    .A2(net1945));
 sg13g2_nand2_1 _06616_ (.Y(_02146_),
    .A(net2687),
    .B(net1944));
 sg13g2_o21ai_1 _06617_ (.B1(_02146_),
    .Y(_01063_),
    .A1(net2546),
    .A2(net1944));
 sg13g2_nand2_1 _06618_ (.Y(_02147_),
    .A(net2936),
    .B(net1944));
 sg13g2_o21ai_1 _06619_ (.B1(_02147_),
    .Y(_01064_),
    .A1(net2542),
    .A2(net1944));
 sg13g2_nand2_1 _06620_ (.Y(_02148_),
    .A(net3237),
    .B(net1946));
 sg13g2_o21ai_1 _06621_ (.B1(_02148_),
    .Y(_01065_),
    .A1(net2536),
    .A2(net1945));
 sg13g2_nand2_1 _06622_ (.Y(_02149_),
    .A(net1739),
    .B(net1944));
 sg13g2_o21ai_1 _06623_ (.B1(_02149_),
    .Y(_01066_),
    .A1(net2530),
    .A2(net1944));
 sg13g2_nand2_1 _06624_ (.Y(_02150_),
    .A(net1424),
    .B(net1944));
 sg13g2_o21ai_1 _06625_ (.B1(_02150_),
    .Y(_01067_),
    .A1(net2526),
    .A2(net1944));
 sg13g2_nand2_1 _06626_ (.Y(_02151_),
    .A(net3203),
    .B(net1943));
 sg13g2_o21ai_1 _06627_ (.B1(_02151_),
    .Y(_01068_),
    .A1(net2521),
    .A2(net1943));
 sg13g2_nand2_1 _06628_ (.Y(_02152_),
    .A(net3188),
    .B(net1943));
 sg13g2_o21ai_1 _06629_ (.B1(_02152_),
    .Y(_01069_),
    .A1(net2514),
    .A2(net1943));
 sg13g2_nand2_1 _06630_ (.Y(_02153_),
    .A(net2959),
    .B(net1943));
 sg13g2_o21ai_1 _06631_ (.B1(_02153_),
    .Y(_01070_),
    .A1(net2509),
    .A2(net1943));
 sg13g2_nand2_1 _06632_ (.Y(_02154_),
    .A(net1635),
    .B(net1942));
 sg13g2_o21ai_1 _06633_ (.B1(_02154_),
    .Y(_01071_),
    .A1(net2505),
    .A2(net1942));
 sg13g2_nand2_1 _06634_ (.Y(_02155_),
    .A(net2798),
    .B(net1943));
 sg13g2_o21ai_1 _06635_ (.B1(_02155_),
    .Y(_01072_),
    .A1(net2501),
    .A2(net1943));
 sg13g2_nand2_1 _06636_ (.Y(_02156_),
    .A(net3199),
    .B(net1945));
 sg13g2_o21ai_1 _06637_ (.B1(_02156_),
    .Y(_01073_),
    .A1(net2493),
    .A2(net1945));
 sg13g2_nand2_1 _06638_ (.Y(_02157_),
    .A(net3289),
    .B(net1938));
 sg13g2_o21ai_1 _06639_ (.B1(_02157_),
    .Y(_01074_),
    .A1(net2489),
    .A2(net1941));
 sg13g2_nand2_1 _06640_ (.Y(_02158_),
    .A(net3091),
    .B(net1942));
 sg13g2_o21ai_1 _06641_ (.B1(_02158_),
    .Y(_01075_),
    .A1(net2483),
    .A2(net1942));
 sg13g2_nand2_1 _06642_ (.Y(_02159_),
    .A(net3129),
    .B(net1942));
 sg13g2_o21ai_1 _06643_ (.B1(_02159_),
    .Y(_01076_),
    .A1(net2477),
    .A2(net1942));
 sg13g2_nand2_1 _06644_ (.Y(_02160_),
    .A(net2676),
    .B(net1938));
 sg13g2_o21ai_1 _06645_ (.B1(_02160_),
    .Y(_01077_),
    .A1(net2472),
    .A2(net1938));
 sg13g2_nand2_1 _06646_ (.Y(_02161_),
    .A(net1715),
    .B(net1942));
 sg13g2_o21ai_1 _06647_ (.B1(_02161_),
    .Y(_01078_),
    .A1(net2466),
    .A2(net1942));
 sg13g2_nand2_1 _06648_ (.Y(_02162_),
    .A(net1432),
    .B(net1937));
 sg13g2_o21ai_1 _06649_ (.B1(_02162_),
    .Y(_01079_),
    .A1(net2460),
    .A2(net1937));
 sg13g2_nand2_1 _06650_ (.Y(_02163_),
    .A(net2935),
    .B(net1938));
 sg13g2_o21ai_1 _06651_ (.B1(_02163_),
    .Y(_01080_),
    .A1(net2458),
    .A2(net1938));
 sg13g2_nand2_1 _06652_ (.Y(_02164_),
    .A(net3324),
    .B(net1940));
 sg13g2_o21ai_1 _06653_ (.B1(_02164_),
    .Y(_01081_),
    .A1(net2451),
    .A2(net1941));
 sg13g2_nand2_1 _06654_ (.Y(_02165_),
    .A(net1664),
    .B(net1945));
 sg13g2_o21ai_1 _06655_ (.B1(_02165_),
    .Y(_01082_),
    .A1(net2447),
    .A2(net1945));
 sg13g2_nand2_1 _06656_ (.Y(_02166_),
    .A(net1499),
    .B(net1939));
 sg13g2_o21ai_1 _06657_ (.B1(_02166_),
    .Y(_01083_),
    .A1(net2442),
    .A2(net1939));
 sg13g2_nand2_1 _06658_ (.Y(_02167_),
    .A(net3204),
    .B(net1940));
 sg13g2_o21ai_1 _06659_ (.B1(_02167_),
    .Y(_01084_),
    .A1(net2438),
    .A2(net1940));
 sg13g2_nand2_1 _06660_ (.Y(_02168_),
    .A(net2827),
    .B(net1939));
 sg13g2_o21ai_1 _06661_ (.B1(_02168_),
    .Y(_01085_),
    .A1(net2431),
    .A2(net1939));
 sg13g2_nand2_1 _06662_ (.Y(_02169_),
    .A(net1677),
    .B(net1940));
 sg13g2_o21ai_1 _06663_ (.B1(_02169_),
    .Y(_01086_),
    .A1(net2424),
    .A2(net1940));
 sg13g2_nand2_1 _06664_ (.Y(_02170_),
    .A(net2815),
    .B(net1939));
 sg13g2_o21ai_1 _06665_ (.B1(_02170_),
    .Y(_01087_),
    .A1(net2420),
    .A2(net1939));
 sg13g2_nand2_1 _06666_ (.Y(_02171_),
    .A(net2902),
    .B(net1939));
 sg13g2_o21ai_1 _06667_ (.B1(_02171_),
    .Y(_01088_),
    .A1(net2416),
    .A2(net1939));
 sg13g2_nand2_1 _06668_ (.Y(_02172_),
    .A(net1466),
    .B(net1937));
 sg13g2_o21ai_1 _06669_ (.B1(_02172_),
    .Y(_01089_),
    .A1(net2411),
    .A2(net1937));
 sg13g2_nand2_1 _06670_ (.Y(_02173_),
    .A(net2691),
    .B(net1937));
 sg13g2_o21ai_1 _06671_ (.B1(_02173_),
    .Y(_01090_),
    .A1(net2405),
    .A2(net1937));
 sg13g2_nand2_1 _06672_ (.Y(_02174_),
    .A(net2889),
    .B(net1937));
 sg13g2_o21ai_1 _06673_ (.B1(_02174_),
    .Y(_01091_),
    .A1(net2400),
    .A2(net1937));
 sg13g2_nand2_2 _06674_ (.Y(_02175_),
    .A(_01678_),
    .B(_01716_));
 sg13g2_nand2_1 _06675_ (.Y(_02176_),
    .A(net2711),
    .B(net1927));
 sg13g2_o21ai_1 _06676_ (.B1(_02176_),
    .Y(_01092_),
    .A1(net2560),
    .A2(net1927));
 sg13g2_nand2_1 _06677_ (.Y(_02177_),
    .A(net1589),
    .B(net1929));
 sg13g2_o21ai_1 _06678_ (.B1(_02177_),
    .Y(_01093_),
    .A1(net2557),
    .A2(net1929));
 sg13g2_nand2_1 _06679_ (.Y(_02178_),
    .A(net3096),
    .B(net1934));
 sg13g2_o21ai_1 _06680_ (.B1(_02178_),
    .Y(_01094_),
    .A1(net2553),
    .A2(net1935));
 sg13g2_nand2_1 _06681_ (.Y(_02179_),
    .A(net2901),
    .B(net1935));
 sg13g2_o21ai_1 _06682_ (.B1(_02179_),
    .Y(_01095_),
    .A1(net2547),
    .A2(net1935));
 sg13g2_nand2_1 _06683_ (.Y(_02180_),
    .A(net2777),
    .B(net1934));
 sg13g2_o21ai_1 _06684_ (.B1(_02180_),
    .Y(_01096_),
    .A1(net2539),
    .A2(net1935));
 sg13g2_nand2_1 _06685_ (.Y(_02181_),
    .A(net3028),
    .B(net1935));
 sg13g2_o21ai_1 _06686_ (.B1(_02181_),
    .Y(_01097_),
    .A1(net2535),
    .A2(net1935));
 sg13g2_nand2_1 _06687_ (.Y(_02182_),
    .A(net1681),
    .B(net1936));
 sg13g2_o21ai_1 _06688_ (.B1(_02182_),
    .Y(_01098_),
    .A1(net2531),
    .A2(net1936));
 sg13g2_nand2_1 _06689_ (.Y(_02183_),
    .A(net2622),
    .B(net1935));
 sg13g2_o21ai_1 _06690_ (.B1(_02183_),
    .Y(_01099_),
    .A1(net2526),
    .A2(net1936));
 sg13g2_nand2_1 _06691_ (.Y(_02184_),
    .A(net2866),
    .B(net1933));
 sg13g2_o21ai_1 _06692_ (.B1(_02184_),
    .Y(_01100_),
    .A1(net2522),
    .A2(net1933));
 sg13g2_nand2_1 _06693_ (.Y(_02185_),
    .A(net1518),
    .B(net1933));
 sg13g2_o21ai_1 _06694_ (.B1(_02185_),
    .Y(_01101_),
    .A1(net2515),
    .A2(net1933));
 sg13g2_nand2_1 _06695_ (.Y(_02186_),
    .A(net3215),
    .B(net1932));
 sg13g2_o21ai_1 _06696_ (.B1(_02186_),
    .Y(_01102_),
    .A1(net2510),
    .A2(net1932));
 sg13g2_nand2_1 _06697_ (.Y(_02187_),
    .A(net3290),
    .B(net1932));
 sg13g2_o21ai_1 _06698_ (.B1(_02187_),
    .Y(_01103_),
    .A1(net2505),
    .A2(net1932));
 sg13g2_nand2_1 _06699_ (.Y(_02188_),
    .A(net2761),
    .B(net1933));
 sg13g2_o21ai_1 _06700_ (.B1(_02188_),
    .Y(_01104_),
    .A1(net2500),
    .A2(net1933));
 sg13g2_nand2_1 _06701_ (.Y(_02189_),
    .A(net2956),
    .B(net1934));
 sg13g2_o21ai_1 _06702_ (.B1(_02189_),
    .Y(_01105_),
    .A1(net2494),
    .A2(net1934));
 sg13g2_nand2_1 _06703_ (.Y(_02190_),
    .A(net1539),
    .B(net1931));
 sg13g2_o21ai_1 _06704_ (.B1(_02190_),
    .Y(_01106_),
    .A1(net2487),
    .A2(net1931));
 sg13g2_nand2_1 _06705_ (.Y(_02191_),
    .A(net1624),
    .B(net1928));
 sg13g2_o21ai_1 _06706_ (.B1(_02191_),
    .Y(_01107_),
    .A1(net2481),
    .A2(net1928));
 sg13g2_nand2_1 _06707_ (.Y(_02192_),
    .A(net2652),
    .B(net1932));
 sg13g2_o21ai_1 _06708_ (.B1(_02192_),
    .Y(_01108_),
    .A1(net2475),
    .A2(net1932));
 sg13g2_nand2_1 _06709_ (.Y(_02193_),
    .A(net1452),
    .B(net1928));
 sg13g2_o21ai_1 _06710_ (.B1(_02193_),
    .Y(_01109_),
    .A1(net2473),
    .A2(net1928));
 sg13g2_nand2_1 _06711_ (.Y(_02194_),
    .A(net1549),
    .B(net1932));
 sg13g2_o21ai_1 _06712_ (.B1(_02194_),
    .Y(_01110_),
    .A1(net2467),
    .A2(net1932));
 sg13g2_nand2_1 _06713_ (.Y(_02195_),
    .A(net3311),
    .B(net1926));
 sg13g2_o21ai_1 _06714_ (.B1(_02195_),
    .Y(_01111_),
    .A1(net2461),
    .A2(net1926));
 sg13g2_nand2_1 _06715_ (.Y(_02196_),
    .A(net1567),
    .B(net1928));
 sg13g2_o21ai_1 _06716_ (.B1(_02196_),
    .Y(_01112_),
    .A1(net2455),
    .A2(net1928));
 sg13g2_nand2_1 _06717_ (.Y(_02197_),
    .A(net3030),
    .B(net1930));
 sg13g2_o21ai_1 _06718_ (.B1(_02197_),
    .Y(_01113_),
    .A1(net2453),
    .A2(net1930));
 sg13g2_nand2_1 _06719_ (.Y(_02198_),
    .A(net2892),
    .B(net1934));
 sg13g2_o21ai_1 _06720_ (.B1(_02198_),
    .Y(_01114_),
    .A1(net2448),
    .A2(net1934));
 sg13g2_nand2_1 _06721_ (.Y(_02199_),
    .A(net3241),
    .B(net1927));
 sg13g2_o21ai_1 _06722_ (.B1(_02199_),
    .Y(_01115_),
    .A1(net2441),
    .A2(net1927));
 sg13g2_nand2_1 _06723_ (.Y(_02200_),
    .A(net3106),
    .B(net1934));
 sg13g2_o21ai_1 _06724_ (.B1(_02200_),
    .Y(_01116_),
    .A1(net2436),
    .A2(net1934));
 sg13g2_nand2_1 _06725_ (.Y(_02201_),
    .A(net3072),
    .B(net1930));
 sg13g2_o21ai_1 _06726_ (.B1(_02201_),
    .Y(_01117_),
    .A1(net2432),
    .A2(net1930));
 sg13g2_nand2_1 _06727_ (.Y(_02202_),
    .A(net2964),
    .B(net1929));
 sg13g2_o21ai_1 _06728_ (.B1(_02202_),
    .Y(_01118_),
    .A1(net2427),
    .A2(net1929));
 sg13g2_nand2_1 _06729_ (.Y(_02203_),
    .A(net2721),
    .B(net1929));
 sg13g2_o21ai_1 _06730_ (.B1(_02203_),
    .Y(_01119_),
    .A1(net2422),
    .A2(net1929));
 sg13g2_nand2_1 _06731_ (.Y(_02204_),
    .A(net2891),
    .B(net1929));
 sg13g2_o21ai_1 _06732_ (.B1(_02204_),
    .Y(_01120_),
    .A1(net2416),
    .A2(net1929));
 sg13g2_nand2_1 _06733_ (.Y(_02205_),
    .A(net1586),
    .B(net1926));
 sg13g2_o21ai_1 _06734_ (.B1(_02205_),
    .Y(_01121_),
    .A1(net2409),
    .A2(net1926));
 sg13g2_nand2_1 _06735_ (.Y(_02206_),
    .A(net1582),
    .B(net1926));
 sg13g2_o21ai_1 _06736_ (.B1(_02206_),
    .Y(_01122_),
    .A1(net2405),
    .A2(net1926));
 sg13g2_nand2_1 _06737_ (.Y(_02207_),
    .A(net3126),
    .B(net1926));
 sg13g2_o21ai_1 _06738_ (.B1(_02207_),
    .Y(_01123_),
    .A1(net2398),
    .A2(net1926));
 sg13g2_nand2_2 _06739_ (.Y(_02208_),
    .A(_01616_),
    .B(_01678_));
 sg13g2_nand2_1 _06740_ (.Y(_02209_),
    .A(net1630),
    .B(net1917));
 sg13g2_o21ai_1 _06741_ (.B1(_02209_),
    .Y(_01124_),
    .A1(net2564),
    .A2(net1917));
 sg13g2_nand2_1 _06742_ (.Y(_02210_),
    .A(net3060),
    .B(net1919));
 sg13g2_o21ai_1 _06743_ (.B1(_02210_),
    .Y(_01125_),
    .A1(net2559),
    .A2(net1919));
 sg13g2_nand2_1 _06744_ (.Y(_02211_),
    .A(net2981),
    .B(net1923));
 sg13g2_o21ai_1 _06745_ (.B1(_02211_),
    .Y(_01126_),
    .A1(net2553),
    .A2(net1924));
 sg13g2_nand2_1 _06746_ (.Y(_02212_),
    .A(net3083),
    .B(net1924));
 sg13g2_o21ai_1 _06747_ (.B1(_02212_),
    .Y(_01127_),
    .A1(net2546),
    .A2(net1924));
 sg13g2_nand2_1 _06748_ (.Y(_02213_),
    .A(net1639),
    .B(net1923));
 sg13g2_o21ai_1 _06749_ (.B1(_02213_),
    .Y(_01128_),
    .A1(net2538),
    .A2(net1924));
 sg13g2_nand2_1 _06750_ (.Y(_02214_),
    .A(net2861),
    .B(net1924));
 sg13g2_o21ai_1 _06751_ (.B1(_02214_),
    .Y(_01129_),
    .A1(net2535),
    .A2(net1924));
 sg13g2_nand2_1 _06752_ (.Y(_02215_),
    .A(net2605),
    .B(net1925));
 sg13g2_o21ai_1 _06753_ (.B1(_02215_),
    .Y(_01130_),
    .A1(net2530),
    .A2(net1925));
 sg13g2_nand2_1 _06754_ (.Y(_02216_),
    .A(net3075),
    .B(net1924));
 sg13g2_o21ai_1 _06755_ (.B1(_02216_),
    .Y(_01131_),
    .A1(net2526),
    .A2(net1925));
 sg13g2_nand2_1 _06756_ (.Y(_02217_),
    .A(net1495),
    .B(net1922));
 sg13g2_o21ai_1 _06757_ (.B1(_02217_),
    .Y(_01132_),
    .A1(net2521),
    .A2(net1922));
 sg13g2_nand2_1 _06758_ (.Y(_02218_),
    .A(net3222),
    .B(net1922));
 sg13g2_o21ai_1 _06759_ (.B1(_02218_),
    .Y(_01133_),
    .A1(net2515),
    .A2(net1922));
 sg13g2_nand2_1 _06760_ (.Y(_02219_),
    .A(net1733),
    .B(net1921));
 sg13g2_o21ai_1 _06761_ (.B1(_02219_),
    .Y(_01134_),
    .A1(net2510),
    .A2(net1921));
 sg13g2_nand2_1 _06762_ (.Y(_02220_),
    .A(net1483),
    .B(net1921));
 sg13g2_o21ai_1 _06763_ (.B1(_02220_),
    .Y(_01135_),
    .A1(net2505),
    .A2(net1921));
 sg13g2_nand2_1 _06764_ (.Y(_02221_),
    .A(net1680),
    .B(net1922));
 sg13g2_o21ai_1 _06765_ (.B1(_02221_),
    .Y(_01136_),
    .A1(net2500),
    .A2(net1922));
 sg13g2_nand2_1 _06766_ (.Y(_02222_),
    .A(net3150),
    .B(net1923));
 sg13g2_o21ai_1 _06767_ (.B1(_02222_),
    .Y(_01137_),
    .A1(net2494),
    .A2(net1923));
 sg13g2_nand2_1 _06768_ (.Y(_02223_),
    .A(net1534),
    .B(net1920));
 sg13g2_o21ai_1 _06769_ (.B1(_02223_),
    .Y(_01138_),
    .A1(net2490),
    .A2(net1920));
 sg13g2_nand2_1 _06770_ (.Y(_02224_),
    .A(net1672),
    .B(net1917));
 sg13g2_o21ai_1 _06771_ (.B1(_02224_),
    .Y(_01139_),
    .A1(net2481),
    .A2(net1917));
 sg13g2_nand2_1 _06772_ (.Y(_02225_),
    .A(net1665),
    .B(net1921));
 sg13g2_o21ai_1 _06773_ (.B1(_02225_),
    .Y(_01140_),
    .A1(net2477),
    .A2(net1921));
 sg13g2_nand2_1 _06774_ (.Y(_02226_),
    .A(net1729),
    .B(net1917));
 sg13g2_o21ai_1 _06775_ (.B1(_02226_),
    .Y(_01141_),
    .A1(net2474),
    .A2(net1917));
 sg13g2_nand2_1 _06776_ (.Y(_02227_),
    .A(net2983),
    .B(net1921));
 sg13g2_o21ai_1 _06777_ (.B1(_02227_),
    .Y(_01142_),
    .A1(net2467),
    .A2(net1921));
 sg13g2_nand2_1 _06778_ (.Y(_02228_),
    .A(net3212),
    .B(net1916));
 sg13g2_o21ai_1 _06779_ (.B1(_02228_),
    .Y(_01143_),
    .A1(net2461),
    .A2(net1916));
 sg13g2_nand2_1 _06780_ (.Y(_02229_),
    .A(net3074),
    .B(net1917));
 sg13g2_o21ai_1 _06781_ (.B1(_02229_),
    .Y(_01144_),
    .A1(net2456),
    .A2(net1920));
 sg13g2_nand2_1 _06782_ (.Y(_02230_),
    .A(net3259),
    .B(net1919));
 sg13g2_o21ai_1 _06783_ (.B1(_02230_),
    .Y(_01145_),
    .A1(net2454),
    .A2(net1919));
 sg13g2_nand2_1 _06784_ (.Y(_02231_),
    .A(net3024),
    .B(net1923));
 sg13g2_o21ai_1 _06785_ (.B1(_02231_),
    .Y(_01146_),
    .A1(net2448),
    .A2(net1923));
 sg13g2_nand2_1 _06786_ (.Y(_02232_),
    .A(net1694),
    .B(net1918));
 sg13g2_o21ai_1 _06787_ (.B1(_02232_),
    .Y(_01147_),
    .A1(net2441),
    .A2(net1918));
 sg13g2_nand2_1 _06788_ (.Y(_02233_),
    .A(net2940),
    .B(net1923));
 sg13g2_o21ai_1 _06789_ (.B1(_02233_),
    .Y(_01148_),
    .A1(net2437),
    .A2(net1923));
 sg13g2_nand2_1 _06790_ (.Y(_02234_),
    .A(net2752),
    .B(net1918));
 sg13g2_o21ai_1 _06791_ (.B1(_02234_),
    .Y(_01149_),
    .A1(net2432),
    .A2(net1918));
 sg13g2_nand2_1 _06792_ (.Y(_02235_),
    .A(net2937),
    .B(net1918));
 sg13g2_o21ai_1 _06793_ (.B1(_02235_),
    .Y(_01150_),
    .A1(net2427),
    .A2(net1918));
 sg13g2_nand2_1 _06794_ (.Y(_02236_),
    .A(net1563),
    .B(net1919));
 sg13g2_o21ai_1 _06795_ (.B1(_02236_),
    .Y(_01151_),
    .A1(net2422),
    .A2(net1919));
 sg13g2_nand2_1 _06796_ (.Y(_02237_),
    .A(net1704),
    .B(net1918));
 sg13g2_o21ai_1 _06797_ (.B1(_02237_),
    .Y(_01152_),
    .A1(net2417),
    .A2(net1918));
 sg13g2_nand2_1 _06798_ (.Y(_02238_),
    .A(net1438),
    .B(net1916));
 sg13g2_o21ai_1 _06799_ (.B1(_02238_),
    .Y(_01153_),
    .A1(net2411),
    .A2(net1916));
 sg13g2_nand2_1 _06800_ (.Y(_02239_),
    .A(net2684),
    .B(net1916));
 sg13g2_o21ai_1 _06801_ (.B1(_02239_),
    .Y(_01154_),
    .A1(net2405),
    .A2(net1916));
 sg13g2_nand2_1 _06802_ (.Y(_02240_),
    .A(net1668),
    .B(net1916));
 sg13g2_o21ai_1 _06803_ (.B1(_02240_),
    .Y(_01155_),
    .A1(net2400),
    .A2(net1916));
 sg13g2_nand2_1 _06804_ (.Y(_02241_),
    .A(_01547_),
    .B(_01825_));
 sg13g2_nand2_1 _06805_ (.Y(_02242_),
    .A(net3202),
    .B(net1906));
 sg13g2_o21ai_1 _06806_ (.B1(_02242_),
    .Y(_01156_),
    .A1(net2561),
    .A2(net1906));
 sg13g2_nand2_1 _06807_ (.Y(_02243_),
    .A(net2768),
    .B(net1907));
 sg13g2_o21ai_1 _06808_ (.B1(_02243_),
    .Y(_01157_),
    .A1(net2558),
    .A2(net1907));
 sg13g2_nand2_1 _06809_ (.Y(_02244_),
    .A(net3299),
    .B(net1914));
 sg13g2_o21ai_1 _06810_ (.B1(_02244_),
    .Y(_01158_),
    .A1(net2552),
    .A2(net1914));
 sg13g2_nand2_1 _06811_ (.Y(_02245_),
    .A(net2657),
    .B(net1915));
 sg13g2_o21ai_1 _06812_ (.B1(_02245_),
    .Y(_01159_),
    .A1(net2548),
    .A2(net1914));
 sg13g2_nand2_1 _06813_ (.Y(_02246_),
    .A(net2961),
    .B(net1913));
 sg13g2_o21ai_1 _06814_ (.B1(_02246_),
    .Y(_01160_),
    .A1(net2543),
    .A2(net1913));
 sg13g2_nand2_1 _06815_ (.Y(_02247_),
    .A(net3207),
    .B(net1913));
 sg13g2_o21ai_1 _06816_ (.B1(_02247_),
    .Y(_01161_),
    .A1(net2534),
    .A2(net1913));
 sg13g2_nand2_1 _06817_ (.Y(_02248_),
    .A(net2988),
    .B(net1913));
 sg13g2_o21ai_1 _06818_ (.B1(_02248_),
    .Y(_01162_),
    .A1(net2529),
    .A2(net1913));
 sg13g2_nand2_1 _06819_ (.Y(_02249_),
    .A(net3101),
    .B(net1913));
 sg13g2_o21ai_1 _06820_ (.B1(_02249_),
    .Y(_01163_),
    .A1(net2525),
    .A2(net1913));
 sg13g2_nand2_1 _06821_ (.Y(_02250_),
    .A(net3122),
    .B(net1911));
 sg13g2_o21ai_1 _06822_ (.B1(_02250_),
    .Y(_01164_),
    .A1(net2522),
    .A2(net1911));
 sg13g2_nand2_1 _06823_ (.Y(_02251_),
    .A(net1571),
    .B(net1910));
 sg13g2_o21ai_1 _06824_ (.B1(_02251_),
    .Y(_01165_),
    .A1(net2513),
    .A2(net1910));
 sg13g2_nand2_1 _06825_ (.Y(_02252_),
    .A(net3320),
    .B(net1910));
 sg13g2_o21ai_1 _06826_ (.B1(_02252_),
    .Y(_01166_),
    .A1(net2508),
    .A2(net1910));
 sg13g2_nand2_1 _06827_ (.Y(_02253_),
    .A(net2635),
    .B(net1910));
 sg13g2_o21ai_1 _06828_ (.B1(_02253_),
    .Y(_01167_),
    .A1(net2505),
    .A2(net1910));
 sg13g2_nand2_1 _06829_ (.Y(_02254_),
    .A(net1474),
    .B(net1910));
 sg13g2_o21ai_1 _06830_ (.B1(_02254_),
    .Y(_01168_),
    .A1(net2499),
    .A2(net1910));
 sg13g2_nand2_1 _06831_ (.Y(_02255_),
    .A(net3117),
    .B(net1911));
 sg13g2_o21ai_1 _06832_ (.B1(_02255_),
    .Y(_01169_),
    .A1(net2493),
    .A2(net1911));
 sg13g2_nand2_1 _06833_ (.Y(_02256_),
    .A(net3201),
    .B(net1906));
 sg13g2_o21ai_1 _06834_ (.B1(_02256_),
    .Y(_01170_),
    .A1(net2490),
    .A2(net1906));
 sg13g2_nand2_1 _06835_ (.Y(_02257_),
    .A(net3270),
    .B(net1912));
 sg13g2_o21ai_1 _06836_ (.B1(_02257_),
    .Y(_01171_),
    .A1(net2482),
    .A2(net1912));
 sg13g2_nand2_1 _06837_ (.Y(_02258_),
    .A(net3079),
    .B(net1912));
 sg13g2_o21ai_1 _06838_ (.B1(_02258_),
    .Y(_01172_),
    .A1(net2475),
    .A2(net1912));
 sg13g2_nand2_1 _06839_ (.Y(_02259_),
    .A(net1720),
    .B(net1906));
 sg13g2_o21ai_1 _06840_ (.B1(_02259_),
    .Y(_01173_),
    .A1(net2473),
    .A2(net1906));
 sg13g2_nand2_1 _06841_ (.Y(_02260_),
    .A(net1748),
    .B(net1912));
 sg13g2_o21ai_1 _06842_ (.B1(_02260_),
    .Y(_01174_),
    .A1(net2465),
    .A2(net1912));
 sg13g2_nand2_1 _06843_ (.Y(_02261_),
    .A(net1511),
    .B(net1909));
 sg13g2_o21ai_1 _06844_ (.B1(_02261_),
    .Y(_01175_),
    .A1(net2463),
    .A2(net1909));
 sg13g2_nand2_1 _06845_ (.Y(_02262_),
    .A(net3239),
    .B(net1906));
 sg13g2_o21ai_1 _06846_ (.B1(_02262_),
    .Y(_01176_),
    .A1(net2459),
    .A2(net1909));
 sg13g2_nand2_1 _06847_ (.Y(_02263_),
    .A(net1625),
    .B(net1908));
 sg13g2_o21ai_1 _06848_ (.B1(_02263_),
    .Y(_01177_),
    .A1(net2454),
    .A2(net1908));
 sg13g2_nand2_1 _06849_ (.Y(_02264_),
    .A(net3302),
    .B(net1914));
 sg13g2_o21ai_1 _06850_ (.B1(_02264_),
    .Y(_01178_),
    .A1(net2446),
    .A2(net1914));
 sg13g2_nand2_1 _06851_ (.Y(_02265_),
    .A(net3317),
    .B(net1905));
 sg13g2_o21ai_1 _06852_ (.B1(_02265_),
    .Y(_01179_),
    .A1(net2439),
    .A2(net1905));
 sg13g2_nand2_1 _06853_ (.Y(_02266_),
    .A(net1699),
    .B(net1914));
 sg13g2_o21ai_1 _06854_ (.B1(_02266_),
    .Y(_01180_),
    .A1(net2434),
    .A2(net1914));
 sg13g2_nand2_1 _06855_ (.Y(_02267_),
    .A(net2616),
    .B(net1907));
 sg13g2_o21ai_1 _06856_ (.B1(_02267_),
    .Y(_01181_),
    .A1(net2430),
    .A2(net1907));
 sg13g2_nand2_1 _06857_ (.Y(_02268_),
    .A(net2628),
    .B(net1908));
 sg13g2_o21ai_1 _06858_ (.B1(_02268_),
    .Y(_01182_),
    .A1(net2427),
    .A2(net1908));
 sg13g2_nand2_1 _06859_ (.Y(_02269_),
    .A(net3048),
    .B(net1907));
 sg13g2_o21ai_1 _06860_ (.B1(_02269_),
    .Y(_01183_),
    .A1(net2421),
    .A2(net1907));
 sg13g2_nand2_1 _06861_ (.Y(_02270_),
    .A(net2679),
    .B(net1907));
 sg13g2_o21ai_1 _06862_ (.B1(_02270_),
    .Y(_01184_),
    .A1(net2413),
    .A2(net1907));
 sg13g2_nand2_1 _06863_ (.Y(_02271_),
    .A(net1448),
    .B(net1905));
 sg13g2_o21ai_1 _06864_ (.B1(_02271_),
    .Y(_01185_),
    .A1(net2408),
    .A2(net1905));
 sg13g2_nand2_1 _06865_ (.Y(_02272_),
    .A(net2834),
    .B(net1905));
 sg13g2_o21ai_1 _06866_ (.B1(_02272_),
    .Y(_01186_),
    .A1(net2405),
    .A2(net1905));
 sg13g2_nand2_1 _06867_ (.Y(_02273_),
    .A(net1731),
    .B(net1905));
 sg13g2_o21ai_1 _06868_ (.B1(_02273_),
    .Y(_01187_),
    .A1(net2398),
    .A2(net1905));
 sg13g2_nand2_1 _06869_ (.Y(_02274_),
    .A(_01547_),
    .B(_01713_));
 sg13g2_nand2_1 _06870_ (.Y(_02275_),
    .A(net3021),
    .B(net1896));
 sg13g2_o21ai_1 _06871_ (.B1(_02275_),
    .Y(_01188_),
    .A1(net2564),
    .A2(net1895));
 sg13g2_nand2_1 _06872_ (.Y(_02276_),
    .A(net1570),
    .B(net1898));
 sg13g2_o21ai_1 _06873_ (.B1(_02276_),
    .Y(_01189_),
    .A1(net2556),
    .A2(net1898));
 sg13g2_nand2_1 _06874_ (.Y(_02277_),
    .A(net3019),
    .B(net1903));
 sg13g2_o21ai_1 _06875_ (.B1(_02277_),
    .Y(_01190_),
    .A1(net2550),
    .A2(net1903));
 sg13g2_nand2_1 _06876_ (.Y(_02278_),
    .A(net3206),
    .B(net1901));
 sg13g2_o21ai_1 _06877_ (.B1(_02278_),
    .Y(_01191_),
    .A1(net2544),
    .A2(net1901));
 sg13g2_nand2_1 _06878_ (.Y(_02279_),
    .A(net2888),
    .B(net1902));
 sg13g2_o21ai_1 _06879_ (.B1(_02279_),
    .Y(_01192_),
    .A1(net2540),
    .A2(net1902));
 sg13g2_nand2_1 _06880_ (.Y(_02280_),
    .A(net1591),
    .B(net1902));
 sg13g2_o21ai_1 _06881_ (.B1(_02280_),
    .Y(_01193_),
    .A1(net2533),
    .A2(net1902));
 sg13g2_nand2_1 _06882_ (.Y(_02281_),
    .A(net1506),
    .B(net1901));
 sg13g2_o21ai_1 _06883_ (.B1(_02281_),
    .Y(_01194_),
    .A1(net2528),
    .A2(net1901));
 sg13g2_nand2_1 _06884_ (.Y(_02282_),
    .A(net1525),
    .B(net1901));
 sg13g2_o21ai_1 _06885_ (.B1(_02282_),
    .Y(_01195_),
    .A1(net2523),
    .A2(net1901));
 sg13g2_nand2_1 _06886_ (.Y(_02283_),
    .A(net2775),
    .B(net1899));
 sg13g2_o21ai_1 _06887_ (.B1(_02283_),
    .Y(_01196_),
    .A1(net2518),
    .A2(net1899));
 sg13g2_nand2_1 _06888_ (.Y(_02284_),
    .A(net2716),
    .B(net1899));
 sg13g2_o21ai_1 _06889_ (.B1(_02284_),
    .Y(_01197_),
    .A1(net2512),
    .A2(net1899));
 sg13g2_nand2_1 _06890_ (.Y(_02285_),
    .A(net3279),
    .B(net1904));
 sg13g2_o21ai_1 _06891_ (.B1(_02285_),
    .Y(_01198_),
    .A1(net2507),
    .A2(net1900));
 sg13g2_nand2_1 _06892_ (.Y(_02286_),
    .A(net3174),
    .B(net1899));
 sg13g2_o21ai_1 _06893_ (.B1(_02286_),
    .Y(_01199_),
    .A1(net2503),
    .A2(net1899));
 sg13g2_nand2_1 _06894_ (.Y(_02287_),
    .A(net1670),
    .B(net1899));
 sg13g2_o21ai_1 _06895_ (.B1(_02287_),
    .Y(_01200_),
    .A1(net2496),
    .A2(net1899));
 sg13g2_nand2_1 _06896_ (.Y(_02288_),
    .A(net2911),
    .B(net1901));
 sg13g2_o21ai_1 _06897_ (.B1(_02288_),
    .Y(_01201_),
    .A1(net2494),
    .A2(net1901));
 sg13g2_nand2_1 _06898_ (.Y(_02289_),
    .A(net2695),
    .B(net1896));
 sg13g2_o21ai_1 _06899_ (.B1(_02289_),
    .Y(_01202_),
    .A1(net2488),
    .A2(net1896));
 sg13g2_nand2_1 _06900_ (.Y(_02290_),
    .A(net2734),
    .B(net1900));
 sg13g2_o21ai_1 _06901_ (.B1(_02290_),
    .Y(_01203_),
    .A1(net2484),
    .A2(net1900));
 sg13g2_nand2_1 _06902_ (.Y(_02291_),
    .A(net2806),
    .B(net1902));
 sg13g2_o21ai_1 _06903_ (.B1(_02291_),
    .Y(_01204_),
    .A1(net2478),
    .A2(net1902));
 sg13g2_nand2_1 _06904_ (.Y(_02292_),
    .A(net2989),
    .B(net1900));
 sg13g2_o21ai_1 _06905_ (.B1(_02292_),
    .Y(_01205_),
    .A1(net2473),
    .A2(net1900));
 sg13g2_nand2_1 _06906_ (.Y(_02293_),
    .A(net2760),
    .B(net1900));
 sg13g2_o21ai_1 _06907_ (.B1(_02293_),
    .Y(_01206_),
    .A1(net2465),
    .A2(net1900));
 sg13g2_nand2_1 _06908_ (.Y(_02294_),
    .A(net1580),
    .B(net1896));
 sg13g2_o21ai_1 _06909_ (.B1(_02294_),
    .Y(_01207_),
    .A1(net2462),
    .A2(net1896));
 sg13g2_nand2_1 _06910_ (.Y(_02295_),
    .A(net2905),
    .B(net1896));
 sg13g2_o21ai_1 _06911_ (.B1(_02295_),
    .Y(_01208_),
    .A1(net2455),
    .A2(net1896));
 sg13g2_nand2_1 _06912_ (.Y(_02296_),
    .A(net2802),
    .B(net1898));
 sg13g2_o21ai_1 _06913_ (.B1(_02296_),
    .Y(_01209_),
    .A1(net2450),
    .A2(net1898));
 sg13g2_nand2_1 _06914_ (.Y(_02297_),
    .A(net2604),
    .B(net1903));
 sg13g2_o21ai_1 _06915_ (.B1(_02297_),
    .Y(_01210_),
    .A1(net2446),
    .A2(net1903));
 sg13g2_nand2_1 _06916_ (.Y(_02298_),
    .A(net2883),
    .B(net1897));
 sg13g2_o21ai_1 _06917_ (.B1(_02298_),
    .Y(_01211_),
    .A1(net2439),
    .A2(net1895));
 sg13g2_nand2_1 _06918_ (.Y(_02299_),
    .A(net2787),
    .B(net1903));
 sg13g2_o21ai_1 _06919_ (.B1(_02299_),
    .Y(_01212_),
    .A1(net2434),
    .A2(net1903));
 sg13g2_nand2_1 _06920_ (.Y(_02300_),
    .A(net2875),
    .B(net1897));
 sg13g2_o21ai_1 _06921_ (.B1(_02300_),
    .Y(_01213_),
    .A1(net2428),
    .A2(net1897));
 sg13g2_nand2_1 _06922_ (.Y(_02301_),
    .A(net2943),
    .B(net1897));
 sg13g2_o21ai_1 _06923_ (.B1(_02301_),
    .Y(_01214_),
    .A1(net2423),
    .A2(net1898));
 sg13g2_nand2_1 _06924_ (.Y(_02302_),
    .A(net2688),
    .B(net1897));
 sg13g2_o21ai_1 _06925_ (.B1(_02302_),
    .Y(_01215_),
    .A1(net2419),
    .A2(net1897));
 sg13g2_nand2_1 _06926_ (.Y(_02303_),
    .A(net3183),
    .B(net1897));
 sg13g2_o21ai_1 _06927_ (.B1(_02303_),
    .Y(_01216_),
    .A1(net2415),
    .A2(net1897));
 sg13g2_nand2_1 _06928_ (.Y(_02304_),
    .A(net2925),
    .B(net1895));
 sg13g2_o21ai_1 _06929_ (.B1(_02304_),
    .Y(_01217_),
    .A1(net2411),
    .A2(net1895));
 sg13g2_nand2_1 _06930_ (.Y(_02305_),
    .A(net1531),
    .B(net1895));
 sg13g2_o21ai_1 _06931_ (.B1(_02305_),
    .Y(_01218_),
    .A1(net2403),
    .A2(net1895));
 sg13g2_nand2_1 _06932_ (.Y(_02306_),
    .A(net2975),
    .B(net1895));
 sg13g2_o21ai_1 _06933_ (.B1(_02306_),
    .Y(_01219_),
    .A1(net2399),
    .A2(net1895));
 sg13g2_nand2b_2 _06934_ (.Y(_02307_),
    .B(_01616_),
    .A_N(net2307));
 sg13g2_nand2_1 _06935_ (.Y(_02308_),
    .A(net2839),
    .B(net1885));
 sg13g2_o21ai_1 _06936_ (.B1(_02308_),
    .Y(_01220_),
    .A1(net2560),
    .A2(net1885));
 sg13g2_nand2_1 _06937_ (.Y(_02309_),
    .A(net1709),
    .B(net1894));
 sg13g2_o21ai_1 _06938_ (.B1(_02309_),
    .Y(_01221_),
    .A1(net2557),
    .A2(net1888));
 sg13g2_nand2_1 _06939_ (.Y(_02310_),
    .A(net2831),
    .B(net1893));
 sg13g2_o21ai_1 _06940_ (.B1(_02310_),
    .Y(_01222_),
    .A1(net2554),
    .A2(net1893));
 sg13g2_nand2_1 _06941_ (.Y(_02311_),
    .A(net2607),
    .B(net1892));
 sg13g2_o21ai_1 _06942_ (.B1(_02311_),
    .Y(_01223_),
    .A1(net2544),
    .A2(net1893));
 sg13g2_nand2_1 _06943_ (.Y(_02312_),
    .A(net1482),
    .B(net1892));
 sg13g2_o21ai_1 _06944_ (.B1(_02312_),
    .Y(_01224_),
    .A1(net2538),
    .A2(net1893));
 sg13g2_nand2_1 _06945_ (.Y(_02313_),
    .A(net2625),
    .B(net1893));
 sg13g2_o21ai_1 _06946_ (.B1(_02313_),
    .Y(_01225_),
    .A1(net2534),
    .A2(net1893));
 sg13g2_nand2_1 _06947_ (.Y(_02314_),
    .A(net1463),
    .B(net1892));
 sg13g2_o21ai_1 _06948_ (.B1(_02314_),
    .Y(_01226_),
    .A1(net2528),
    .A2(net1892));
 sg13g2_nand2_1 _06949_ (.Y(_02315_),
    .A(net2845),
    .B(net1892));
 sg13g2_o21ai_1 _06950_ (.B1(_02315_),
    .Y(_01227_),
    .A1(net2523),
    .A2(net1892));
 sg13g2_nand2_1 _06951_ (.Y(_02316_),
    .A(net1656),
    .B(net1889));
 sg13g2_o21ai_1 _06952_ (.B1(_02316_),
    .Y(_01228_),
    .A1(net2518),
    .A2(net1889));
 sg13g2_nand2_1 _06953_ (.Y(_02317_),
    .A(net1477),
    .B(net1889));
 sg13g2_o21ai_1 _06954_ (.B1(_02317_),
    .Y(_01229_),
    .A1(net2513),
    .A2(net1889));
 sg13g2_nand2_1 _06955_ (.Y(_02318_),
    .A(net1550),
    .B(net1890));
 sg13g2_o21ai_1 _06956_ (.B1(_02318_),
    .Y(_01230_),
    .A1(net2507),
    .A2(net1890));
 sg13g2_nand2_1 _06957_ (.Y(_02319_),
    .A(net3170),
    .B(net1889));
 sg13g2_o21ai_1 _06958_ (.B1(_02319_),
    .Y(_01231_),
    .A1(net2502),
    .A2(net1889));
 sg13g2_nand2_1 _06959_ (.Y(_02320_),
    .A(net2844),
    .B(net1889));
 sg13g2_o21ai_1 _06960_ (.B1(_02320_),
    .Y(_01232_),
    .A1(net2496),
    .A2(net1889));
 sg13g2_nand2_1 _06961_ (.Y(_02321_),
    .A(net2859),
    .B(net1890));
 sg13g2_o21ai_1 _06962_ (.B1(_02321_),
    .Y(_01233_),
    .A1(net2492),
    .A2(net1890));
 sg13g2_nand2_1 _06963_ (.Y(_02322_),
    .A(net3071),
    .B(net1886));
 sg13g2_o21ai_1 _06964_ (.B1(_02322_),
    .Y(_01234_),
    .A1(net2486),
    .A2(net1886));
 sg13g2_nand2_1 _06965_ (.Y(_02323_),
    .A(net3141),
    .B(net1891));
 sg13g2_o21ai_1 _06966_ (.B1(_02323_),
    .Y(_01235_),
    .A1(net2482),
    .A2(net1891));
 sg13g2_nand2_1 _06967_ (.Y(_02324_),
    .A(net2653),
    .B(net1892));
 sg13g2_o21ai_1 _06968_ (.B1(_02324_),
    .Y(_01236_),
    .A1(net2478),
    .A2(net1892));
 sg13g2_nand2_1 _06969_ (.Y(_02325_),
    .A(net1444),
    .B(net1891));
 sg13g2_o21ai_1 _06970_ (.B1(_02325_),
    .Y(_01237_),
    .A1(net2470),
    .A2(net1891));
 sg13g2_nand2_1 _06971_ (.Y(_02326_),
    .A(net2780),
    .B(net1891));
 sg13g2_o21ai_1 _06972_ (.B1(_02326_),
    .Y(_01238_),
    .A1(net2465),
    .A2(net1891));
 sg13g2_nand2_1 _06973_ (.Y(_02327_),
    .A(net1566),
    .B(net1886));
 sg13g2_o21ai_1 _06974_ (.B1(_02327_),
    .Y(_01239_),
    .A1(net2463),
    .A2(net1886));
 sg13g2_nand2_1 _06975_ (.Y(_02328_),
    .A(net2786),
    .B(net1886));
 sg13g2_o21ai_1 _06976_ (.B1(_02328_),
    .Y(_01240_),
    .A1(net2455),
    .A2(net1886));
 sg13g2_nand2_1 _06977_ (.Y(_02329_),
    .A(net1443),
    .B(net1887));
 sg13g2_o21ai_1 _06978_ (.B1(_02329_),
    .Y(_01241_),
    .A1(net2450),
    .A2(net1887));
 sg13g2_nand2_1 _06979_ (.Y(_02330_),
    .A(net2931),
    .B(net1894));
 sg13g2_o21ai_1 _06980_ (.B1(_02330_),
    .Y(_01242_),
    .A1(net2445),
    .A2(net1894));
 sg13g2_nand2_1 _06981_ (.Y(_02331_),
    .A(net1606),
    .B(net1886));
 sg13g2_o21ai_1 _06982_ (.B1(_02331_),
    .Y(_01243_),
    .A1(net2439),
    .A2(net1886));
 sg13g2_nand2_1 _06983_ (.Y(_02332_),
    .A(net1556),
    .B(net1894));
 sg13g2_o21ai_1 _06984_ (.B1(_02332_),
    .Y(_01244_),
    .A1(net2436),
    .A2(net1894));
 sg13g2_nand2_1 _06985_ (.Y(_02333_),
    .A(net2950),
    .B(net1887));
 sg13g2_o21ai_1 _06986_ (.B1(_02333_),
    .Y(_01245_),
    .A1(net2429),
    .A2(net1887));
 sg13g2_nand2_1 _06987_ (.Y(_02334_),
    .A(net3031),
    .B(net1888));
 sg13g2_o21ai_1 _06988_ (.B1(_02334_),
    .Y(_01246_),
    .A1(net2425),
    .A2(net1888));
 sg13g2_nand2_1 _06989_ (.Y(_02335_),
    .A(net2779),
    .B(net1887));
 sg13g2_o21ai_1 _06990_ (.B1(_02335_),
    .Y(_01247_),
    .A1(net2418),
    .A2(net1887));
 sg13g2_nand2_1 _06991_ (.Y(_02336_),
    .A(net2689),
    .B(net1887));
 sg13g2_o21ai_1 _06992_ (.B1(_02336_),
    .Y(_01248_),
    .A1(net2413),
    .A2(net1887));
 sg13g2_nand2_1 _06993_ (.Y(_02337_),
    .A(net2611),
    .B(net1885));
 sg13g2_o21ai_1 _06994_ (.B1(_02337_),
    .Y(_01249_),
    .A1(net2410),
    .A2(net1885));
 sg13g2_nand2_1 _06995_ (.Y(_02338_),
    .A(net1421),
    .B(net1885));
 sg13g2_o21ai_1 _06996_ (.B1(_02338_),
    .Y(_01250_),
    .A1(net2403),
    .A2(net1885));
 sg13g2_nand2_1 _06997_ (.Y(_02339_),
    .A(net1478),
    .B(net1885));
 sg13g2_o21ai_1 _06998_ (.B1(_02339_),
    .Y(_01251_),
    .A1(net2397),
    .A2(net1885));
 sg13g2_nand2b_2 _06999_ (.Y(_02340_),
    .B(_01535_),
    .A_N(_01538_));
 sg13g2_nor2_2 _07000_ (.A(net2325),
    .B(_02340_),
    .Y(_02341_));
 sg13g2_or2_1 _07001_ (.X(_02342_),
    .B(_02340_),
    .A(_01533_));
 sg13g2_nand2_2 _07002_ (.Y(_02343_),
    .A(_01547_),
    .B(_02341_));
 sg13g2_nand2_1 _07003_ (.Y(_02344_),
    .A(net3337),
    .B(net1877));
 sg13g2_o21ai_1 _07004_ (.B1(_02344_),
    .Y(_01252_),
    .A1(net2563),
    .A2(net1877));
 sg13g2_nand2_1 _07005_ (.Y(_02345_),
    .A(net3268),
    .B(net1879));
 sg13g2_o21ai_1 _07006_ (.B1(_02345_),
    .Y(_01253_),
    .A1(net2555),
    .A2(net1879));
 sg13g2_nand2_1 _07007_ (.Y(_02346_),
    .A(net1737),
    .B(net1883));
 sg13g2_o21ai_1 _07008_ (.B1(_02346_),
    .Y(_01254_),
    .A1(net2551),
    .A2(net1883));
 sg13g2_nand2_1 _07009_ (.Y(_02347_),
    .A(net2958),
    .B(net1882));
 sg13g2_o21ai_1 _07010_ (.B1(_02347_),
    .Y(_01255_),
    .A1(net2547),
    .A2(net1882));
 sg13g2_nand2_1 _07011_ (.Y(_02348_),
    .A(net1551),
    .B(net1882));
 sg13g2_o21ai_1 _07012_ (.B1(_02348_),
    .Y(_01256_),
    .A1(net2541),
    .A2(net1882));
 sg13g2_nand2_1 _07013_ (.Y(_02349_),
    .A(net2640),
    .B(net1882));
 sg13g2_o21ai_1 _07014_ (.B1(_02349_),
    .Y(_01257_),
    .A1(net2537),
    .A2(net1884));
 sg13g2_nand2_1 _07015_ (.Y(_02350_),
    .A(net3112),
    .B(net1884));
 sg13g2_o21ai_1 _07016_ (.B1(_02350_),
    .Y(_01258_),
    .A1(net2530),
    .A2(net1883));
 sg13g2_nand2_1 _07017_ (.Y(_02351_),
    .A(net1735),
    .B(net1882));
 sg13g2_o21ai_1 _07018_ (.B1(_02351_),
    .Y(_01259_),
    .A1(net2527),
    .A2(net1882));
 sg13g2_nand2_1 _07019_ (.Y(_02352_),
    .A(net2930),
    .B(net1882));
 sg13g2_o21ai_1 _07020_ (.B1(_02352_),
    .Y(_01260_),
    .A1(net2521),
    .A2(net1880));
 sg13g2_nand2_1 _07021_ (.Y(_02353_),
    .A(net3321),
    .B(net1881));
 sg13g2_o21ai_1 _07022_ (.B1(_02353_),
    .Y(_01261_),
    .A1(net2514),
    .A2(net1881));
 sg13g2_nand2_1 _07023_ (.Y(_02354_),
    .A(net1647),
    .B(net1881));
 sg13g2_o21ai_1 _07024_ (.B1(_02354_),
    .Y(_01262_),
    .A1(net2509),
    .A2(net1881));
 sg13g2_nand2_1 _07025_ (.Y(_02355_),
    .A(net1693),
    .B(net1880));
 sg13g2_o21ai_1 _07026_ (.B1(_02355_),
    .Y(_01263_),
    .A1(net2502),
    .A2(net1880));
 sg13g2_nand2_1 _07027_ (.Y(_02356_),
    .A(net2757),
    .B(net1881));
 sg13g2_o21ai_1 _07028_ (.B1(_02356_),
    .Y(_01264_),
    .A1(net2496),
    .A2(net1881));
 sg13g2_nand2_1 _07029_ (.Y(_02357_),
    .A(net2854),
    .B(net1880));
 sg13g2_o21ai_1 _07030_ (.B1(_02357_),
    .Y(_01265_),
    .A1(net2491),
    .A2(net1880));
 sg13g2_nand2_1 _07031_ (.Y(_02358_),
    .A(net3151),
    .B(net1875));
 sg13g2_o21ai_1 _07032_ (.B1(_02358_),
    .Y(_01266_),
    .A1(net2486),
    .A2(net1875));
 sg13g2_nand2_1 _07033_ (.Y(_02359_),
    .A(net2962),
    .B(net1880));
 sg13g2_o21ai_1 _07034_ (.B1(_02359_),
    .Y(_01267_),
    .A1(net2483),
    .A2(net1875));
 sg13g2_nand2_1 _07035_ (.Y(_02360_),
    .A(net2926),
    .B(net1883));
 sg13g2_o21ai_1 _07036_ (.B1(_02360_),
    .Y(_01268_),
    .A1(net2475),
    .A2(net1883));
 sg13g2_nand2_1 _07037_ (.Y(_02361_),
    .A(net2909),
    .B(net1875));
 sg13g2_o21ai_1 _07038_ (.B1(_02361_),
    .Y(_01269_),
    .A1(net2471),
    .A2(net1875));
 sg13g2_nand2_1 _07039_ (.Y(_02362_),
    .A(net3248),
    .B(net1880));
 sg13g2_o21ai_1 _07040_ (.B1(_02362_),
    .Y(_01270_),
    .A1(net2466),
    .A2(net1880));
 sg13g2_nand2_1 _07041_ (.Y(_02363_),
    .A(net2860),
    .B(net1876));
 sg13g2_o21ai_1 _07042_ (.B1(_02363_),
    .Y(_01271_),
    .A1(net2462),
    .A2(net1875));
 sg13g2_nand2_1 _07043_ (.Y(_02364_),
    .A(net1659),
    .B(net1875));
 sg13g2_o21ai_1 _07044_ (.B1(_02364_),
    .Y(_01272_),
    .A1(net2458),
    .A2(net1875));
 sg13g2_nand2_1 _07045_ (.Y(_02365_),
    .A(net2870),
    .B(net1879));
 sg13g2_o21ai_1 _07046_ (.B1(_02365_),
    .Y(_01273_),
    .A1(net2453),
    .A2(net1879));
 sg13g2_nand2_1 _07047_ (.Y(_02366_),
    .A(net1598),
    .B(net1883));
 sg13g2_o21ai_1 _07048_ (.B1(_02366_),
    .Y(_01274_),
    .A1(net2444),
    .A2(net1883));
 sg13g2_nand2_1 _07049_ (.Y(_02367_),
    .A(net1558),
    .B(net1877));
 sg13g2_o21ai_1 _07050_ (.B1(_02367_),
    .Y(_01275_),
    .A1(net2443),
    .A2(net1877));
 sg13g2_nand2_1 _07051_ (.Y(_02368_),
    .A(net2655),
    .B(net1879));
 sg13g2_o21ai_1 _07052_ (.B1(_02368_),
    .Y(_01276_),
    .A1(net2435),
    .A2(net1879));
 sg13g2_nand2_1 _07053_ (.Y(_02369_),
    .A(net1698),
    .B(net1878));
 sg13g2_o21ai_1 _07054_ (.B1(_02369_),
    .Y(_01277_),
    .A1(net2431),
    .A2(net1878));
 sg13g2_nand2_1 _07055_ (.Y(_02370_),
    .A(net2984),
    .B(net1877));
 sg13g2_o21ai_1 _07056_ (.B1(_02370_),
    .Y(_01278_),
    .A1(net2426),
    .A2(net1877));
 sg13g2_nand2_1 _07057_ (.Y(_02371_),
    .A(net1574),
    .B(net1878));
 sg13g2_o21ai_1 _07058_ (.B1(_02371_),
    .Y(_01279_),
    .A1(net2420),
    .A2(net1878));
 sg13g2_nand2_1 _07059_ (.Y(_02372_),
    .A(net3110),
    .B(net1877));
 sg13g2_o21ai_1 _07060_ (.B1(_02372_),
    .Y(_01280_),
    .A1(net2416),
    .A2(net1877));
 sg13g2_nand2_1 _07061_ (.Y(_02373_),
    .A(net3053),
    .B(net1876));
 sg13g2_o21ai_1 _07062_ (.B1(_02373_),
    .Y(_01281_),
    .A1(net2412),
    .A2(net1876));
 sg13g2_nand2_1 _07063_ (.Y(_02374_),
    .A(net3076),
    .B(net1876));
 sg13g2_o21ai_1 _07064_ (.B1(_02374_),
    .Y(_01282_),
    .A1(net2402),
    .A2(net1876));
 sg13g2_nand2_1 _07065_ (.Y(_02375_),
    .A(net3029),
    .B(net1876));
 sg13g2_o21ai_1 _07066_ (.B1(_02375_),
    .Y(_01283_),
    .A1(net2399),
    .A2(net1876));
 sg13g2_nand2_1 _07067_ (.Y(_02376_),
    .A(_01616_),
    .B(_01713_));
 sg13g2_nand2_1 _07068_ (.Y(_02377_),
    .A(net2829),
    .B(net1865));
 sg13g2_o21ai_1 _07069_ (.B1(_02377_),
    .Y(_01284_),
    .A1(net2564),
    .A2(net1865));
 sg13g2_nand2_1 _07070_ (.Y(_02378_),
    .A(net2800),
    .B(net1866));
 sg13g2_o21ai_1 _07071_ (.B1(_02378_),
    .Y(_01285_),
    .A1(net2559),
    .A2(net1867));
 sg13g2_nand2_1 _07072_ (.Y(_02379_),
    .A(net3011),
    .B(net1873));
 sg13g2_o21ai_1 _07073_ (.B1(_02379_),
    .Y(_01286_),
    .A1(net2550),
    .A2(net1873));
 sg13g2_nand2_1 _07074_ (.Y(_02380_),
    .A(net1561),
    .B(net1871));
 sg13g2_o21ai_1 _07075_ (.B1(_02380_),
    .Y(_01287_),
    .A1(net2544),
    .A2(net1871));
 sg13g2_nand2_1 _07076_ (.Y(_02381_),
    .A(net1718),
    .B(net1872));
 sg13g2_o21ai_1 _07077_ (.B1(_02381_),
    .Y(_01288_),
    .A1(net2540),
    .A2(net1872));
 sg13g2_nand2_1 _07078_ (.Y(_02382_),
    .A(net1649),
    .B(net1872));
 sg13g2_o21ai_1 _07079_ (.B1(_02382_),
    .Y(_01289_),
    .A1(net2533),
    .A2(net1872));
 sg13g2_nand2_1 _07080_ (.Y(_02383_),
    .A(net1684),
    .B(net1871));
 sg13g2_o21ai_1 _07081_ (.B1(_02383_),
    .Y(_01290_),
    .A1(net2528),
    .A2(net1871));
 sg13g2_nand2_1 _07082_ (.Y(_02384_),
    .A(net2867),
    .B(net1871));
 sg13g2_o21ai_1 _07083_ (.B1(_02384_),
    .Y(_01291_),
    .A1(net2523),
    .A2(net1871));
 sg13g2_nand2_1 _07084_ (.Y(_02385_),
    .A(net2794),
    .B(net1869));
 sg13g2_o21ai_1 _07085_ (.B1(_02385_),
    .Y(_01292_),
    .A1(net2518),
    .A2(net1869));
 sg13g2_nand2_1 _07086_ (.Y(_02386_),
    .A(net2998),
    .B(net1869));
 sg13g2_o21ai_1 _07087_ (.B1(_02386_),
    .Y(_01293_),
    .A1(net2512),
    .A2(net1869));
 sg13g2_nand2_1 _07088_ (.Y(_02387_),
    .A(net3388),
    .B(net1874));
 sg13g2_o21ai_1 _07089_ (.B1(_02387_),
    .Y(_01294_),
    .A1(net2507),
    .A2(net1870));
 sg13g2_nand2_1 _07090_ (.Y(_02388_),
    .A(net1486),
    .B(net1869));
 sg13g2_o21ai_1 _07091_ (.B1(_02388_),
    .Y(_01295_),
    .A1(net2503),
    .A2(net1869));
 sg13g2_nand2_1 _07092_ (.Y(_02389_),
    .A(net1420),
    .B(net1869));
 sg13g2_o21ai_1 _07093_ (.B1(_02389_),
    .Y(_01296_),
    .A1(net2496),
    .A2(net1869));
 sg13g2_nand2_1 _07094_ (.Y(_02390_),
    .A(net3119),
    .B(net1871));
 sg13g2_o21ai_1 _07095_ (.B1(_02390_),
    .Y(_01297_),
    .A1(net2494),
    .A2(net1871));
 sg13g2_nand2_1 _07096_ (.Y(_02391_),
    .A(net1456),
    .B(net1865));
 sg13g2_o21ai_1 _07097_ (.B1(_02391_),
    .Y(_01298_),
    .A1(net2488),
    .A2(net1868));
 sg13g2_nand2_1 _07098_ (.Y(_02392_),
    .A(net3171),
    .B(net1870));
 sg13g2_o21ai_1 _07099_ (.B1(_02392_),
    .Y(_01299_),
    .A1(net2484),
    .A2(net1870));
 sg13g2_nand2_1 _07100_ (.Y(_02393_),
    .A(net2828),
    .B(net1872));
 sg13g2_o21ai_1 _07101_ (.B1(_02393_),
    .Y(_01300_),
    .A1(net2479),
    .A2(net1872));
 sg13g2_nand2_1 _07102_ (.Y(_02394_),
    .A(net2970),
    .B(net1870));
 sg13g2_o21ai_1 _07103_ (.B1(_02394_),
    .Y(_01301_),
    .A1(net2473),
    .A2(net1870));
 sg13g2_nand2_1 _07104_ (.Y(_02395_),
    .A(net2835),
    .B(net1870));
 sg13g2_o21ai_1 _07105_ (.B1(_02395_),
    .Y(_01302_),
    .A1(net2467),
    .A2(net1870));
 sg13g2_nand2_1 _07106_ (.Y(_02396_),
    .A(net2978),
    .B(net1865));
 sg13g2_o21ai_1 _07107_ (.B1(_02396_),
    .Y(_01303_),
    .A1(net2462),
    .A2(net1865));
 sg13g2_nand2_1 _07108_ (.Y(_02397_),
    .A(net1602),
    .B(net1865));
 sg13g2_o21ai_1 _07109_ (.B1(_02397_),
    .Y(_01304_),
    .A1(net2457),
    .A2(net1865));
 sg13g2_nand2_1 _07110_ (.Y(_02398_),
    .A(net3194),
    .B(net1867));
 sg13g2_o21ai_1 _07111_ (.B1(_02398_),
    .Y(_01305_),
    .A1(net2453),
    .A2(net1867));
 sg13g2_nand2_1 _07112_ (.Y(_02399_),
    .A(net3219),
    .B(net1873));
 sg13g2_o21ai_1 _07113_ (.B1(_02399_),
    .Y(_01306_),
    .A1(net2446),
    .A2(net1873));
 sg13g2_nand2_1 _07114_ (.Y(_02400_),
    .A(net3224),
    .B(net1864));
 sg13g2_o21ai_1 _07115_ (.B1(_02400_),
    .Y(_01307_),
    .A1(net2439),
    .A2(net1864));
 sg13g2_nand2_1 _07116_ (.Y(_02401_),
    .A(net2879),
    .B(net1873));
 sg13g2_o21ai_1 _07117_ (.B1(_02401_),
    .Y(_01308_),
    .A1(net2434),
    .A2(net1873));
 sg13g2_nand2_1 _07118_ (.Y(_02402_),
    .A(net1425),
    .B(net1866));
 sg13g2_o21ai_1 _07119_ (.B1(_02402_),
    .Y(_01309_),
    .A1(net2428),
    .A2(net1866));
 sg13g2_nand2_1 _07120_ (.Y(_02403_),
    .A(net1459),
    .B(net1867));
 sg13g2_o21ai_1 _07121_ (.B1(_02403_),
    .Y(_01310_),
    .A1(net2423),
    .A2(net1866));
 sg13g2_nand2_1 _07122_ (.Y(_02404_),
    .A(net3228),
    .B(net1866));
 sg13g2_o21ai_1 _07123_ (.B1(_02404_),
    .Y(_01311_),
    .A1(net2419),
    .A2(net1866));
 sg13g2_nand2_1 _07124_ (.Y(_02405_),
    .A(net2920),
    .B(net1866));
 sg13g2_o21ai_1 _07125_ (.B1(_02405_),
    .Y(_01312_),
    .A1(net2415),
    .A2(net1866));
 sg13g2_nand2_1 _07126_ (.Y(_02406_),
    .A(net1455),
    .B(net1864));
 sg13g2_o21ai_1 _07127_ (.B1(_02406_),
    .Y(_01313_),
    .A1(net2411),
    .A2(net1864));
 sg13g2_nand2_1 _07128_ (.Y(_02407_),
    .A(net2765),
    .B(net1864));
 sg13g2_o21ai_1 _07129_ (.B1(_02407_),
    .Y(_01314_),
    .A1(net2403),
    .A2(net1864));
 sg13g2_nand2_1 _07130_ (.Y(_02408_),
    .A(net1473),
    .B(net1864));
 sg13g2_o21ai_1 _07131_ (.B1(_02408_),
    .Y(_01315_),
    .A1(net2399),
    .A2(net1864));
 sg13g2_nand2_2 _07132_ (.Y(_02409_),
    .A(_01616_),
    .B(_02341_));
 sg13g2_nand2_1 _07133_ (.Y(_02410_),
    .A(net3251),
    .B(net1856));
 sg13g2_o21ai_1 _07134_ (.B1(_02410_),
    .Y(_01316_),
    .A1(net2563),
    .A2(net1856));
 sg13g2_nand2_1 _07135_ (.Y(_02411_),
    .A(net2710),
    .B(net1858));
 sg13g2_o21ai_1 _07136_ (.B1(_02411_),
    .Y(_01317_),
    .A1(net2555),
    .A2(net1858));
 sg13g2_nand2_1 _07137_ (.Y(_02412_),
    .A(net2776),
    .B(net1862));
 sg13g2_o21ai_1 _07138_ (.B1(_02412_),
    .Y(_01318_),
    .A1(net2551),
    .A2(net1862));
 sg13g2_nand2_1 _07139_ (.Y(_02413_),
    .A(net3243),
    .B(net1861));
 sg13g2_o21ai_1 _07140_ (.B1(_02413_),
    .Y(_01319_),
    .A1(net2547),
    .A2(net1861));
 sg13g2_nand2_1 _07141_ (.Y(_02414_),
    .A(net2969),
    .B(net1861));
 sg13g2_o21ai_1 _07142_ (.B1(_02414_),
    .Y(_01320_),
    .A1(net2541),
    .A2(net1861));
 sg13g2_nand2_1 _07143_ (.Y(_02415_),
    .A(net1690),
    .B(net1861));
 sg13g2_o21ai_1 _07144_ (.B1(_02415_),
    .Y(_01321_),
    .A1(net2537),
    .A2(net1863));
 sg13g2_nand2_1 _07145_ (.Y(_02416_),
    .A(net2697),
    .B(net1863));
 sg13g2_o21ai_1 _07146_ (.B1(_02416_),
    .Y(_01322_),
    .A1(net2530),
    .A2(net1862));
 sg13g2_nand2_1 _07147_ (.Y(_02417_),
    .A(net2885),
    .B(net1861));
 sg13g2_o21ai_1 _07148_ (.B1(_02417_),
    .Y(_01323_),
    .A1(net2527),
    .A2(net1861));
 sg13g2_nand2_1 _07149_ (.Y(_02418_),
    .A(net1746),
    .B(net1861));
 sg13g2_o21ai_1 _07150_ (.B1(_02418_),
    .Y(_01324_),
    .A1(net2521),
    .A2(net1859));
 sg13g2_nand2_1 _07151_ (.Y(_02419_),
    .A(net1540),
    .B(net1860));
 sg13g2_o21ai_1 _07152_ (.B1(_02419_),
    .Y(_01325_),
    .A1(net2514),
    .A2(net1860));
 sg13g2_nand2_1 _07153_ (.Y(_02420_),
    .A(net2896),
    .B(net1860));
 sg13g2_o21ai_1 _07154_ (.B1(_02420_),
    .Y(_01326_),
    .A1(net2509),
    .A2(net1860));
 sg13g2_nand2_1 _07155_ (.Y(_02421_),
    .A(net2947),
    .B(net1859));
 sg13g2_o21ai_1 _07156_ (.B1(_02421_),
    .Y(_01327_),
    .A1(net2502),
    .A2(net1859));
 sg13g2_nand2_1 _07157_ (.Y(_02422_),
    .A(net2946),
    .B(net1860));
 sg13g2_o21ai_1 _07158_ (.B1(_02422_),
    .Y(_01328_),
    .A1(net2496),
    .A2(net1860));
 sg13g2_nand2_1 _07159_ (.Y(_02423_),
    .A(net1481),
    .B(net1859));
 sg13g2_o21ai_1 _07160_ (.B1(_02423_),
    .Y(_01329_),
    .A1(net2491),
    .A2(net1859));
 sg13g2_nand2_1 _07161_ (.Y(_02424_),
    .A(net3046),
    .B(net1854));
 sg13g2_o21ai_1 _07162_ (.B1(_02424_),
    .Y(_01330_),
    .A1(net2486),
    .A2(net1854));
 sg13g2_nand2_1 _07163_ (.Y(_02425_),
    .A(net1530),
    .B(net1859));
 sg13g2_o21ai_1 _07164_ (.B1(_02425_),
    .Y(_01331_),
    .A1(net2483),
    .A2(net1854));
 sg13g2_nand2_1 _07165_ (.Y(_02426_),
    .A(net2632),
    .B(net1862));
 sg13g2_o21ai_1 _07166_ (.B1(_02426_),
    .Y(_01332_),
    .A1(net2476),
    .A2(net1862));
 sg13g2_nand2_1 _07167_ (.Y(_02427_),
    .A(net3002),
    .B(net1854));
 sg13g2_o21ai_1 _07168_ (.B1(_02427_),
    .Y(_00072_),
    .A1(net2471),
    .A2(net1854));
 sg13g2_nand2_1 _07169_ (.Y(_02428_),
    .A(net1514),
    .B(net1859));
 sg13g2_o21ai_1 _07170_ (.B1(_02428_),
    .Y(_00073_),
    .A1(net2466),
    .A2(net1859));
 sg13g2_nand2_1 _07171_ (.Y(_02429_),
    .A(net3009),
    .B(net1855));
 sg13g2_o21ai_1 _07172_ (.B1(_02429_),
    .Y(_00074_),
    .A1(net2462),
    .A2(net1854));
 sg13g2_nand2_1 _07173_ (.Y(_02430_),
    .A(net2813),
    .B(net1854));
 sg13g2_o21ai_1 _07174_ (.B1(_02430_),
    .Y(_00075_),
    .A1(net2458),
    .A2(net1854));
 sg13g2_nand2_1 _07175_ (.Y(_02431_),
    .A(net2769),
    .B(net1858));
 sg13g2_o21ai_1 _07176_ (.B1(_02431_),
    .Y(_00076_),
    .A1(net2453),
    .A2(net1858));
 sg13g2_nand2_1 _07177_ (.Y(_02432_),
    .A(net2972),
    .B(net1862));
 sg13g2_o21ai_1 _07178_ (.B1(_02432_),
    .Y(_00077_),
    .A1(net2444),
    .A2(net1862));
 sg13g2_nand2_1 _07179_ (.Y(_02433_),
    .A(net2921),
    .B(net1856));
 sg13g2_o21ai_1 _07180_ (.B1(_02433_),
    .Y(_00078_),
    .A1(net2443),
    .A2(net1856));
 sg13g2_nand2_1 _07181_ (.Y(_02434_),
    .A(net2656),
    .B(net1858));
 sg13g2_o21ai_1 _07182_ (.B1(_02434_),
    .Y(_00079_),
    .A1(net2435),
    .A2(net1858));
 sg13g2_nand2_1 _07183_ (.Y(_02435_),
    .A(net1678),
    .B(net1857));
 sg13g2_o21ai_1 _07184_ (.B1(_02435_),
    .Y(_00080_),
    .A1(net2431),
    .A2(net1857));
 sg13g2_nand2_1 _07185_ (.Y(_02436_),
    .A(net1520),
    .B(net1856));
 sg13g2_o21ai_1 _07186_ (.B1(_02436_),
    .Y(_00081_),
    .A1(net2426),
    .A2(net1856));
 sg13g2_nand2_1 _07187_ (.Y(_02437_),
    .A(net1738),
    .B(net1857));
 sg13g2_o21ai_1 _07188_ (.B1(_02437_),
    .Y(_00082_),
    .A1(net2420),
    .A2(net1857));
 sg13g2_nand2_1 _07189_ (.Y(_02438_),
    .A(net3077),
    .B(net1856));
 sg13g2_o21ai_1 _07190_ (.B1(_02438_),
    .Y(_00083_),
    .A1(net2416),
    .A2(net1856));
 sg13g2_nand2_1 _07191_ (.Y(_02439_),
    .A(net2887),
    .B(net1855));
 sg13g2_o21ai_1 _07192_ (.B1(_02439_),
    .Y(_00084_),
    .A1(net2412),
    .A2(net1855));
 sg13g2_nand2_1 _07193_ (.Y(_02440_),
    .A(net1553),
    .B(net1855));
 sg13g2_o21ai_1 _07194_ (.B1(_02440_),
    .Y(_00085_),
    .A1(net2402),
    .A2(net1855));
 sg13g2_nand2_1 _07195_ (.Y(_02441_),
    .A(net1617),
    .B(net1855));
 sg13g2_o21ai_1 _07196_ (.B1(_02441_),
    .Y(_00086_),
    .A1(net2399),
    .A2(net1855));
 sg13g2_nand2_1 _07197_ (.Y(_02442_),
    .A(_01716_),
    .B(_02341_));
 sg13g2_nand2_1 _07198_ (.Y(_02443_),
    .A(net2807),
    .B(net1844));
 sg13g2_o21ai_1 _07199_ (.B1(_02443_),
    .Y(_00087_),
    .A1(net2563),
    .A2(net1844));
 sg13g2_nand2_1 _07200_ (.Y(_02444_),
    .A(net3128),
    .B(net1846));
 sg13g2_o21ai_1 _07201_ (.B1(_02444_),
    .Y(_00088_),
    .A1(net2556),
    .A2(net1846));
 sg13g2_nand2_1 _07202_ (.Y(_02445_),
    .A(net2917),
    .B(net1852));
 sg13g2_o21ai_1 _07203_ (.B1(_02445_),
    .Y(_00089_),
    .A1(net2551),
    .A2(net1852));
 sg13g2_nand2_1 _07204_ (.Y(_02446_),
    .A(net3264),
    .B(net1850));
 sg13g2_o21ai_1 _07205_ (.B1(_02446_),
    .Y(_00090_),
    .A1(net2548),
    .A2(net1850));
 sg13g2_nand2_1 _07206_ (.Y(_02447_),
    .A(net2772),
    .B(net1850));
 sg13g2_o21ai_1 _07207_ (.B1(_02447_),
    .Y(_00091_),
    .A1(net2541),
    .A2(net1850));
 sg13g2_nand2_1 _07208_ (.Y(_02448_),
    .A(net2713),
    .B(net1851));
 sg13g2_o21ai_1 _07209_ (.B1(_02448_),
    .Y(_00092_),
    .A1(net2537),
    .A2(net1851));
 sg13g2_nand2_1 _07210_ (.Y(_02449_),
    .A(net2890),
    .B(net1851));
 sg13g2_o21ai_1 _07211_ (.B1(_02449_),
    .Y(_00093_),
    .A1(net2531),
    .A2(net1851));
 sg13g2_nand2_1 _07212_ (.Y(_02450_),
    .A(net1562),
    .B(net1850));
 sg13g2_o21ai_1 _07213_ (.B1(_02450_),
    .Y(_00094_),
    .A1(net2527),
    .A2(net1850));
 sg13g2_nand2_1 _07214_ (.Y(_02451_),
    .A(net1657),
    .B(net1850));
 sg13g2_o21ai_1 _07215_ (.B1(_02451_),
    .Y(_00095_),
    .A1(net2520),
    .A2(net1850));
 sg13g2_nand2_1 _07216_ (.Y(_02452_),
    .A(net2621),
    .B(net1849));
 sg13g2_o21ai_1 _07217_ (.B1(_02452_),
    .Y(_00096_),
    .A1(net2514),
    .A2(net1849));
 sg13g2_nand2_1 _07218_ (.Y(_02453_),
    .A(net1687),
    .B(net1849));
 sg13g2_o21ai_1 _07219_ (.B1(_02453_),
    .Y(_00097_),
    .A1(net2509),
    .A2(net1849));
 sg13g2_nand2_1 _07220_ (.Y(_02454_),
    .A(net2948),
    .B(net1849));
 sg13g2_o21ai_1 _07221_ (.B1(_02454_),
    .Y(_00098_),
    .A1(net2502),
    .A2(net1848));
 sg13g2_nand2_1 _07222_ (.Y(_02455_),
    .A(net3008),
    .B(net1849));
 sg13g2_o21ai_1 _07223_ (.B1(_02455_),
    .Y(_00099_),
    .A1(net2501),
    .A2(net1849));
 sg13g2_nand2_1 _07224_ (.Y(_02456_),
    .A(net1701),
    .B(net1848));
 sg13g2_o21ai_1 _07225_ (.B1(_02456_),
    .Y(_00100_),
    .A1(net2491),
    .A2(net1848));
 sg13g2_nand2_1 _07226_ (.Y(_02457_),
    .A(net3269),
    .B(net1847));
 sg13g2_o21ai_1 _07227_ (.B1(_02457_),
    .Y(_00101_),
    .A1(net2486),
    .A2(net1847));
 sg13g2_nand2_1 _07228_ (.Y(_02458_),
    .A(net3307),
    .B(net1848));
 sg13g2_o21ai_1 _07229_ (.B1(_02458_),
    .Y(_00102_),
    .A1(net2483),
    .A2(net1848));
 sg13g2_nand2_1 _07230_ (.Y(_02459_),
    .A(net3218),
    .B(net1852));
 sg13g2_o21ai_1 _07231_ (.B1(_02459_),
    .Y(_00103_),
    .A1(net2476),
    .A2(net1852));
 sg13g2_nand2_1 _07232_ (.Y(_02460_),
    .A(net2771),
    .B(net1848));
 sg13g2_o21ai_1 _07233_ (.B1(_02460_),
    .Y(_00104_),
    .A1(net2471),
    .A2(net1843));
 sg13g2_nand2_1 _07234_ (.Y(_02461_),
    .A(net3138),
    .B(net1848));
 sg13g2_o21ai_1 _07235_ (.B1(_02461_),
    .Y(_00105_),
    .A1(net2468),
    .A2(net1848));
 sg13g2_nand2_1 _07236_ (.Y(_02462_),
    .A(net1524),
    .B(net1847));
 sg13g2_o21ai_1 _07237_ (.B1(_02462_),
    .Y(_00106_),
    .A1(net2462),
    .A2(net1843));
 sg13g2_nand2_1 _07238_ (.Y(_02463_),
    .A(net3231),
    .B(net1845));
 sg13g2_o21ai_1 _07239_ (.B1(_02463_),
    .Y(_00107_),
    .A1(net2458),
    .A2(net1845));
 sg13g2_nand2_1 _07240_ (.Y(_02464_),
    .A(net2797),
    .B(net1845));
 sg13g2_o21ai_1 _07241_ (.B1(_02464_),
    .Y(_00108_),
    .A1(net2453),
    .A2(net1845));
 sg13g2_nand2_1 _07242_ (.Y(_02465_),
    .A(net3260),
    .B(net1852));
 sg13g2_o21ai_1 _07243_ (.B1(_02465_),
    .Y(_00109_),
    .A1(net2444),
    .A2(net1852));
 sg13g2_nand2_1 _07244_ (.Y(_02466_),
    .A(net2630),
    .B(net1845));
 sg13g2_o21ai_1 _07245_ (.B1(_02466_),
    .Y(_00110_),
    .A1(net2443),
    .A2(net1845));
 sg13g2_nand2_1 _07246_ (.Y(_02467_),
    .A(net2755),
    .B(net1845));
 sg13g2_o21ai_1 _07247_ (.B1(_02467_),
    .Y(_00111_),
    .A1(net2435),
    .A2(net1845));
 sg13g2_nand2_1 _07248_ (.Y(_02468_),
    .A(net2743),
    .B(net1846));
 sg13g2_o21ai_1 _07249_ (.B1(_02468_),
    .Y(_00112_),
    .A1(net2432),
    .A2(net1846));
 sg13g2_nand2_1 _07250_ (.Y(_02469_),
    .A(net1584),
    .B(net1844));
 sg13g2_o21ai_1 _07251_ (.B1(_02469_),
    .Y(_00113_),
    .A1(net2425),
    .A2(net1844));
 sg13g2_nand2_1 _07252_ (.Y(_02470_),
    .A(net2764),
    .B(net1844));
 sg13g2_o21ai_1 _07253_ (.B1(_02470_),
    .Y(_00114_),
    .A1(net2418),
    .A2(net1844));
 sg13g2_nand2_1 _07254_ (.Y(_02471_),
    .A(net1609),
    .B(net1844));
 sg13g2_o21ai_1 _07255_ (.B1(_02471_),
    .Y(_00115_),
    .A1(net2415),
    .A2(net1844));
 sg13g2_nand2_1 _07256_ (.Y(_02472_),
    .A(net2748),
    .B(net1843));
 sg13g2_o21ai_1 _07257_ (.B1(_02472_),
    .Y(_00116_),
    .A1(net2410),
    .A2(net1843));
 sg13g2_nand2_1 _07258_ (.Y(_02473_),
    .A(net3088),
    .B(net1843));
 sg13g2_o21ai_1 _07259_ (.B1(_02473_),
    .Y(_00117_),
    .A1(net2402),
    .A2(net1843));
 sg13g2_nand2_1 _07260_ (.Y(_02474_),
    .A(net3235),
    .B(net1843));
 sg13g2_o21ai_1 _07261_ (.B1(_02474_),
    .Y(_00118_),
    .A1(net2397),
    .A2(net1843));
 sg13g2_nand2_1 _07262_ (.Y(_02475_),
    .A(_01751_),
    .B(_02341_));
 sg13g2_nand2_1 _07263_ (.Y(_02476_),
    .A(net1636),
    .B(net1833));
 sg13g2_o21ai_1 _07264_ (.B1(_02476_),
    .Y(_00119_),
    .A1(net2563),
    .A2(net1833));
 sg13g2_nand2_1 _07265_ (.Y(_02477_),
    .A(net1537),
    .B(net1835));
 sg13g2_o21ai_1 _07266_ (.B1(_02477_),
    .Y(_00120_),
    .A1(net2556),
    .A2(net1835));
 sg13g2_nand2_1 _07267_ (.Y(_02478_),
    .A(net1654),
    .B(net1841));
 sg13g2_o21ai_1 _07268_ (.B1(_02478_),
    .Y(_00121_),
    .A1(net2551),
    .A2(net1841));
 sg13g2_nand2_1 _07269_ (.Y(_02479_),
    .A(net3335),
    .B(net1839));
 sg13g2_o21ai_1 _07270_ (.B1(_02479_),
    .Y(_00122_),
    .A1(net2548),
    .A2(net1839));
 sg13g2_nand2_1 _07271_ (.Y(_02480_),
    .A(net2742),
    .B(net1839));
 sg13g2_o21ai_1 _07272_ (.B1(_02480_),
    .Y(_00123_),
    .A1(net2541),
    .A2(net1839));
 sg13g2_nand2_1 _07273_ (.Y(_02481_),
    .A(net2968),
    .B(net1840));
 sg13g2_o21ai_1 _07274_ (.B1(_02481_),
    .Y(_00124_),
    .A1(net2537),
    .A2(net1840));
 sg13g2_nand2_1 _07275_ (.Y(_02482_),
    .A(net3226),
    .B(net1840));
 sg13g2_o21ai_1 _07276_ (.B1(_02482_),
    .Y(_00125_),
    .A1(net2531),
    .A2(net1840));
 sg13g2_nand2_1 _07277_ (.Y(_02483_),
    .A(net3173),
    .B(net1839));
 sg13g2_o21ai_1 _07278_ (.B1(_02483_),
    .Y(_00126_),
    .A1(net2527),
    .A2(net1839));
 sg13g2_nand2_1 _07279_ (.Y(_02484_),
    .A(net1433),
    .B(net1839));
 sg13g2_o21ai_1 _07280_ (.B1(_02484_),
    .Y(_00127_),
    .A1(net2521),
    .A2(net1839));
 sg13g2_nand2_1 _07281_ (.Y(_02485_),
    .A(net2708),
    .B(net1838));
 sg13g2_o21ai_1 _07282_ (.B1(_02485_),
    .Y(_00128_),
    .A1(net2514),
    .A2(net1838));
 sg13g2_nand2_1 _07283_ (.Y(_02486_),
    .A(net1462),
    .B(net1838));
 sg13g2_o21ai_1 _07284_ (.B1(_02486_),
    .Y(_00129_),
    .A1(net2509),
    .A2(net1838));
 sg13g2_nand2_1 _07285_ (.Y(_02487_),
    .A(net1454),
    .B(net1838));
 sg13g2_o21ai_1 _07286_ (.B1(_02487_),
    .Y(_00130_),
    .A1(net2502),
    .A2(net1837));
 sg13g2_nand2_1 _07287_ (.Y(_02488_),
    .A(net1467),
    .B(net1838));
 sg13g2_o21ai_1 _07288_ (.B1(_02488_),
    .Y(_00131_),
    .A1(net2501),
    .A2(net1838));
 sg13g2_nand2_1 _07289_ (.Y(_02489_),
    .A(net3294),
    .B(net1837));
 sg13g2_o21ai_1 _07290_ (.B1(_02489_),
    .Y(_00132_),
    .A1(net2491),
    .A2(net1837));
 sg13g2_nand2_1 _07291_ (.Y(_02490_),
    .A(net1436),
    .B(net1836));
 sg13g2_o21ai_1 _07292_ (.B1(_02490_),
    .Y(_00133_),
    .A1(net2486),
    .A2(net1836));
 sg13g2_nand2_1 _07293_ (.Y(_02491_),
    .A(net2645),
    .B(net1837));
 sg13g2_o21ai_1 _07294_ (.B1(_02491_),
    .Y(_00134_),
    .A1(net2483),
    .A2(net1837));
 sg13g2_nand2_1 _07295_ (.Y(_02492_),
    .A(net1493),
    .B(net1841));
 sg13g2_o21ai_1 _07296_ (.B1(_02492_),
    .Y(_00135_),
    .A1(net2480),
    .A2(net1841));
 sg13g2_nand2_1 _07297_ (.Y(_02493_),
    .A(net3107),
    .B(net1837));
 sg13g2_o21ai_1 _07298_ (.B1(_02493_),
    .Y(_00136_),
    .A1(net2471),
    .A2(net1832));
 sg13g2_nand2_1 _07299_ (.Y(_02494_),
    .A(net2884),
    .B(net1837));
 sg13g2_o21ai_1 _07300_ (.B1(_02494_),
    .Y(_00137_),
    .A1(net2468),
    .A2(net1837));
 sg13g2_nand2_1 _07301_ (.Y(_02495_),
    .A(net2729),
    .B(net1836));
 sg13g2_o21ai_1 _07302_ (.B1(_02495_),
    .Y(_00138_),
    .A1(net2462),
    .A2(net1832));
 sg13g2_nand2_1 _07303_ (.Y(_02496_),
    .A(net3118),
    .B(net1834));
 sg13g2_o21ai_1 _07304_ (.B1(_02496_),
    .Y(_00139_),
    .A1(net2458),
    .A2(net1834));
 sg13g2_nand2_1 _07305_ (.Y(_02497_),
    .A(net1583),
    .B(net1834));
 sg13g2_o21ai_1 _07306_ (.B1(_02497_),
    .Y(_00140_),
    .A1(net2453),
    .A2(net1834));
 sg13g2_nand2_1 _07307_ (.Y(_02498_),
    .A(net3297),
    .B(net1841));
 sg13g2_o21ai_1 _07308_ (.B1(_02498_),
    .Y(_00141_),
    .A1(net2444),
    .A2(net1841));
 sg13g2_nand2_1 _07309_ (.Y(_02499_),
    .A(net3105),
    .B(net1834));
 sg13g2_o21ai_1 _07310_ (.B1(_02499_),
    .Y(_00142_),
    .A1(net2442),
    .A2(net1834));
 sg13g2_nand2_1 _07311_ (.Y(_02500_),
    .A(net1662),
    .B(net1834));
 sg13g2_o21ai_1 _07312_ (.B1(_02500_),
    .Y(_00143_),
    .A1(net2435),
    .A2(net1834));
 sg13g2_nand2_1 _07313_ (.Y(_02501_),
    .A(net2986),
    .B(net1833));
 sg13g2_o21ai_1 _07314_ (.B1(_02501_),
    .Y(_00144_),
    .A1(net2432),
    .A2(net1835));
 sg13g2_nand2_1 _07315_ (.Y(_02502_),
    .A(net1517),
    .B(net1833));
 sg13g2_o21ai_1 _07316_ (.B1(_02502_),
    .Y(_00145_),
    .A1(net2426),
    .A2(net1833));
 sg13g2_nand2_1 _07317_ (.Y(_02503_),
    .A(net2730),
    .B(net1833));
 sg13g2_o21ai_1 _07318_ (.B1(_02503_),
    .Y(_00146_),
    .A1(net2419),
    .A2(net1835));
 sg13g2_nand2_1 _07319_ (.Y(_02504_),
    .A(net1613),
    .B(net1833));
 sg13g2_o21ai_1 _07320_ (.B1(_02504_),
    .Y(_00147_),
    .A1(net2415),
    .A2(net1833));
 sg13g2_nand2_1 _07321_ (.Y(_02505_),
    .A(net2876),
    .B(net1832));
 sg13g2_o21ai_1 _07322_ (.B1(_02505_),
    .Y(_00148_),
    .A1(net2410),
    .A2(net1832));
 sg13g2_nand2_1 _07323_ (.Y(_02506_),
    .A(net2678),
    .B(net1832));
 sg13g2_o21ai_1 _07324_ (.B1(_02506_),
    .Y(_00149_),
    .A1(net2402),
    .A2(net1832));
 sg13g2_nand2_1 _07325_ (.Y(_02507_),
    .A(net2865),
    .B(net1832));
 sg13g2_o21ai_1 _07326_ (.B1(_02507_),
    .Y(_00150_),
    .A1(net2397),
    .A2(net1832));
 sg13g2_nand2b_2 _07327_ (.Y(_02508_),
    .B(_01716_),
    .A_N(net2307));
 sg13g2_nand2_1 _07328_ (.Y(_02509_),
    .A(net2740),
    .B(net1821));
 sg13g2_o21ai_1 _07329_ (.B1(_02509_),
    .Y(_00151_),
    .A1(net2560),
    .A2(net1821));
 sg13g2_nand2_1 _07330_ (.Y(_02510_),
    .A(net3223),
    .B(net1823));
 sg13g2_o21ai_1 _07331_ (.B1(_02510_),
    .Y(_00152_),
    .A1(net2556),
    .A2(net1824));
 sg13g2_nand2_1 _07332_ (.Y(_02511_),
    .A(net3045),
    .B(net1831));
 sg13g2_o21ai_1 _07333_ (.B1(_02511_),
    .Y(_00153_),
    .A1(net2554),
    .A2(net1831));
 sg13g2_nand2_1 _07334_ (.Y(_02512_),
    .A(net2665),
    .B(net1829));
 sg13g2_o21ai_1 _07335_ (.B1(_02512_),
    .Y(_00154_),
    .A1(net2544),
    .A2(net1829));
 sg13g2_nand2_1 _07336_ (.Y(_02513_),
    .A(net2663),
    .B(net1830));
 sg13g2_o21ai_1 _07337_ (.B1(_02513_),
    .Y(_00155_),
    .A1(net2538),
    .A2(net1830));
 sg13g2_nand2_1 _07338_ (.Y(_02514_),
    .A(net1713),
    .B(net1830));
 sg13g2_o21ai_1 _07339_ (.B1(_02514_),
    .Y(_00156_),
    .A1(net2533),
    .A2(net1830));
 sg13g2_nand2_1 _07340_ (.Y(_02515_),
    .A(net2682),
    .B(net1829));
 sg13g2_o21ai_1 _07341_ (.B1(_02515_),
    .Y(_00157_),
    .A1(net2529),
    .A2(net1829));
 sg13g2_nand2_1 _07342_ (.Y(_02516_),
    .A(net3180),
    .B(net1829));
 sg13g2_o21ai_1 _07343_ (.B1(_02516_),
    .Y(_00158_),
    .A1(net2523),
    .A2(net1829));
 sg13g2_nand2_1 _07344_ (.Y(_02517_),
    .A(net2644),
    .B(net1826));
 sg13g2_o21ai_1 _07345_ (.B1(_02517_),
    .Y(_00159_),
    .A1(net2518),
    .A2(net1826));
 sg13g2_nand2_1 _07346_ (.Y(_02518_),
    .A(net2738),
    .B(net1826));
 sg13g2_o21ai_1 _07347_ (.B1(_02518_),
    .Y(_00160_),
    .A1(net2513),
    .A2(net1826));
 sg13g2_nand2_1 _07348_ (.Y(_02519_),
    .A(net3196),
    .B(net1827));
 sg13g2_o21ai_1 _07349_ (.B1(_02519_),
    .Y(_00161_),
    .A1(net2507),
    .A2(net1827));
 sg13g2_nand2_1 _07350_ (.Y(_02520_),
    .A(net3109),
    .B(net1826));
 sg13g2_o21ai_1 _07351_ (.B1(_02520_),
    .Y(_00162_),
    .A1(net2502),
    .A2(net1826));
 sg13g2_nand2_1 _07352_ (.Y(_02521_),
    .A(net1734),
    .B(net1826));
 sg13g2_o21ai_1 _07353_ (.B1(_02521_),
    .Y(_00163_),
    .A1(net2496),
    .A2(net1826));
 sg13g2_nand2_1 _07354_ (.Y(_02522_),
    .A(net2727),
    .B(net1827));
 sg13g2_o21ai_1 _07355_ (.B1(_02522_),
    .Y(_00164_),
    .A1(net2492),
    .A2(net1827));
 sg13g2_nand2_1 _07356_ (.Y(_02523_),
    .A(net3081),
    .B(net1822));
 sg13g2_o21ai_1 _07357_ (.B1(_02523_),
    .Y(_00165_),
    .A1(net2486),
    .A2(net1822));
 sg13g2_nand2_1 _07358_ (.Y(_02524_),
    .A(net3191),
    .B(net1828));
 sg13g2_o21ai_1 _07359_ (.B1(_02524_),
    .Y(_00166_),
    .A1(net2481),
    .A2(net1828));
 sg13g2_nand2_1 _07360_ (.Y(_02525_),
    .A(net2745),
    .B(net1829));
 sg13g2_o21ai_1 _07361_ (.B1(_02525_),
    .Y(_00167_),
    .A1(net2479),
    .A2(net1829));
 sg13g2_nand2_1 _07362_ (.Y(_02526_),
    .A(net3242),
    .B(net1828));
 sg13g2_o21ai_1 _07363_ (.B1(_02526_),
    .Y(_00168_),
    .A1(net2470),
    .A2(net1828));
 sg13g2_nand2_1 _07364_ (.Y(_02527_),
    .A(net3178),
    .B(net1828));
 sg13g2_o21ai_1 _07365_ (.B1(_02527_),
    .Y(_00169_),
    .A1(net2466),
    .A2(net1828));
 sg13g2_nand2_1 _07366_ (.Y(_02528_),
    .A(net2941),
    .B(net1822));
 sg13g2_o21ai_1 _07367_ (.B1(_02528_),
    .Y(_00170_),
    .A1(net2464),
    .A2(net1822));
 sg13g2_nand2_1 _07368_ (.Y(_02529_),
    .A(net1732),
    .B(net1822));
 sg13g2_o21ai_1 _07369_ (.B1(_02529_),
    .Y(_00171_),
    .A1(net2455),
    .A2(net1822));
 sg13g2_nand2_1 _07370_ (.Y(_02530_),
    .A(net1711),
    .B(net1823));
 sg13g2_o21ai_1 _07371_ (.B1(_02530_),
    .Y(_00172_),
    .A1(net2450),
    .A2(net1824));
 sg13g2_nand2_1 _07372_ (.Y(_02531_),
    .A(net3322),
    .B(net1831));
 sg13g2_o21ai_1 _07373_ (.B1(_02531_),
    .Y(_00173_),
    .A1(net2445),
    .A2(net1831));
 sg13g2_nand2_1 _07374_ (.Y(_02532_),
    .A(net3052),
    .B(net1822));
 sg13g2_o21ai_1 _07375_ (.B1(_02532_),
    .Y(_00174_),
    .A1(net2439),
    .A2(net1822));
 sg13g2_nand2_1 _07376_ (.Y(_02533_),
    .A(net2733),
    .B(net1831));
 sg13g2_o21ai_1 _07377_ (.B1(_02533_),
    .Y(_00175_),
    .A1(net2436),
    .A2(net1831));
 sg13g2_nand2_1 _07378_ (.Y(_02534_),
    .A(net1626),
    .B(net1823));
 sg13g2_o21ai_1 _07379_ (.B1(_02534_),
    .Y(_00176_),
    .A1(net2428),
    .A2(net1823));
 sg13g2_nand2_1 _07380_ (.Y(_02535_),
    .A(net3098),
    .B(net1824));
 sg13g2_o21ai_1 _07381_ (.B1(_02535_),
    .Y(_00177_),
    .A1(net2425),
    .A2(net1824));
 sg13g2_nand2_1 _07382_ (.Y(_02536_),
    .A(net2735),
    .B(net1823));
 sg13g2_o21ai_1 _07383_ (.B1(_02536_),
    .Y(_00178_),
    .A1(net2418),
    .A2(net1823));
 sg13g2_nand2_1 _07384_ (.Y(_02537_),
    .A(net2985),
    .B(net1823));
 sg13g2_o21ai_1 _07385_ (.B1(_02537_),
    .Y(_00179_),
    .A1(net2413),
    .A2(net1823));
 sg13g2_nand2_1 _07386_ (.Y(_02538_),
    .A(net1595),
    .B(net1821));
 sg13g2_o21ai_1 _07387_ (.B1(_02538_),
    .Y(_00180_),
    .A1(net2410),
    .A2(net1821));
 sg13g2_nand2_1 _07388_ (.Y(_02539_),
    .A(net1532),
    .B(net1821));
 sg13g2_o21ai_1 _07389_ (.B1(_02539_),
    .Y(_00181_),
    .A1(net2403),
    .A2(net1821));
 sg13g2_nand2_1 _07390_ (.Y(_02540_),
    .A(net3172),
    .B(net1821));
 sg13g2_o21ai_1 _07391_ (.B1(_02540_),
    .Y(_00182_),
    .A1(net2397),
    .A2(net1821));
 sg13g2_nor2_1 _07392_ (.A(_01532_),
    .B(_02340_),
    .Y(_02541_));
 sg13g2_nand2b_1 _07393_ (.Y(_02542_),
    .B(net2325),
    .A_N(_02340_));
 sg13g2_nand2_1 _07394_ (.Y(_02543_),
    .A(_01616_),
    .B(_02541_));
 sg13g2_nand2_1 _07395_ (.Y(_02544_),
    .A(net1575),
    .B(net1811));
 sg13g2_o21ai_1 _07396_ (.B1(_02544_),
    .Y(_00183_),
    .A1(net2560),
    .A2(net1811));
 sg13g2_nand2_1 _07397_ (.Y(_02545_),
    .A(net3316),
    .B(net1814));
 sg13g2_o21ai_1 _07398_ (.B1(_02545_),
    .Y(_00184_),
    .A1(net2558),
    .A2(net1814));
 sg13g2_nand2_1 _07399_ (.Y(_02546_),
    .A(net2791),
    .B(net1818));
 sg13g2_o21ai_1 _07400_ (.B1(_02546_),
    .Y(_00185_),
    .A1(net2551),
    .A2(net1818));
 sg13g2_nand2_1 _07401_ (.Y(_02547_),
    .A(net3133),
    .B(net1819));
 sg13g2_o21ai_1 _07402_ (.B1(_02547_),
    .Y(_00186_),
    .A1(net2548),
    .A2(net1819));
 sg13g2_nand2_1 _07403_ (.Y(_02548_),
    .A(net1522),
    .B(net1819));
 sg13g2_o21ai_1 _07404_ (.B1(_02548_),
    .Y(_00187_),
    .A1(net2538),
    .A2(net1819));
 sg13g2_nand2_1 _07405_ (.Y(_02549_),
    .A(net2788),
    .B(net1819));
 sg13g2_o21ai_1 _07406_ (.B1(_02549_),
    .Y(_00188_),
    .A1(net2535),
    .A2(net1819));
 sg13g2_nand2_1 _07407_ (.Y(_02550_),
    .A(net3054),
    .B(net1819));
 sg13g2_o21ai_1 _07408_ (.B1(_02550_),
    .Y(_00189_),
    .A1(net2529),
    .A2(net1819));
 sg13g2_nand2_1 _07409_ (.Y(_02551_),
    .A(net2822),
    .B(net1816));
 sg13g2_o21ai_1 _07410_ (.B1(_02551_),
    .Y(_00190_),
    .A1(net2525),
    .A2(net1816));
 sg13g2_nand2_1 _07411_ (.Y(_02552_),
    .A(net1488),
    .B(net1816));
 sg13g2_o21ai_1 _07412_ (.B1(_02552_),
    .Y(_00191_),
    .A1(net2520),
    .A2(net1816));
 sg13g2_nand2_1 _07413_ (.Y(_02553_),
    .A(net1472),
    .B(net1815));
 sg13g2_o21ai_1 _07414_ (.B1(_02553_),
    .Y(_00192_),
    .A1(net2517),
    .A2(net1815));
 sg13g2_nand2_1 _07415_ (.Y(_02554_),
    .A(net3256),
    .B(net1815));
 sg13g2_o21ai_1 _07416_ (.B1(_02554_),
    .Y(_00193_),
    .A1(net2511),
    .A2(net1815));
 sg13g2_nand2_1 _07417_ (.Y(_02555_),
    .A(net1485),
    .B(net1817));
 sg13g2_o21ai_1 _07418_ (.B1(_02555_),
    .Y(_00194_),
    .A1(net2504),
    .A2(net1817));
 sg13g2_nand2_1 _07419_ (.Y(_02556_),
    .A(net1427),
    .B(net1815));
 sg13g2_o21ai_1 _07420_ (.B1(_02556_),
    .Y(_00195_),
    .A1(net2499),
    .A2(net1815));
 sg13g2_nand2_1 _07421_ (.Y(_02557_),
    .A(net3200),
    .B(net1815));
 sg13g2_o21ai_1 _07422_ (.B1(_02557_),
    .Y(_00196_),
    .A1(net2492),
    .A2(net1815));
 sg13g2_nand2_1 _07423_ (.Y(_02558_),
    .A(net1736),
    .B(net1812));
 sg13g2_o21ai_1 _07424_ (.B1(_02558_),
    .Y(_00197_),
    .A1(net2489),
    .A2(net1812));
 sg13g2_nand2_1 _07425_ (.Y(_02559_),
    .A(net1431),
    .B(net1812));
 sg13g2_o21ai_1 _07426_ (.B1(_02559_),
    .Y(_00198_),
    .A1(net2482),
    .A2(net1812));
 sg13g2_nand2_1 _07427_ (.Y(_02560_),
    .A(net3181),
    .B(net1818));
 sg13g2_o21ai_1 _07428_ (.B1(_02560_),
    .Y(_00199_),
    .A1(net2478),
    .A2(net1818));
 sg13g2_nand2_1 _07429_ (.Y(_02561_),
    .A(net2756),
    .B(net1817));
 sg13g2_o21ai_1 _07430_ (.B1(_02561_),
    .Y(_00200_),
    .A1(net2474),
    .A2(net1817));
 sg13g2_nand2_1 _07431_ (.Y(_02562_),
    .A(net1437),
    .B(net1817));
 sg13g2_o21ai_1 _07432_ (.B1(_02562_),
    .Y(_00201_),
    .A1(net2468),
    .A2(net1817));
 sg13g2_nand2_1 _07433_ (.Y(_02563_),
    .A(net1526),
    .B(net1812));
 sg13g2_o21ai_1 _07434_ (.B1(_02563_),
    .Y(_00202_),
    .A1(net2460),
    .A2(net1812));
 sg13g2_nand2_1 _07435_ (.Y(_02564_),
    .A(net2979),
    .B(net1812));
 sg13g2_o21ai_1 _07436_ (.B1(_02564_),
    .Y(_00203_),
    .A1(net2456),
    .A2(net1812));
 sg13g2_nand2_1 _07437_ (.Y(_02565_),
    .A(net1541),
    .B(net1814));
 sg13g2_o21ai_1 _07438_ (.B1(_02565_),
    .Y(_00204_),
    .A1(net2451),
    .A2(net1814));
 sg13g2_nand2_1 _07439_ (.Y(_02566_),
    .A(net3027),
    .B(net1818));
 sg13g2_o21ai_1 _07440_ (.B1(_02566_),
    .Y(_00205_),
    .A1(net2444),
    .A2(net1818));
 sg13g2_nand2_1 _07441_ (.Y(_02567_),
    .A(net3124),
    .B(net1813));
 sg13g2_o21ai_1 _07442_ (.B1(_02567_),
    .Y(_00206_),
    .A1(net2441),
    .A2(net1813));
 sg13g2_nand2_1 _07443_ (.Y(_02568_),
    .A(net2746),
    .B(net1818));
 sg13g2_o21ai_1 _07444_ (.B1(_02568_),
    .Y(_00207_),
    .A1(net2438),
    .A2(net1818));
 sg13g2_nand2_1 _07445_ (.Y(_02569_),
    .A(net3078),
    .B(net1813));
 sg13g2_o21ai_1 _07446_ (.B1(_02569_),
    .Y(_00208_),
    .A1(net2429),
    .A2(net1813));
 sg13g2_nand2_1 _07447_ (.Y(_02570_),
    .A(net3161),
    .B(net1813));
 sg13g2_o21ai_1 _07448_ (.B1(_02570_),
    .Y(_00209_),
    .A1(net2426),
    .A2(net1813));
 sg13g2_nand2_1 _07449_ (.Y(_02571_),
    .A(net3120),
    .B(net1814));
 sg13g2_o21ai_1 _07450_ (.B1(_02571_),
    .Y(_00210_),
    .A1(net2421),
    .A2(net1814));
 sg13g2_nand2_1 _07451_ (.Y(_02572_),
    .A(net1505),
    .B(net1813));
 sg13g2_o21ai_1 _07452_ (.B1(_02572_),
    .Y(_00211_),
    .A1(net2414),
    .A2(net1813));
 sg13g2_nand2_1 _07453_ (.Y(_02573_),
    .A(net3232),
    .B(net1811));
 sg13g2_o21ai_1 _07454_ (.B1(_02573_),
    .Y(_00212_),
    .A1(net2408),
    .A2(net1811));
 sg13g2_nand2_1 _07455_ (.Y(_02574_),
    .A(net1439),
    .B(net1811));
 sg13g2_o21ai_1 _07456_ (.B1(_02574_),
    .Y(_00213_),
    .A1(net2406),
    .A2(net1811));
 sg13g2_nand2_1 _07457_ (.Y(_02575_),
    .A(net1470),
    .B(net1811));
 sg13g2_o21ai_1 _07458_ (.B1(_02575_),
    .Y(_00214_),
    .A1(net2398),
    .A2(net1811));
 sg13g2_nand2_1 _07459_ (.Y(_02576_),
    .A(_01716_),
    .B(_02541_));
 sg13g2_nand2_1 _07460_ (.Y(_02577_),
    .A(net3271),
    .B(net1801));
 sg13g2_o21ai_1 _07461_ (.B1(_02577_),
    .Y(_00215_),
    .A1(net2560),
    .A2(net1801));
 sg13g2_nand2_1 _07462_ (.Y(_02578_),
    .A(net3005),
    .B(net1804));
 sg13g2_o21ai_1 _07463_ (.B1(_02578_),
    .Y(_00216_),
    .A1(net2558),
    .A2(net1804));
 sg13g2_nand2_1 _07464_ (.Y(_02579_),
    .A(net2634),
    .B(net1808));
 sg13g2_o21ai_1 _07465_ (.B1(_02579_),
    .Y(_00217_),
    .A1(net2551),
    .A2(net1808));
 sg13g2_nand2_1 _07466_ (.Y(_02580_),
    .A(net3152),
    .B(net1809));
 sg13g2_o21ai_1 _07467_ (.B1(_02580_),
    .Y(_00218_),
    .A1(net2546),
    .A2(net1809));
 sg13g2_nand2_1 _07468_ (.Y(_02581_),
    .A(net2650),
    .B(net1809));
 sg13g2_o21ai_1 _07469_ (.B1(_02581_),
    .Y(_00219_),
    .A1(net2538),
    .A2(net1809));
 sg13g2_nand2_1 _07470_ (.Y(_02582_),
    .A(net3067),
    .B(net1809));
 sg13g2_o21ai_1 _07471_ (.B1(_02582_),
    .Y(_00220_),
    .A1(net2535),
    .A2(net1809));
 sg13g2_nand2_1 _07472_ (.Y(_02583_),
    .A(net2812),
    .B(net1809));
 sg13g2_o21ai_1 _07473_ (.B1(_02583_),
    .Y(_00221_),
    .A1(net2529),
    .A2(net1809));
 sg13g2_nand2_1 _07474_ (.Y(_02584_),
    .A(net2704),
    .B(net1805));
 sg13g2_o21ai_1 _07475_ (.B1(_02584_),
    .Y(_00222_),
    .A1(net2525),
    .A2(net1805));
 sg13g2_nand2_1 _07476_ (.Y(_02585_),
    .A(net3387),
    .B(net1806));
 sg13g2_o21ai_1 _07477_ (.B1(_02585_),
    .Y(_00223_),
    .A1(net2520),
    .A2(net1806));
 sg13g2_nand2_1 _07478_ (.Y(_02586_),
    .A(net3108),
    .B(net1805));
 sg13g2_o21ai_1 _07479_ (.B1(_02586_),
    .Y(_00224_),
    .A1(net2512),
    .A2(net1805));
 sg13g2_nand2_1 _07480_ (.Y(_02587_),
    .A(net3149),
    .B(net1805));
 sg13g2_o21ai_1 _07481_ (.B1(_02587_),
    .Y(_00225_),
    .A1(net2511),
    .A2(net1805));
 sg13g2_nand2_1 _07482_ (.Y(_02588_),
    .A(net3063),
    .B(net1807));
 sg13g2_o21ai_1 _07483_ (.B1(_02588_),
    .Y(_00226_),
    .A1(net2504),
    .A2(net1807));
 sg13g2_nand2_1 _07484_ (.Y(_02589_),
    .A(net2924),
    .B(net1805));
 sg13g2_o21ai_1 _07485_ (.B1(_02589_),
    .Y(_00227_),
    .A1(net2499),
    .A2(net1805));
 sg13g2_nand2_1 _07486_ (.Y(_02590_),
    .A(net3245),
    .B(net1806));
 sg13g2_o21ai_1 _07487_ (.B1(_02590_),
    .Y(_00228_),
    .A1(net2492),
    .A2(net1806));
 sg13g2_nand2_1 _07488_ (.Y(_02591_),
    .A(net2826),
    .B(net1802));
 sg13g2_o21ai_1 _07489_ (.B1(_02591_),
    .Y(_00229_),
    .A1(net2488),
    .A2(net1802));
 sg13g2_nand2_1 _07490_ (.Y(_02592_),
    .A(net1503),
    .B(net1802));
 sg13g2_o21ai_1 _07491_ (.B1(_02592_),
    .Y(_00230_),
    .A1(net2482),
    .A2(net1802));
 sg13g2_nand2_1 _07492_ (.Y(_02593_),
    .A(net2773),
    .B(net1808));
 sg13g2_o21ai_1 _07493_ (.B1(_02593_),
    .Y(_00231_),
    .A1(net2478),
    .A2(net1808));
 sg13g2_nand2_1 _07494_ (.Y(_02594_),
    .A(net3038),
    .B(net1807));
 sg13g2_o21ai_1 _07495_ (.B1(_02594_),
    .Y(_00232_),
    .A1(net2474),
    .A2(net1807));
 sg13g2_nand2_1 _07496_ (.Y(_02595_),
    .A(net2615),
    .B(net1807));
 sg13g2_o21ai_1 _07497_ (.B1(_02595_),
    .Y(_00233_),
    .A1(net2468),
    .A2(net1807));
 sg13g2_nand2_1 _07498_ (.Y(_02596_),
    .A(net2801),
    .B(net1802));
 sg13g2_o21ai_1 _07499_ (.B1(_02596_),
    .Y(_00234_),
    .A1(net2460),
    .A2(net1802));
 sg13g2_nand2_1 _07500_ (.Y(_02597_),
    .A(net3244),
    .B(net1802));
 sg13g2_o21ai_1 _07501_ (.B1(_02597_),
    .Y(_00235_),
    .A1(net2456),
    .A2(net1802));
 sg13g2_nand2_1 _07502_ (.Y(_02598_),
    .A(net3177),
    .B(net1804));
 sg13g2_o21ai_1 _07503_ (.B1(_02598_),
    .Y(_00236_),
    .A1(net2451),
    .A2(net1804));
 sg13g2_nand2_1 _07504_ (.Y(_02599_),
    .A(net2805),
    .B(net1808));
 sg13g2_o21ai_1 _07505_ (.B1(_02599_),
    .Y(_00237_),
    .A1(net2444),
    .A2(net1808));
 sg13g2_nand2_1 _07506_ (.Y(_02600_),
    .A(net2863),
    .B(net1803));
 sg13g2_o21ai_1 _07507_ (.B1(_02600_),
    .Y(_00238_),
    .A1(net2441),
    .A2(net1803));
 sg13g2_nand2_1 _07508_ (.Y(_02601_),
    .A(net1603),
    .B(net1808));
 sg13g2_o21ai_1 _07509_ (.B1(_02601_),
    .Y(_00239_),
    .A1(net2437),
    .A2(net1808));
 sg13g2_nand2_1 _07510_ (.Y(_02602_),
    .A(net2873),
    .B(net1803));
 sg13g2_o21ai_1 _07511_ (.B1(_02602_),
    .Y(_00240_),
    .A1(net2429),
    .A2(net1803));
 sg13g2_nand2_1 _07512_ (.Y(_02603_),
    .A(net1587),
    .B(net1803));
 sg13g2_o21ai_1 _07513_ (.B1(_02603_),
    .Y(_00241_),
    .A1(net2426),
    .A2(net1803));
 sg13g2_nand2_1 _07514_ (.Y(_02604_),
    .A(net2818),
    .B(net1804));
 sg13g2_o21ai_1 _07515_ (.B1(_02604_),
    .Y(_00242_),
    .A1(net2421),
    .A2(net1804));
 sg13g2_nand2_1 _07516_ (.Y(_02605_),
    .A(net2966),
    .B(net1803));
 sg13g2_o21ai_1 _07517_ (.B1(_02605_),
    .Y(_00243_),
    .A1(net2414),
    .A2(net1803));
 sg13g2_nand2_1 _07518_ (.Y(_02606_),
    .A(net3066),
    .B(net1801));
 sg13g2_o21ai_1 _07519_ (.B1(_02606_),
    .Y(_00244_),
    .A1(net2408),
    .A2(net1801));
 sg13g2_nand2_1 _07520_ (.Y(_02607_),
    .A(net1740),
    .B(net1801));
 sg13g2_o21ai_1 _07521_ (.B1(_02607_),
    .Y(_00245_),
    .A1(net2406),
    .A2(net1801));
 sg13g2_nand2_1 _07522_ (.Y(_02608_),
    .A(net2862),
    .B(net1801));
 sg13g2_o21ai_1 _07523_ (.B1(_02608_),
    .Y(_00246_),
    .A1(net2401),
    .A2(net1801));
 sg13g2_nand2_1 _07524_ (.Y(_02609_),
    .A(_01751_),
    .B(_02541_));
 sg13g2_nand2_1 _07525_ (.Y(_02610_),
    .A(net1696),
    .B(net1791));
 sg13g2_o21ai_1 _07526_ (.B1(_02610_),
    .Y(_00247_),
    .A1(net2560),
    .A2(net1791));
 sg13g2_nand2_1 _07527_ (.Y(_02611_),
    .A(net3175),
    .B(net1794));
 sg13g2_o21ai_1 _07528_ (.B1(_02611_),
    .Y(_00248_),
    .A1(net2558),
    .A2(net1794));
 sg13g2_nand2_1 _07529_ (.Y(_02612_),
    .A(net2664),
    .B(net1798));
 sg13g2_o21ai_1 _07530_ (.B1(_02612_),
    .Y(_00249_),
    .A1(net2551),
    .A2(net1798));
 sg13g2_nand2_1 _07531_ (.Y(_02613_),
    .A(net3184),
    .B(net1799));
 sg13g2_o21ai_1 _07532_ (.B1(_02613_),
    .Y(_00250_),
    .A1(net2546),
    .A2(net1799));
 sg13g2_nand2_1 _07533_ (.Y(_02614_),
    .A(net2903),
    .B(net1799));
 sg13g2_o21ai_1 _07534_ (.B1(_02614_),
    .Y(_00251_),
    .A1(net2538),
    .A2(net1798));
 sg13g2_nand2_1 _07535_ (.Y(_02615_),
    .A(net1726),
    .B(net1799));
 sg13g2_o21ai_1 _07536_ (.B1(_02615_),
    .Y(_00252_),
    .A1(net2535),
    .A2(net1799));
 sg13g2_nand2_1 _07537_ (.Y(_02616_),
    .A(net1430),
    .B(net1800));
 sg13g2_o21ai_1 _07538_ (.B1(_02616_),
    .Y(_00253_),
    .A1(net2529),
    .A2(net1799));
 sg13g2_nand2_1 _07539_ (.Y(_02617_),
    .A(net2763),
    .B(net1795));
 sg13g2_o21ai_1 _07540_ (.B1(_02617_),
    .Y(_00254_),
    .A1(net2525),
    .A2(net1795));
 sg13g2_nand2_1 _07541_ (.Y(_02618_),
    .A(net3344),
    .B(net1796));
 sg13g2_o21ai_1 _07542_ (.B1(_02618_),
    .Y(_00255_),
    .A1(net2520),
    .A2(net1796));
 sg13g2_nand2_1 _07543_ (.Y(_02619_),
    .A(net1692),
    .B(net1795));
 sg13g2_o21ai_1 _07544_ (.B1(_02619_),
    .Y(_00256_),
    .A1(net2512),
    .A2(net1795));
 sg13g2_nand2_1 _07545_ (.Y(_02620_),
    .A(net2945),
    .B(net1795));
 sg13g2_o21ai_1 _07546_ (.B1(_02620_),
    .Y(_00257_),
    .A1(net2511),
    .A2(net1795));
 sg13g2_nand2_1 _07547_ (.Y(_02621_),
    .A(net3040),
    .B(net1797));
 sg13g2_o21ai_1 _07548_ (.B1(_02621_),
    .Y(_00258_),
    .A1(net2504),
    .A2(net1797));
 sg13g2_nand2_1 _07549_ (.Y(_02622_),
    .A(net2671),
    .B(net1795));
 sg13g2_o21ai_1 _07550_ (.B1(_02622_),
    .Y(_00259_),
    .A1(net2499),
    .A2(net1795));
 sg13g2_nand2_1 _07551_ (.Y(_02623_),
    .A(net2619),
    .B(net1796));
 sg13g2_o21ai_1 _07552_ (.B1(_02623_),
    .Y(_00260_),
    .A1(net2492),
    .A2(net1796));
 sg13g2_nand2_1 _07553_ (.Y(_02624_),
    .A(net3084),
    .B(net1792));
 sg13g2_o21ai_1 _07554_ (.B1(_02624_),
    .Y(_00261_),
    .A1(net2488),
    .A2(net1792));
 sg13g2_nand2_1 _07555_ (.Y(_02625_),
    .A(net1640),
    .B(net1792));
 sg13g2_o21ai_1 _07556_ (.B1(_02625_),
    .Y(_00262_),
    .A1(net2485),
    .A2(net1792));
 sg13g2_nand2_1 _07557_ (.Y(_02626_),
    .A(net1688),
    .B(net1798));
 sg13g2_o21ai_1 _07558_ (.B1(_02626_),
    .Y(_00263_),
    .A1(net2478),
    .A2(net1798));
 sg13g2_nand2_1 _07559_ (.Y(_02627_),
    .A(net2643),
    .B(net1797));
 sg13g2_o21ai_1 _07560_ (.B1(_02627_),
    .Y(_00264_),
    .A1(net2474),
    .A2(net1797));
 sg13g2_nand2_1 _07561_ (.Y(_02628_),
    .A(net1435),
    .B(net1797));
 sg13g2_o21ai_1 _07562_ (.B1(_02628_),
    .Y(_00265_),
    .A1(net2468),
    .A2(net1797));
 sg13g2_nand2_1 _07563_ (.Y(_02629_),
    .A(net1508),
    .B(net1792));
 sg13g2_o21ai_1 _07564_ (.B1(_02629_),
    .Y(_00266_),
    .A1(net2460),
    .A2(net1792));
 sg13g2_nand2_1 _07565_ (.Y(_02630_),
    .A(net3082),
    .B(net1792));
 sg13g2_o21ai_1 _07566_ (.B1(_02630_),
    .Y(_00267_),
    .A1(net2456),
    .A2(net1792));
 sg13g2_nand2_1 _07567_ (.Y(_02631_),
    .A(net3068),
    .B(net1794));
 sg13g2_o21ai_1 _07568_ (.B1(_02631_),
    .Y(_00268_),
    .A1(net2451),
    .A2(net1794));
 sg13g2_nand2_1 _07569_ (.Y(_02632_),
    .A(net2641),
    .B(net1798));
 sg13g2_o21ai_1 _07570_ (.B1(_02632_),
    .Y(_00269_),
    .A1(net2444),
    .A2(net1798));
 sg13g2_nand2_1 _07571_ (.Y(_02633_),
    .A(net1741),
    .B(net1793));
 sg13g2_o21ai_1 _07572_ (.B1(_02633_),
    .Y(_00270_),
    .A1(net2442),
    .A2(net1793));
 sg13g2_nand2_1 _07573_ (.Y(_02634_),
    .A(net2675),
    .B(net1798));
 sg13g2_o21ai_1 _07574_ (.B1(_02634_),
    .Y(_00271_),
    .A1(net2437),
    .A2(net1799));
 sg13g2_nand2_1 _07575_ (.Y(_02635_),
    .A(net1544),
    .B(net1793));
 sg13g2_o21ai_1 _07576_ (.B1(_02635_),
    .Y(_00272_),
    .A1(net2429),
    .A2(net1793));
 sg13g2_nand2_1 _07577_ (.Y(_02636_),
    .A(net2654),
    .B(net1793));
 sg13g2_o21ai_1 _07578_ (.B1(_02636_),
    .Y(_00273_),
    .A1(net2426),
    .A2(net1793));
 sg13g2_nand2_1 _07579_ (.Y(_02637_),
    .A(net2685),
    .B(net1794));
 sg13g2_o21ai_1 _07580_ (.B1(_02637_),
    .Y(_00274_),
    .A1(net2421),
    .A2(net1794));
 sg13g2_nand2_1 _07581_ (.Y(_02638_),
    .A(net2782),
    .B(net1793));
 sg13g2_o21ai_1 _07582_ (.B1(_02638_),
    .Y(_00275_),
    .A1(net2414),
    .A2(net1793));
 sg13g2_nand2_1 _07583_ (.Y(_02639_),
    .A(net1457),
    .B(net1791));
 sg13g2_o21ai_1 _07584_ (.B1(_02639_),
    .Y(_00276_),
    .A1(net2408),
    .A2(net1791));
 sg13g2_nand2_1 _07585_ (.Y(_02640_),
    .A(net3131),
    .B(net1791));
 sg13g2_o21ai_1 _07586_ (.B1(_02640_),
    .Y(_00277_),
    .A1(net2406),
    .A2(net1791));
 sg13g2_nand2_1 _07587_ (.Y(_02641_),
    .A(net3051),
    .B(net1791));
 sg13g2_o21ai_1 _07588_ (.B1(_02641_),
    .Y(_00278_),
    .A1(net2401),
    .A2(net1791));
 sg13g2_nand2_1 _07589_ (.Y(_02642_),
    .A(_01547_),
    .B(_02541_));
 sg13g2_nand2_1 _07590_ (.Y(_02643_),
    .A(net1666),
    .B(net1780));
 sg13g2_o21ai_1 _07591_ (.B1(_02643_),
    .Y(_00279_),
    .A1(net2561),
    .A2(net1780));
 sg13g2_nand2_1 _07592_ (.Y(_02644_),
    .A(net2963),
    .B(net1783));
 sg13g2_o21ai_1 _07593_ (.B1(_02644_),
    .Y(_00280_),
    .A1(net2558),
    .A2(net1783));
 sg13g2_nand2_1 _07594_ (.Y(_02645_),
    .A(net1700),
    .B(net1787));
 sg13g2_o21ai_1 _07595_ (.B1(_02645_),
    .Y(_00281_),
    .A1(net2551),
    .A2(net1787));
 sg13g2_nand2_1 _07596_ (.Y(_02646_),
    .A(net2750),
    .B(net1788));
 sg13g2_o21ai_1 _07597_ (.B1(_02646_),
    .Y(_00282_),
    .A1(net2548),
    .A2(net1788));
 sg13g2_nand2_1 _07598_ (.Y(_02647_),
    .A(net3217),
    .B(net1787));
 sg13g2_o21ai_1 _07599_ (.B1(_02647_),
    .Y(_00283_),
    .A1(net2539),
    .A2(net1787));
 sg13g2_nand2_1 _07600_ (.Y(_02648_),
    .A(net2996),
    .B(net1788));
 sg13g2_o21ai_1 _07601_ (.B1(_02648_),
    .Y(_00284_),
    .A1(net2535),
    .A2(net1788));
 sg13g2_nand2_1 _07602_ (.Y(_02649_),
    .A(net2851),
    .B(net1788));
 sg13g2_o21ai_1 _07603_ (.B1(_02649_),
    .Y(_00285_),
    .A1(net2532),
    .A2(net1788));
 sg13g2_nand2_1 _07604_ (.Y(_02650_),
    .A(net3257),
    .B(net1785));
 sg13g2_o21ai_1 _07605_ (.B1(_02650_),
    .Y(_00286_),
    .A1(net2525),
    .A2(net1785));
 sg13g2_nand2_1 _07606_ (.Y(_02651_),
    .A(net3187),
    .B(net1785));
 sg13g2_o21ai_1 _07607_ (.B1(_02651_),
    .Y(_00287_),
    .A1(net2520),
    .A2(net1785));
 sg13g2_nand2_1 _07608_ (.Y(_02652_),
    .A(net3292),
    .B(net1784));
 sg13g2_o21ai_1 _07609_ (.B1(_02652_),
    .Y(_00288_),
    .A1(net2517),
    .A2(net1784));
 sg13g2_nand2_1 _07610_ (.Y(_02653_),
    .A(net1682),
    .B(net1784));
 sg13g2_o21ai_1 _07611_ (.B1(_02653_),
    .Y(_00289_),
    .A1(net2511),
    .A2(net1784));
 sg13g2_nand2_1 _07612_ (.Y(_02654_),
    .A(net2747),
    .B(net1786));
 sg13g2_o21ai_1 _07613_ (.B1(_02654_),
    .Y(_00290_),
    .A1(net2504),
    .A2(net1786));
 sg13g2_nand2_1 _07614_ (.Y(_02655_),
    .A(net3233),
    .B(net1784));
 sg13g2_o21ai_1 _07615_ (.B1(_02655_),
    .Y(_00291_),
    .A1(net2499),
    .A2(net1784));
 sg13g2_nand2_1 _07616_ (.Y(_02656_),
    .A(net3103),
    .B(net1784));
 sg13g2_o21ai_1 _07617_ (.B1(_02656_),
    .Y(_00292_),
    .A1(net2492),
    .A2(net1784));
 sg13g2_nand2_1 _07618_ (.Y(_02657_),
    .A(net3102),
    .B(net1781));
 sg13g2_o21ai_1 _07619_ (.B1(_02657_),
    .Y(_00293_),
    .A1(net2489),
    .A2(net1781));
 sg13g2_nand2_1 _07620_ (.Y(_02658_),
    .A(net1451),
    .B(net1781));
 sg13g2_o21ai_1 _07621_ (.B1(_02658_),
    .Y(_00294_),
    .A1(net2482),
    .A2(net1781));
 sg13g2_nand2_1 _07622_ (.Y(_02659_),
    .A(net1615),
    .B(net1786));
 sg13g2_o21ai_1 _07623_ (.B1(_02659_),
    .Y(_00295_),
    .A1(net2478),
    .A2(net1786));
 sg13g2_nand2_1 _07624_ (.Y(_02660_),
    .A(net3336),
    .B(net1786));
 sg13g2_o21ai_1 _07625_ (.B1(_02660_),
    .Y(_00296_),
    .A1(net2474),
    .A2(net1786));
 sg13g2_nand2_1 _07626_ (.Y(_02661_),
    .A(net3195),
    .B(net1786));
 sg13g2_o21ai_1 _07627_ (.B1(_02661_),
    .Y(_00297_),
    .A1(net2468),
    .A2(net1786));
 sg13g2_nand2_1 _07628_ (.Y(_02662_),
    .A(net3286),
    .B(net1781));
 sg13g2_o21ai_1 _07629_ (.B1(_02662_),
    .Y(_00298_),
    .A1(net2460),
    .A2(net1781));
 sg13g2_nand2_1 _07630_ (.Y(_02663_),
    .A(net3306),
    .B(net1781));
 sg13g2_o21ai_1 _07631_ (.B1(_02663_),
    .Y(_00299_),
    .A1(net2456),
    .A2(net1781));
 sg13g2_nand2_1 _07632_ (.Y(_02664_),
    .A(net3025),
    .B(net1783));
 sg13g2_o21ai_1 _07633_ (.B1(_02664_),
    .Y(_00300_),
    .A1(net2451),
    .A2(net1783));
 sg13g2_nand2_1 _07634_ (.Y(_02665_),
    .A(net1727),
    .B(net1787));
 sg13g2_o21ai_1 _07635_ (.B1(_02665_),
    .Y(_00301_),
    .A1(net2444),
    .A2(net1787));
 sg13g2_nand2_1 _07636_ (.Y(_02666_),
    .A(net1577),
    .B(net1782));
 sg13g2_o21ai_1 _07637_ (.B1(_02666_),
    .Y(_00302_),
    .A1(net2442),
    .A2(net1782));
 sg13g2_nand2_1 _07638_ (.Y(_02667_),
    .A(net3159),
    .B(net1787));
 sg13g2_o21ai_1 _07639_ (.B1(_02667_),
    .Y(_00303_),
    .A1(net2438),
    .A2(net1787));
 sg13g2_nand2_1 _07640_ (.Y(_02668_),
    .A(net1652),
    .B(net1782));
 sg13g2_o21ai_1 _07641_ (.B1(_02668_),
    .Y(_00304_),
    .A1(net2429),
    .A2(net1782));
 sg13g2_nand2_1 _07642_ (.Y(_02669_),
    .A(net2932),
    .B(net1782));
 sg13g2_o21ai_1 _07643_ (.B1(_02669_),
    .Y(_00305_),
    .A1(net2426),
    .A2(net1782));
 sg13g2_nand2_1 _07644_ (.Y(_02670_),
    .A(net3313),
    .B(net1783));
 sg13g2_o21ai_1 _07645_ (.B1(_02670_),
    .Y(_00306_),
    .A1(net2421),
    .A2(net1783));
 sg13g2_nand2_1 _07646_ (.Y(_02671_),
    .A(net1705),
    .B(net1782));
 sg13g2_o21ai_1 _07647_ (.B1(_02671_),
    .Y(_00307_),
    .A1(net2414),
    .A2(net1782));
 sg13g2_nand2_1 _07648_ (.Y(_02672_),
    .A(net3407),
    .B(net1780));
 sg13g2_o21ai_1 _07649_ (.B1(_02672_),
    .Y(_00308_),
    .A1(net2408),
    .A2(net1780));
 sg13g2_nand2_1 _07650_ (.Y(_02673_),
    .A(net2855),
    .B(net1780));
 sg13g2_o21ai_1 _07651_ (.B1(_02673_),
    .Y(_00309_),
    .A1(net2406),
    .A2(net1780));
 sg13g2_nand2_1 _07652_ (.Y(_02674_),
    .A(net3310),
    .B(net1780));
 sg13g2_o21ai_1 _07653_ (.B1(_02674_),
    .Y(_00310_),
    .A1(net2401),
    .A2(net1780));
 sg13g2_and2_1 _07654_ (.A(_01427_),
    .B(net2376),
    .X(_02675_));
 sg13g2_nand2_1 _07655_ (.Y(_02676_),
    .A(_01427_),
    .B(net2376));
 sg13g2_o21ai_1 _07656_ (.B1(_02676_),
    .Y(_02677_),
    .A1(_01346_),
    .A2(_01651_));
 sg13g2_o21ai_1 _07657_ (.B1(_02677_),
    .Y(_02678_),
    .A1(_01346_),
    .A2(_01467_));
 sg13g2_a21o_1 _07658_ (.A2(_01454_),
    .A1(_01451_),
    .B1(net2572),
    .X(_02679_));
 sg13g2_a21oi_2 _07659_ (.B1(_01785_),
    .Y(_02680_),
    .A2(net2391),
    .A1(_01406_));
 sg13g2_o21ai_1 _07660_ (.B1(net2357),
    .Y(_02681_),
    .A1(_01458_),
    .A2(_02678_));
 sg13g2_a21oi_2 _07661_ (.B1(_02681_),
    .Y(_02682_),
    .A2(_02679_),
    .A1(_02675_));
 sg13g2_nand2_1 _07662_ (.Y(_02683_),
    .A(_01406_),
    .B(net2393));
 sg13g2_inv_2 _07663_ (.Y(_00471_),
    .A(net2366));
 sg13g2_nand3_1 _07664_ (.B(_02682_),
    .C(net2366),
    .A(net2602),
    .Y(_02684_));
 sg13g2_nor2_1 _07665_ (.A(net3340),
    .B(_02684_),
    .Y(_00311_));
 sg13g2_and3_1 _07666_ (.X(_02685_),
    .A(net3340),
    .B(net3818),
    .C(net3261));
 sg13g2_a21oi_1 _07667_ (.A1(\cpu.rf_ram_if.rcnt[0] ),
    .A2(\cpu.rf_ram_if.rcnt[1] ),
    .Y(_02686_),
    .B1(net3261));
 sg13g2_nor3_1 _07668_ (.A(_02684_),
    .B(_02685_),
    .C(net3262),
    .Y(_00312_));
 sg13g2_and2_1 _07669_ (.A(net3619),
    .B(_02685_),
    .X(_02687_));
 sg13g2_nor2_1 _07670_ (.A(net3619),
    .B(_02685_),
    .Y(_02688_));
 sg13g2_nor3_1 _07671_ (.A(_02684_),
    .B(_02687_),
    .C(net3620),
    .Y(_00313_));
 sg13g2_xnor2_1 _07672_ (.Y(_02689_),
    .A(net3723),
    .B(_02687_));
 sg13g2_nor2_1 _07673_ (.A(_02684_),
    .B(_02689_),
    .Y(_00314_));
 sg13g2_nand2_1 _07674_ (.Y(_02690_),
    .A(_01374_),
    .B(_01379_));
 sg13g2_a21oi_1 _07675_ (.A1(net2596),
    .A2(_02690_),
    .Y(_02691_),
    .B1(net2362));
 sg13g2_nand2_1 _07676_ (.Y(_02692_),
    .A(net2375),
    .B(net2318));
 sg13g2_a22oi_1 _07677_ (.Y(_02693_),
    .B1(net2318),
    .B2(net3586),
    .A2(net2360),
    .A1(\cpu.arbiter.i_wb_mem_rdt[15] ));
 sg13g2_nor2_1 _07678_ (.A(net3494),
    .B(net2129),
    .Y(_02694_));
 sg13g2_a21oi_1 _07679_ (.A1(net2129),
    .A2(net3587),
    .Y(_00315_),
    .B1(_02694_));
 sg13g2_nand2_1 _07680_ (.Y(_02695_),
    .A(net3494),
    .B(net2359));
 sg13g2_o21ai_1 _07681_ (.B1(net2317),
    .Y(_02696_),
    .A1(\cpu.arbiter.i_wb_cpu_dbus_dat[17] ),
    .A2(net2374));
 sg13g2_nor2_1 _07682_ (.A(net3485),
    .B(net2128),
    .Y(_02697_));
 sg13g2_a21oi_1 _07683_ (.A1(_02695_),
    .A2(_02696_),
    .Y(_00316_),
    .B1(_02697_));
 sg13g2_nand2_1 _07684_ (.Y(_02698_),
    .A(net3485),
    .B(net2359));
 sg13g2_o21ai_1 _07685_ (.B1(net2316),
    .Y(_02699_),
    .A1(\cpu.arbiter.i_wb_cpu_dbus_dat[18] ),
    .A2(net2374));
 sg13g2_nor2_1 _07686_ (.A(\cpu.arbiter.i_wb_mem_rdt[18] ),
    .B(net2128),
    .Y(_02700_));
 sg13g2_a21oi_1 _07687_ (.A1(_02698_),
    .A2(_02699_),
    .Y(_00317_),
    .B1(_02700_));
 sg13g2_nand2_1 _07688_ (.Y(_02701_),
    .A(net3565),
    .B(net2358));
 sg13g2_o21ai_1 _07689_ (.B1(net2316),
    .Y(_02702_),
    .A1(\cpu.arbiter.i_wb_cpu_dbus_dat[19] ),
    .A2(net2374));
 sg13g2_nor2_1 _07690_ (.A(\cpu.arbiter.i_wb_mem_rdt[19] ),
    .B(net2127),
    .Y(_02703_));
 sg13g2_a21oi_1 _07691_ (.A1(_02701_),
    .A2(_02702_),
    .Y(_00318_),
    .B1(_02703_));
 sg13g2_a22oi_1 _07692_ (.Y(_02704_),
    .B1(net2316),
    .B2(net3521),
    .A2(net2358),
    .A1(net3653));
 sg13g2_nor2_1 _07693_ (.A(net3558),
    .B(net2127),
    .Y(_02705_));
 sg13g2_a21oi_1 _07694_ (.A1(net2127),
    .A2(_02704_),
    .Y(_00319_),
    .B1(_02705_));
 sg13g2_nand2_1 _07695_ (.Y(_02706_),
    .A(net3558),
    .B(net2358));
 sg13g2_o21ai_1 _07696_ (.B1(net2316),
    .Y(_02707_),
    .A1(net3519),
    .A2(net2374));
 sg13g2_nor2_1 _07697_ (.A(\cpu.arbiter.i_wb_mem_rdt[21] ),
    .B(net2128),
    .Y(_02708_));
 sg13g2_a21oi_1 _07698_ (.A1(_02706_),
    .A2(_02707_),
    .Y(_00320_),
    .B1(_02708_));
 sg13g2_a22oi_1 _07699_ (.Y(_02709_),
    .B1(net2317),
    .B2(net3550),
    .A2(net2359),
    .A1(net3707));
 sg13g2_nor2_1 _07700_ (.A(net3680),
    .B(net2128),
    .Y(_02710_));
 sg13g2_a21oi_1 _07701_ (.A1(net2127),
    .A2(_02709_),
    .Y(_00321_),
    .B1(_02710_));
 sg13g2_nand2_1 _07702_ (.Y(_02711_),
    .A(net3680),
    .B(net2360));
 sg13g2_o21ai_1 _07703_ (.B1(net2317),
    .Y(_02712_),
    .A1(net3650),
    .A2(net2375));
 sg13g2_nor2_1 _07704_ (.A(\cpu.arbiter.i_wb_mem_rdt[23] ),
    .B(net2128),
    .Y(_02713_));
 sg13g2_a21oi_1 _07705_ (.A1(net3681),
    .A2(_02712_),
    .Y(_00322_),
    .B1(_02713_));
 sg13g2_a22oi_1 _07706_ (.Y(_02714_),
    .B1(net2317),
    .B2(\cpu.arbiter.i_wb_cpu_dbus_dat[24] ),
    .A2(net2359),
    .A1(net3728));
 sg13g2_nor2_1 _07707_ (.A(net3584),
    .B(net2128),
    .Y(_02715_));
 sg13g2_a21oi_1 _07708_ (.A1(net2129),
    .A2(net3729),
    .Y(_00323_),
    .B1(_02715_));
 sg13g2_nand2_1 _07709_ (.Y(_02716_),
    .A(net3584),
    .B(net2358));
 sg13g2_o21ai_1 _07710_ (.B1(net2316),
    .Y(_02717_),
    .A1(\cpu.arbiter.i_wb_cpu_dbus_dat[25] ),
    .A2(net2374));
 sg13g2_nor2_1 _07711_ (.A(net3556),
    .B(net2127),
    .Y(_02718_));
 sg13g2_a21oi_1 _07712_ (.A1(_02716_),
    .A2(_02717_),
    .Y(_00324_),
    .B1(_02718_));
 sg13g2_nand2_1 _07713_ (.Y(_02719_),
    .A(net3556),
    .B(net2358));
 sg13g2_o21ai_1 _07714_ (.B1(net2316),
    .Y(_02720_),
    .A1(\cpu.arbiter.i_wb_cpu_dbus_dat[26] ),
    .A2(net2374));
 sg13g2_nor2_1 _07715_ (.A(net3536),
    .B(net2127),
    .Y(_02721_));
 sg13g2_a21oi_1 _07716_ (.A1(_02719_),
    .A2(_02720_),
    .Y(_00325_),
    .B1(_02721_));
 sg13g2_nand2_1 _07717_ (.Y(_02722_),
    .A(net3536),
    .B(net2358));
 sg13g2_o21ai_1 _07718_ (.B1(net2316),
    .Y(_02723_),
    .A1(\cpu.arbiter.i_wb_cpu_dbus_dat[27] ),
    .A2(net2374));
 sg13g2_nor2_1 _07719_ (.A(\cpu.arbiter.i_wb_mem_rdt[27] ),
    .B(net2127),
    .Y(_02724_));
 sg13g2_a21oi_1 _07720_ (.A1(_02722_),
    .A2(_02723_),
    .Y(_00326_),
    .B1(_02724_));
 sg13g2_nand2_1 _07721_ (.Y(_02725_),
    .A(net3602),
    .B(net2358));
 sg13g2_o21ai_1 _07722_ (.B1(net2316),
    .Y(_02726_),
    .A1(\cpu.arbiter.i_wb_cpu_dbus_dat[28] ),
    .A2(net2374));
 sg13g2_nor2_1 _07723_ (.A(\cpu.arbiter.i_wb_mem_rdt[28] ),
    .B(net2127),
    .Y(_02727_));
 sg13g2_a21oi_1 _07724_ (.A1(_02725_),
    .A2(_02726_),
    .Y(_00327_),
    .B1(_02727_));
 sg13g2_nand2_1 _07725_ (.Y(_02728_),
    .A(net3613),
    .B(net2358));
 sg13g2_o21ai_1 _07726_ (.B1(net2317),
    .Y(_02729_),
    .A1(\cpu.arbiter.i_wb_cpu_dbus_dat[29] ),
    .A2(net2375));
 sg13g2_nor2_1 _07727_ (.A(net3591),
    .B(net2128),
    .Y(_02730_));
 sg13g2_a21oi_1 _07728_ (.A1(_02728_),
    .A2(_02729_),
    .Y(_00328_),
    .B1(_02730_));
 sg13g2_nand2_1 _07729_ (.Y(_02731_),
    .A(net3591),
    .B(net2360));
 sg13g2_o21ai_1 _07730_ (.B1(net2318),
    .Y(_02732_),
    .A1(net3450),
    .A2(net2375));
 sg13g2_nor2_1 _07731_ (.A(\cpu.arbiter.i_wb_mem_rdt[30] ),
    .B(net2129),
    .Y(_02733_));
 sg13g2_a21oi_1 _07732_ (.A1(net3592),
    .A2(_02732_),
    .Y(_00329_),
    .B1(_02733_));
 sg13g2_a22oi_1 _07733_ (.Y(_02734_),
    .B1(net2318),
    .B2(net3464),
    .A2(_01415_),
    .A1(\cpu.arbiter.i_wb_mem_rdt[30] ));
 sg13g2_nor2_1 _07734_ (.A(net3688),
    .B(net2129),
    .Y(_02735_));
 sg13g2_a21oi_1 _07735_ (.A1(net2129),
    .A2(_02734_),
    .Y(_00330_),
    .B1(_02735_));
 sg13g2_nor2_1 _07736_ (.A(_01334_),
    .B(_01339_),
    .Y(_00331_));
 sg13g2_nor2_1 _07737_ (.A(_01334_),
    .B(_01338_),
    .Y(_00332_));
 sg13g2_nor2_1 _07738_ (.A(_01334_),
    .B(_01337_),
    .Y(_00333_));
 sg13g2_nor2_1 _07739_ (.A(_01334_),
    .B(_01336_),
    .Y(_00334_));
 sg13g2_and2_1 _07740_ (.A(net2602),
    .B(net2),
    .X(_00335_));
 sg13g2_and2_1 _07741_ (.A(net2602),
    .B(net3),
    .X(_00336_));
 sg13g2_and2_1 _07742_ (.A(net2602),
    .B(net4),
    .X(_00337_));
 sg13g2_and2_1 _07743_ (.A(net2602),
    .B(net5),
    .X(_00338_));
 sg13g2_nand2_2 _07744_ (.Y(_02736_),
    .A(_01547_),
    .B(_01992_));
 sg13g2_nand2_1 _07745_ (.Y(_02737_),
    .A(net2810),
    .B(net1771));
 sg13g2_o21ai_1 _07746_ (.B1(_02737_),
    .Y(_00339_),
    .A1(net2562),
    .A2(net1771));
 sg13g2_nand2_1 _07747_ (.Y(_02738_),
    .A(net3093),
    .B(net1773));
 sg13g2_o21ai_1 _07748_ (.B1(_02738_),
    .Y(_00340_),
    .A1(net2558),
    .A2(net1773));
 sg13g2_nand2_1 _07749_ (.Y(_02739_),
    .A(net3319),
    .B(net1778));
 sg13g2_o21ai_1 _07750_ (.B1(_02739_),
    .Y(_00341_),
    .A1(net2552),
    .A2(net1778));
 sg13g2_nand2_1 _07751_ (.Y(_02740_),
    .A(net3153),
    .B(net1777));
 sg13g2_o21ai_1 _07752_ (.B1(_02740_),
    .Y(_00342_),
    .A1(net2546),
    .A2(net1777));
 sg13g2_nand2_1 _07753_ (.Y(_02741_),
    .A(net2766),
    .B(net1777));
 sg13g2_o21ai_1 _07754_ (.B1(_02741_),
    .Y(_00343_),
    .A1(net2542),
    .A2(net1777));
 sg13g2_nand2_1 _07755_ (.Y(_02742_),
    .A(net3258),
    .B(net1779));
 sg13g2_o21ai_1 _07756_ (.B1(_02742_),
    .Y(_00344_),
    .A1(net2536),
    .A2(net1778));
 sg13g2_nand2_1 _07757_ (.Y(_02743_),
    .A(net2699),
    .B(net1777));
 sg13g2_o21ai_1 _07758_ (.B1(_02743_),
    .Y(_00345_),
    .A1(net2530),
    .A2(net1777));
 sg13g2_nand2_1 _07759_ (.Y(_02744_),
    .A(net1728),
    .B(net1777));
 sg13g2_o21ai_1 _07760_ (.B1(_02744_),
    .Y(_00346_),
    .A1(net2526),
    .A2(net1777));
 sg13g2_nand2_1 _07761_ (.Y(_02745_),
    .A(net2880),
    .B(net1776));
 sg13g2_o21ai_1 _07762_ (.B1(_02745_),
    .Y(_00347_),
    .A1(net2521),
    .A2(net1776));
 sg13g2_nand2_1 _07763_ (.Y(_02746_),
    .A(net1557),
    .B(net1776));
 sg13g2_o21ai_1 _07764_ (.B1(_02746_),
    .Y(_00348_),
    .A1(net2514),
    .A2(net1776));
 sg13g2_nand2_1 _07765_ (.Y(_02747_),
    .A(net3137),
    .B(net1776));
 sg13g2_o21ai_1 _07766_ (.B1(_02747_),
    .Y(_00349_),
    .A1(net2509),
    .A2(net1776));
 sg13g2_nand2_1 _07767_ (.Y(_02748_),
    .A(net1712),
    .B(net1775));
 sg13g2_o21ai_1 _07768_ (.B1(_02748_),
    .Y(_00350_),
    .A1(net2506),
    .A2(net1775));
 sg13g2_nand2_1 _07769_ (.Y(_02749_),
    .A(net3139),
    .B(net1776));
 sg13g2_o21ai_1 _07770_ (.B1(_02749_),
    .Y(_00351_),
    .A1(net2501),
    .A2(net1776));
 sg13g2_nand2_1 _07771_ (.Y(_02750_),
    .A(net2933),
    .B(net1778));
 sg13g2_o21ai_1 _07772_ (.B1(_02750_),
    .Y(_00352_),
    .A1(net2493),
    .A2(net1778));
 sg13g2_nand2_1 _07773_ (.Y(_02751_),
    .A(net2843),
    .B(net1771));
 sg13g2_o21ai_1 _07774_ (.B1(_02751_),
    .Y(_00353_),
    .A1(net2489),
    .A2(net1774));
 sg13g2_nand2_1 _07775_ (.Y(_02752_),
    .A(net2823),
    .B(net1775));
 sg13g2_o21ai_1 _07776_ (.B1(_02752_),
    .Y(_00354_),
    .A1(net2483),
    .A2(net1775));
 sg13g2_nand2_1 _07777_ (.Y(_02753_),
    .A(net2783),
    .B(net1775));
 sg13g2_o21ai_1 _07778_ (.B1(_02753_),
    .Y(_00355_),
    .A1(net2477),
    .A2(net1775));
 sg13g2_nand2_1 _07779_ (.Y(_02754_),
    .A(net3216),
    .B(net1771));
 sg13g2_o21ai_1 _07780_ (.B1(_02754_),
    .Y(_00356_),
    .A1(net2471),
    .A2(net1771));
 sg13g2_nand2_1 _07781_ (.Y(_02755_),
    .A(net1691),
    .B(net1775));
 sg13g2_o21ai_1 _07782_ (.B1(_02755_),
    .Y(_00357_),
    .A1(net2466),
    .A2(net1775));
 sg13g2_nand2_1 _07783_ (.Y(_02756_),
    .A(net1440),
    .B(net1770));
 sg13g2_o21ai_1 _07784_ (.B1(_02756_),
    .Y(_00358_),
    .A1(net2460),
    .A2(net1770));
 sg13g2_nand2_1 _07785_ (.Y(_02757_),
    .A(net3013),
    .B(net1771));
 sg13g2_o21ai_1 _07786_ (.B1(_02757_),
    .Y(_00359_),
    .A1(net2456),
    .A2(net1771));
 sg13g2_nand2_1 _07787_ (.Y(_02758_),
    .A(net3252),
    .B(net1773));
 sg13g2_o21ai_1 _07788_ (.B1(_02758_),
    .Y(_00360_),
    .A1(net2451),
    .A2(net1774));
 sg13g2_nand2_1 _07789_ (.Y(_02759_),
    .A(net1543),
    .B(net1778));
 sg13g2_o21ai_1 _07790_ (.B1(_02759_),
    .Y(_00361_),
    .A1(net2447),
    .A2(net1778));
 sg13g2_nand2_1 _07791_ (.Y(_02760_),
    .A(net2864),
    .B(net1772));
 sg13g2_o21ai_1 _07792_ (.B1(_02760_),
    .Y(_00362_),
    .A1(net2442),
    .A2(net1772));
 sg13g2_nand2_1 _07793_ (.Y(_02761_),
    .A(net1667),
    .B(net1773));
 sg13g2_o21ai_1 _07794_ (.B1(_02761_),
    .Y(_00363_),
    .A1(net2438),
    .A2(net1773));
 sg13g2_nand2_1 _07795_ (.Y(_02762_),
    .A(net2705),
    .B(net1772));
 sg13g2_o21ai_1 _07796_ (.B1(_02762_),
    .Y(_00364_),
    .A1(net2431),
    .A2(net1772));
 sg13g2_nand2_1 _07797_ (.Y(_02763_),
    .A(net2789),
    .B(net1773));
 sg13g2_o21ai_1 _07798_ (.B1(_02763_),
    .Y(_00365_),
    .A1(net2424),
    .A2(net1773));
 sg13g2_nand2_1 _07799_ (.Y(_02764_),
    .A(net2784),
    .B(net1772));
 sg13g2_o21ai_1 _07800_ (.B1(_02764_),
    .Y(_00366_),
    .A1(net2420),
    .A2(net1772));
 sg13g2_nand2_1 _07801_ (.Y(_02765_),
    .A(net1607),
    .B(net1772));
 sg13g2_o21ai_1 _07802_ (.B1(_02765_),
    .Y(_00367_),
    .A1(net2416),
    .A2(net1772));
 sg13g2_nand2_1 _07803_ (.Y(_02766_),
    .A(net2939),
    .B(net1770));
 sg13g2_o21ai_1 _07804_ (.B1(_02766_),
    .Y(_00368_),
    .A1(net2411),
    .A2(net1770));
 sg13g2_nand2_1 _07805_ (.Y(_02767_),
    .A(net2841),
    .B(net1770));
 sg13g2_o21ai_1 _07806_ (.B1(_02767_),
    .Y(_00369_),
    .A1(net2404),
    .A2(net1770));
 sg13g2_nand2_1 _07807_ (.Y(_02768_),
    .A(net3130),
    .B(net1770));
 sg13g2_o21ai_1 _07808_ (.B1(_02768_),
    .Y(_00370_),
    .A1(net2399),
    .A2(net1770));
 sg13g2_nand2_2 _07809_ (.Y(_02769_),
    .A(_01716_),
    .B(_01992_));
 sg13g2_nand2_1 _07810_ (.Y(_02770_),
    .A(net3281),
    .B(net1760));
 sg13g2_o21ai_1 _07811_ (.B1(_02770_),
    .Y(_00371_),
    .A1(net2562),
    .A2(net1760));
 sg13g2_nand2_1 _07812_ (.Y(_02771_),
    .A(net2620),
    .B(net1763));
 sg13g2_o21ai_1 _07813_ (.B1(_02771_),
    .Y(_00372_),
    .A1(net2555),
    .A2(net1763));
 sg13g2_nand2_1 _07814_ (.Y(_02772_),
    .A(net3127),
    .B(net1768));
 sg13g2_o21ai_1 _07815_ (.B1(_02772_),
    .Y(_00373_),
    .A1(net2552),
    .A2(net1768));
 sg13g2_nand2_1 _07816_ (.Y(_02773_),
    .A(net3080),
    .B(net1767));
 sg13g2_o21ai_1 _07817_ (.B1(_02773_),
    .Y(_00374_),
    .A1(net2546),
    .A2(net1767));
 sg13g2_nand2_1 _07818_ (.Y(_02774_),
    .A(net1479),
    .B(net1767));
 sg13g2_o21ai_1 _07819_ (.B1(_02774_),
    .Y(_00375_),
    .A1(net2542),
    .A2(net1767));
 sg13g2_nand2_1 _07820_ (.Y(_02775_),
    .A(net3277),
    .B(net1769));
 sg13g2_o21ai_1 _07821_ (.B1(_02775_),
    .Y(_00376_),
    .A1(net2536),
    .A2(net1768));
 sg13g2_nand2_1 _07822_ (.Y(_02776_),
    .A(net1601),
    .B(net1767));
 sg13g2_o21ai_1 _07823_ (.B1(_02776_),
    .Y(_00377_),
    .A1(net2530),
    .A2(net1767));
 sg13g2_nand2_1 _07824_ (.Y(_02777_),
    .A(net2916),
    .B(net1767));
 sg13g2_o21ai_1 _07825_ (.B1(_02777_),
    .Y(_00378_),
    .A1(net2526),
    .A2(net1767));
 sg13g2_nand2_1 _07826_ (.Y(_02778_),
    .A(net2853),
    .B(net1766));
 sg13g2_o21ai_1 _07827_ (.B1(_02778_),
    .Y(_00379_),
    .A1(net2521),
    .A2(net1766));
 sg13g2_nand2_1 _07828_ (.Y(_02779_),
    .A(net3147),
    .B(net1766));
 sg13g2_o21ai_1 _07829_ (.B1(_02779_),
    .Y(_00380_),
    .A1(net2514),
    .A2(net1766));
 sg13g2_nand2_1 _07830_ (.Y(_02780_),
    .A(net2991),
    .B(net1766));
 sg13g2_o21ai_1 _07831_ (.B1(_02780_),
    .Y(_00381_),
    .A1(net2509),
    .A2(net1766));
 sg13g2_nand2_1 _07832_ (.Y(_02781_),
    .A(net1492),
    .B(net1765));
 sg13g2_o21ai_1 _07833_ (.B1(_02781_),
    .Y(_00382_),
    .A1(net2503),
    .A2(net1765));
 sg13g2_nand2_1 _07834_ (.Y(_02782_),
    .A(net2809),
    .B(net1766));
 sg13g2_o21ai_1 _07835_ (.B1(_02782_),
    .Y(_00383_),
    .A1(net2501),
    .A2(net1766));
 sg13g2_nand2_1 _07836_ (.Y(_02783_),
    .A(net2952),
    .B(net1768));
 sg13g2_o21ai_1 _07837_ (.B1(_02783_),
    .Y(_00384_),
    .A1(net2493),
    .A2(net1768));
 sg13g2_nand2_1 _07838_ (.Y(_02784_),
    .A(net3287),
    .B(net1761));
 sg13g2_o21ai_1 _07839_ (.B1(_02784_),
    .Y(_00385_),
    .A1(net2489),
    .A2(net1764));
 sg13g2_nand2_1 _07840_ (.Y(_02785_),
    .A(net1620),
    .B(net1765));
 sg13g2_o21ai_1 _07841_ (.B1(_02785_),
    .Y(_00386_),
    .A1(net2484),
    .A2(net1765));
 sg13g2_nand2_1 _07842_ (.Y(_02786_),
    .A(net3166),
    .B(net1765));
 sg13g2_o21ai_1 _07843_ (.B1(_02786_),
    .Y(_00387_),
    .A1(net2475),
    .A2(net1765));
 sg13g2_nand2_1 _07844_ (.Y(_02787_),
    .A(net2817),
    .B(net1761));
 sg13g2_o21ai_1 _07845_ (.B1(_02787_),
    .Y(_00388_),
    .A1(net2471),
    .A2(net1761));
 sg13g2_nand2_1 _07846_ (.Y(_02788_),
    .A(net1610),
    .B(net1765));
 sg13g2_o21ai_1 _07847_ (.B1(_02788_),
    .Y(_00389_),
    .A1(net2466),
    .A2(net1765));
 sg13g2_nand2_1 _07848_ (.Y(_02789_),
    .A(net3012),
    .B(net1760));
 sg13g2_o21ai_1 _07849_ (.B1(_02789_),
    .Y(_00390_),
    .A1(net2460),
    .A2(net1760));
 sg13g2_nand2_1 _07850_ (.Y(_02790_),
    .A(net2636),
    .B(net1761));
 sg13g2_o21ai_1 _07851_ (.B1(_02790_),
    .Y(_00391_),
    .A1(net2457),
    .A2(net1761));
 sg13g2_nand2_1 _07852_ (.Y(_02791_),
    .A(net2871),
    .B(net1763));
 sg13g2_o21ai_1 _07853_ (.B1(_02791_),
    .Y(_00392_),
    .A1(net2452),
    .A2(net1764));
 sg13g2_nand2_1 _07854_ (.Y(_02792_),
    .A(net2792),
    .B(net1768));
 sg13g2_o21ai_1 _07855_ (.B1(_02792_),
    .Y(_00393_),
    .A1(net2447),
    .A2(net1768));
 sg13g2_nand2_1 _07856_ (.Y(_02793_),
    .A(net1608),
    .B(net1762));
 sg13g2_o21ai_1 _07857_ (.B1(_02793_),
    .Y(_00394_),
    .A1(net2443),
    .A2(net1762));
 sg13g2_nand2_1 _07858_ (.Y(_02794_),
    .A(net2624),
    .B(net1763));
 sg13g2_o21ai_1 _07859_ (.B1(_02794_),
    .Y(_00395_),
    .A1(net2438),
    .A2(net1763));
 sg13g2_nand2_1 _07860_ (.Y(_02795_),
    .A(net2908),
    .B(net1762));
 sg13g2_o21ai_1 _07861_ (.B1(_02795_),
    .Y(_00396_),
    .A1(net2431),
    .A2(net1762));
 sg13g2_nand2_1 _07862_ (.Y(_02796_),
    .A(net3115),
    .B(net1763));
 sg13g2_o21ai_1 _07863_ (.B1(_02796_),
    .Y(_00397_),
    .A1(net2424),
    .A2(net1763));
 sg13g2_nand2_1 _07864_ (.Y(_02797_),
    .A(net2967),
    .B(net1762));
 sg13g2_o21ai_1 _07865_ (.B1(_02797_),
    .Y(_00398_),
    .A1(net2420),
    .A2(net1762));
 sg13g2_nand2_1 _07866_ (.Y(_02798_),
    .A(net1533),
    .B(net1762));
 sg13g2_o21ai_1 _07867_ (.B1(_02798_),
    .Y(_00399_),
    .A1(net2416),
    .A2(net1762));
 sg13g2_nand2_1 _07868_ (.Y(_02799_),
    .A(net3234),
    .B(net1761));
 sg13g2_o21ai_1 _07869_ (.B1(_02799_),
    .Y(_00400_),
    .A1(net2411),
    .A2(net1761));
 sg13g2_nand2_1 _07870_ (.Y(_02800_),
    .A(net3111),
    .B(net1760));
 sg13g2_o21ai_1 _07871_ (.B1(_02800_),
    .Y(_00401_),
    .A1(net2402),
    .A2(net1760));
 sg13g2_nand2_1 _07872_ (.Y(_02801_),
    .A(net3116),
    .B(net1760));
 sg13g2_o21ai_1 _07873_ (.B1(_02801_),
    .Y(_00402_),
    .A1(net2399),
    .A2(net1760));
 sg13g2_nor2_1 _07874_ (.A(\cpu.arbiter.i_wb_cpu_dbus_adr[3] ),
    .B(net2330),
    .Y(_02802_));
 sg13g2_a21oi_1 _07875_ (.A1(_01355_),
    .A2(net2331),
    .Y(_00403_),
    .B1(_02802_));
 sg13g2_mux2_1 _07876_ (.A0(\cpu.arbiter.i_wb_cpu_dbus_adr[4] ),
    .A1(net3676),
    .S(net2330),
    .X(_00404_));
 sg13g2_mux2_1 _07877_ (.A0(net3670),
    .A1(net3703),
    .S(net2330),
    .X(_00405_));
 sg13g2_mux2_1 _07878_ (.A0(net3654),
    .A1(net3670),
    .S(net2331),
    .X(_00406_));
 sg13g2_mux2_1 _07879_ (.A0(\cpu.arbiter.i_wb_cpu_dbus_adr[7] ),
    .A1(net3654),
    .S(net2331),
    .X(_00407_));
 sg13g2_mux2_1 _07880_ (.A0(net3664),
    .A1(\cpu.arbiter.i_wb_cpu_dbus_adr[7] ),
    .S(net2331),
    .X(_00408_));
 sg13g2_mux2_1 _07881_ (.A0(net3667),
    .A1(net3664),
    .S(net2330),
    .X(_00409_));
 sg13g2_mux2_1 _07882_ (.A0(net3700),
    .A1(net3667),
    .S(net2329),
    .X(_00410_));
 sg13g2_mux2_1 _07883_ (.A0(net3662),
    .A1(\cpu.arbiter.i_wb_cpu_dbus_adr[10] ),
    .S(net2329),
    .X(_00411_));
 sg13g2_mux2_1 _07884_ (.A0(net3685),
    .A1(net3662),
    .S(net2329),
    .X(_00412_));
 sg13g2_mux2_1 _07885_ (.A0(net3712),
    .A1(net3685),
    .S(net2326),
    .X(_00413_));
 sg13g2_mux2_1 _07886_ (.A0(net3671),
    .A1(\cpu.arbiter.i_wb_cpu_dbus_adr[13] ),
    .S(net2328),
    .X(_00414_));
 sg13g2_mux2_1 _07887_ (.A0(net3684),
    .A1(net3671),
    .S(net2326),
    .X(_00415_));
 sg13g2_mux2_1 _07888_ (.A0(net3528),
    .A1(\cpu.arbiter.i_wb_cpu_dbus_adr[15] ),
    .S(net2326),
    .X(_00416_));
 sg13g2_mux2_1 _07889_ (.A0(net3514),
    .A1(\cpu.arbiter.i_wb_cpu_dbus_adr[16] ),
    .S(net2326),
    .X(_00417_));
 sg13g2_mux2_1 _07890_ (.A0(net3541),
    .A1(net3514),
    .S(net2326),
    .X(_00418_));
 sg13g2_mux2_1 _07891_ (.A0(net3564),
    .A1(net3541),
    .S(net2326),
    .X(_00419_));
 sg13g2_mux2_1 _07892_ (.A0(net3622),
    .A1(net3564),
    .S(net2326),
    .X(_00420_));
 sg13g2_mux2_1 _07893_ (.A0(net3563),
    .A1(net3622),
    .S(net2326),
    .X(_00421_));
 sg13g2_mux2_1 _07894_ (.A0(net3561),
    .A1(net3563),
    .S(net2327),
    .X(_00422_));
 sg13g2_mux2_1 _07895_ (.A0(\cpu.arbiter.i_wb_cpu_dbus_adr[23] ),
    .A1(net3561),
    .S(net2327),
    .X(_00423_));
 sg13g2_mux2_1 _07896_ (.A0(net3506),
    .A1(\cpu.arbiter.i_wb_cpu_dbus_adr[23] ),
    .S(net2327),
    .X(_00424_));
 sg13g2_mux2_1 _07897_ (.A0(net3545),
    .A1(net3506),
    .S(net2327),
    .X(_00425_));
 sg13g2_mux2_1 _07898_ (.A0(net3560),
    .A1(net3545),
    .S(net2328),
    .X(_00426_));
 sg13g2_mux2_1 _07899_ (.A0(net3554),
    .A1(net3560),
    .S(net2327),
    .X(_00427_));
 sg13g2_mux2_1 _07900_ (.A0(\cpu.arbiter.i_wb_cpu_dbus_adr[28] ),
    .A1(net3554),
    .S(net2327),
    .X(_00428_));
 sg13g2_mux2_1 _07901_ (.A0(net3508),
    .A1(\cpu.arbiter.i_wb_cpu_dbus_adr[28] ),
    .S(net2327),
    .X(_00429_));
 sg13g2_mux2_1 _07902_ (.A0(net3540),
    .A1(net3508),
    .S(net2327),
    .X(_00430_));
 sg13g2_mux2_1 _07903_ (.A0(net3744),
    .A1(net3540),
    .S(net2331),
    .X(_00431_));
 sg13g2_o21ai_1 _07904_ (.B1(_01482_),
    .Y(_02803_),
    .A1(_01480_),
    .A2(_01481_));
 sg13g2_nand3_1 _07905_ (.B(_01483_),
    .C(_02803_),
    .A(_01455_),
    .Y(_02804_));
 sg13g2_nand2_1 _07906_ (.Y(_02805_),
    .A(net3744),
    .B(\cpu.cpu.bufreg.i_sh_signed ));
 sg13g2_o21ai_1 _07907_ (.B1(_02804_),
    .Y(_02806_),
    .A1(net2376),
    .A2(_02805_));
 sg13g2_mux2_1 _07908_ (.A0(net3744),
    .A1(_02806_),
    .S(_01471_),
    .X(_00432_));
 sg13g2_nor2b_1 _07909_ (.A(net3759),
    .B_N(\cpu.rf_ram_if.rgate ),
    .Y(_02807_));
 sg13g2_a22oi_1 _07910_ (.Y(_02808_),
    .B1(net3768),
    .B2(_02807_),
    .A2(net3606),
    .A1(net2581));
 sg13g2_a22oi_1 _07911_ (.Y(_02809_),
    .B1(net2133),
    .B2(net1572),
    .A2(net2177),
    .A1(net2740));
 sg13g2_a22oi_1 _07912_ (.Y(_02810_),
    .B1(net2221),
    .B2(net2839),
    .A2(net2268),
    .A1(net3032));
 sg13g2_a21oi_1 _07913_ (.A1(_02809_),
    .A2(_02810_),
    .Y(_02811_),
    .B1(net2308));
 sg13g2_a22oi_1 _07914_ (.Y(_02812_),
    .B1(net2133),
    .B2(net1707),
    .A2(net2177),
    .A1(net1685));
 sg13g2_a22oi_1 _07915_ (.Y(_02813_),
    .B1(net2221),
    .B2(net2683),
    .A2(net2268),
    .A1(net3202));
 sg13g2_a21oi_1 _07916_ (.A1(_02812_),
    .A2(_02813_),
    .Y(_02814_),
    .B1(net2082));
 sg13g2_a22oi_1 _07917_ (.Y(_02815_),
    .B1(net2134),
    .B2(net2824),
    .A2(net2178),
    .A1(net3142));
 sg13g2_a22oi_1 _07918_ (.Y(_02816_),
    .B1(net2222),
    .B2(net1446),
    .A2(net2269),
    .A1(net2913));
 sg13g2_a21oi_1 _07919_ (.A1(_02815_),
    .A2(_02816_),
    .Y(_02817_),
    .B1(net2260));
 sg13g2_a22oi_1 _07920_ (.Y(_02818_),
    .B1(net2134),
    .B2(net3144),
    .A2(net2178),
    .A1(net2918));
 sg13g2_a22oi_1 _07921_ (.Y(_02819_),
    .B1(net2222),
    .B2(net2829),
    .A2(net2269),
    .A1(net3021));
 sg13g2_a21oi_1 _07922_ (.A1(_02818_),
    .A2(_02819_),
    .Y(_02820_),
    .B1(net2097));
 sg13g2_a22oi_1 _07923_ (.Y(_02821_),
    .B1(net2134),
    .B2(net3197),
    .A2(net2178),
    .A1(net3281));
 sg13g2_a22oi_1 _07924_ (.Y(_02822_),
    .B1(net2222),
    .B2(net2719),
    .A2(net2269),
    .A1(net3793));
 sg13g2_a21oi_1 _07925_ (.A1(_02821_),
    .A2(_02822_),
    .Y(_02823_),
    .B1(net2077));
 sg13g2_a22oi_1 _07926_ (.Y(_02824_),
    .B1(net2133),
    .B2(net1696),
    .A2(net2177),
    .A1(net3271));
 sg13g2_a22oi_1 _07927_ (.Y(_02825_),
    .B1(net2221),
    .B2(net1575),
    .A2(net2268),
    .A1(net1666));
 sg13g2_a21oi_1 _07928_ (.A1(_02824_),
    .A2(_02825_),
    .Y(_02826_),
    .B1(net2067));
 sg13g2_a22oi_1 _07929_ (.Y(_02827_),
    .B1(net2134),
    .B2(net1636),
    .A2(net2178),
    .A1(net2807));
 sg13g2_a22oi_1 _07930_ (.Y(_02828_),
    .B1(net2222),
    .B2(net3251),
    .A2(net2269),
    .A1(net3337));
 sg13g2_a21oi_1 _07931_ (.A1(_02827_),
    .A2(_02828_),
    .Y(_02829_),
    .B1(net2072));
 sg13g2_a22oi_1 _07932_ (.Y(_02830_),
    .B1(net2133),
    .B2(net2898),
    .A2(net2177),
    .A1(net2711));
 sg13g2_a22oi_1 _07933_ (.Y(_02831_),
    .B1(net2221),
    .B2(net1630),
    .A2(net2268),
    .A1(net3156));
 sg13g2_a21oi_1 _07934_ (.A1(_02830_),
    .A2(_02831_),
    .Y(_02832_),
    .B1(net2102));
 sg13g2_nor4_1 _07935_ (.A(_02811_),
    .B(_02817_),
    .C(_02823_),
    .D(_02826_),
    .Y(_02833_));
 sg13g2_nor4_1 _07936_ (.A(_02814_),
    .B(_02820_),
    .C(_02829_),
    .D(_02832_),
    .Y(_02834_));
 sg13g2_a21oi_1 _07937_ (.A1(_02833_),
    .A2(_02834_),
    .Y(_00433_),
    .B1(net2384));
 sg13g2_a22oi_1 _07938_ (.Y(_02835_),
    .B1(net2150),
    .B2(net1537),
    .A2(net2194),
    .A1(net3128));
 sg13g2_a22oi_1 _07939_ (.Y(_02836_),
    .B1(net2236),
    .B2(net2710),
    .A2(net2281),
    .A1(net3268));
 sg13g2_a21oi_1 _07940_ (.A1(_02835_),
    .A2(_02836_),
    .Y(_02837_),
    .B1(net2073));
 sg13g2_a22oi_1 _07941_ (.Y(_02838_),
    .B1(net2148),
    .B2(net3064),
    .A2(net2192),
    .A1(net2785));
 sg13g2_a22oi_1 _07942_ (.Y(_02839_),
    .B1(net2234),
    .B2(net2707),
    .A2(net2281),
    .A1(net3163));
 sg13g2_a21oi_1 _07943_ (.A1(_02838_),
    .A2(_02839_),
    .Y(_02840_),
    .B1(net2261));
 sg13g2_a22oi_1 _07944_ (.Y(_02841_),
    .B1(net2149),
    .B2(net3303),
    .A2(net2193),
    .A1(net3223));
 sg13g2_a22oi_1 _07945_ (.Y(_02842_),
    .B1(net2235),
    .B2(net1709),
    .A2(net2282),
    .A1(\rf_ram.RAM[3][1] ));
 sg13g2_a21oi_1 _07946_ (.A1(_02841_),
    .A2(_02842_),
    .Y(_02843_),
    .B1(net2307));
 sg13g2_a22oi_1 _07947_ (.Y(_02844_),
    .B1(net2148),
    .B2(net3175),
    .A2(net2192),
    .A1(net3005));
 sg13g2_a22oi_1 _07948_ (.Y(_02845_),
    .B1(net2234),
    .B2(net3316),
    .A2(net2281),
    .A1(net3773));
 sg13g2_a21oi_1 _07949_ (.A1(_02844_),
    .A2(_02845_),
    .Y(_02846_),
    .B1(net2068));
 sg13g2_a22oi_1 _07950_ (.Y(_02847_),
    .B1(net2148),
    .B2(net3155),
    .A2(net2192),
    .A1(net2620));
 sg13g2_a22oi_1 _07951_ (.Y(_02848_),
    .B1(net2234),
    .B2(net1593),
    .A2(net2281),
    .A1(net3093));
 sg13g2_a21oi_1 _07952_ (.A1(_02847_),
    .A2(_02848_),
    .Y(_02849_),
    .B1(net2078));
 sg13g2_a22oi_1 _07953_ (.Y(_02850_),
    .B1(net2149),
    .B2(net1542),
    .A2(net2193),
    .A1(net2662));
 sg13g2_a22oi_1 _07954_ (.Y(_02851_),
    .B1(net2235),
    .B2(net2612),
    .A2(net2282),
    .A1(net2768));
 sg13g2_a21oi_1 _07955_ (.A1(_02850_),
    .A2(_02851_),
    .Y(_02852_),
    .B1(net2083));
 sg13g2_a22oi_1 _07956_ (.Y(_02853_),
    .B1(net2149),
    .B2(net1418),
    .A2(net2193),
    .A1(net1547));
 sg13g2_a22oi_1 _07957_ (.Y(_02854_),
    .B1(net2235),
    .B2(net2800),
    .A2(net2283),
    .A1(net1570));
 sg13g2_a21oi_1 _07958_ (.A1(_02853_),
    .A2(_02854_),
    .Y(_02855_),
    .B1(net2098));
 sg13g2_a22oi_1 _07959_ (.Y(_02856_),
    .B1(net2149),
    .B2(net1461),
    .A2(net2193),
    .A1(net1589));
 sg13g2_a22oi_1 _07960_ (.Y(_02857_),
    .B1(net2235),
    .B2(net3060),
    .A2(net2282),
    .A1(net3225));
 sg13g2_a21oi_1 _07961_ (.A1(_02856_),
    .A2(_02857_),
    .Y(_02858_),
    .B1(net2103));
 sg13g2_nor4_1 _07962_ (.A(_02837_),
    .B(_02840_),
    .C(_02849_),
    .D(_02855_),
    .Y(_02859_));
 sg13g2_nor4_1 _07963_ (.A(_02843_),
    .B(_02846_),
    .C(_02852_),
    .D(_02858_),
    .Y(_02860_));
 sg13g2_a21oi_1 _07964_ (.A1(_02859_),
    .A2(_02860_),
    .Y(_00434_),
    .B1(net2385));
 sg13g2_a22oi_1 _07965_ (.Y(_02861_),
    .B1(net2166),
    .B2(\rf_ram.RAM[18][2] ),
    .A2(net2210),
    .A1(\rf_ram.RAM[17][2] ));
 sg13g2_a22oi_1 _07966_ (.Y(_02862_),
    .B1(net2250),
    .B2(\rf_ram.RAM[16][2] ),
    .A2(net2297),
    .A1(\rf_ram.RAM[19][2] ));
 sg13g2_a21oi_1 _07967_ (.A1(_02861_),
    .A2(_02862_),
    .Y(_02863_),
    .B1(net2075));
 sg13g2_a22oi_1 _07968_ (.Y(_02864_),
    .B1(net2165),
    .B2(\rf_ram.RAM[30][2] ),
    .A2(net2209),
    .A1(\rf_ram.RAM[29][2] ));
 sg13g2_a22oi_1 _07969_ (.Y(_02865_),
    .B1(net2250),
    .B2(\rf_ram.RAM[28][2] ),
    .A2(net2296),
    .A1(\rf_ram.RAM[31][2] ));
 sg13g2_a21oi_1 _07970_ (.A1(_02864_),
    .A2(_02865_),
    .Y(_02866_),
    .B1(net2080));
 sg13g2_a22oi_1 _07971_ (.Y(_02867_),
    .B1(net2164),
    .B2(\rf_ram.RAM[22][2] ),
    .A2(net2208),
    .A1(\rf_ram.RAM[21][2] ));
 sg13g2_a22oi_1 _07972_ (.Y(_02868_),
    .B1(net2251),
    .B2(\rf_ram.RAM[20][2] ),
    .A2(net2296),
    .A1(\rf_ram.RAM[23][2] ));
 sg13g2_a21oi_1 _07973_ (.A1(_02867_),
    .A2(_02868_),
    .Y(_02869_),
    .B1(net2069));
 sg13g2_a22oi_1 _07974_ (.Y(_02870_),
    .B1(net2164),
    .B2(\rf_ram.RAM[2][2] ),
    .A2(net2208),
    .A1(\rf_ram.RAM[1][2] ));
 sg13g2_a22oi_1 _07975_ (.Y(_02871_),
    .B1(net2250),
    .B2(\rf_ram.RAM[0][2] ),
    .A2(net2297),
    .A1(\rf_ram.RAM[3][2] ));
 sg13g2_a21oi_1 _07976_ (.A1(_02870_),
    .A2(_02871_),
    .Y(_02872_),
    .B1(net2310));
 sg13g2_a22oi_1 _07977_ (.Y(_02873_),
    .B1(net2164),
    .B2(\rf_ram.RAM[26][2] ),
    .A2(net2208),
    .A1(\rf_ram.RAM[25][2] ));
 sg13g2_a22oi_1 _07978_ (.Y(_02874_),
    .B1(net2251),
    .B2(\rf_ram.RAM[24][2] ),
    .A2(net2298),
    .A1(\rf_ram.RAM[27][2] ));
 sg13g2_a21oi_1 _07979_ (.A1(_02873_),
    .A2(_02874_),
    .Y(_02875_),
    .B1(net2085));
 sg13g2_a22oi_1 _07980_ (.Y(_02876_),
    .B1(net2165),
    .B2(\rf_ram.RAM[14][2] ),
    .A2(net2209),
    .A1(\rf_ram.RAM[13][2] ));
 sg13g2_a22oi_1 _07981_ (.Y(_02877_),
    .B1(net2252),
    .B2(\rf_ram.RAM[12][2] ),
    .A2(net2298),
    .A1(\rf_ram.RAM[15][2] ));
 sg13g2_a21oi_1 _07982_ (.A1(_02876_),
    .A2(_02877_),
    .Y(_02878_),
    .B1(net2104));
 sg13g2_a22oi_1 _07983_ (.Y(_02879_),
    .B1(net2166),
    .B2(\rf_ram.RAM[6][2] ),
    .A2(net2210),
    .A1(\rf_ram.RAM[5][2] ));
 sg13g2_a22oi_1 _07984_ (.Y(_02880_),
    .B1(net2250),
    .B2(\rf_ram.RAM[4][2] ),
    .A2(net2297),
    .A1(\rf_ram.RAM[7][2] ));
 sg13g2_a21oi_1 _07985_ (.A1(_02879_),
    .A2(_02880_),
    .Y(_02881_),
    .B1(net2262));
 sg13g2_a22oi_1 _07986_ (.Y(_02882_),
    .B1(net2164),
    .B2(net1619),
    .A2(net2208),
    .A1(\rf_ram.RAM[9][2] ));
 sg13g2_a22oi_1 _07987_ (.Y(_02883_),
    .B1(net2251),
    .B2(net3810),
    .A2(net2296),
    .A1(\rf_ram.RAM[11][2] ));
 sg13g2_a21oi_1 _07988_ (.A1(_02882_),
    .A2(_02883_),
    .Y(_02884_),
    .B1(net2099));
 sg13g2_nor4_1 _07989_ (.A(_02863_),
    .B(_02869_),
    .C(_02881_),
    .D(net3811),
    .Y(_02885_));
 sg13g2_nor4_1 _07990_ (.A(_02866_),
    .B(_02872_),
    .C(_02875_),
    .D(_02878_),
    .Y(_02886_));
 sg13g2_a21oi_1 _07991_ (.A1(net3812),
    .A2(_02886_),
    .Y(_00435_),
    .B1(net2387));
 sg13g2_a22oi_1 _07992_ (.Y(_02887_),
    .B1(net2165),
    .B2(\rf_ram.RAM[2][3] ),
    .A2(net2209),
    .A1(\rf_ram.RAM[1][3] ));
 sg13g2_a22oi_1 _07993_ (.Y(_02888_),
    .B1(net2250),
    .B2(\rf_ram.RAM[0][3] ),
    .A2(net2297),
    .A1(\rf_ram.RAM[3][3] ));
 sg13g2_a21oi_1 _07994_ (.A1(_02887_),
    .A2(_02888_),
    .Y(_02889_),
    .B1(net2310));
 sg13g2_a22oi_1 _07995_ (.Y(_02890_),
    .B1(net2166),
    .B2(\rf_ram.RAM[10][3] ),
    .A2(net2210),
    .A1(\rf_ram.RAM[9][3] ));
 sg13g2_a22oi_1 _07996_ (.Y(_02891_),
    .B1(net2250),
    .B2(\rf_ram.RAM[8][3] ),
    .A2(net2297),
    .A1(\rf_ram.RAM[11][3] ));
 sg13g2_a21oi_1 _07997_ (.A1(_02890_),
    .A2(_02891_),
    .Y(_02892_),
    .B1(net2099));
 sg13g2_a22oi_1 _07998_ (.Y(_02893_),
    .B1(net2169),
    .B2(net3335),
    .A2(net2213),
    .A1(net3264));
 sg13g2_a22oi_1 _07999_ (.Y(_02894_),
    .B1(net2255),
    .B2(net3243),
    .A2(net2301),
    .A1(net2958));
 sg13g2_a21oi_1 _08000_ (.A1(_02893_),
    .A2(_02894_),
    .Y(_02895_),
    .B1(net2075));
 sg13g2_a22oi_1 _08001_ (.Y(_02896_),
    .B1(net2169),
    .B2(net1644),
    .A2(net2213),
    .A1(net2901));
 sg13g2_a22oi_1 _08002_ (.Y(_02897_),
    .B1(net2255),
    .B2(net3083),
    .A2(net2301),
    .A1(net3796));
 sg13g2_a21oi_1 _08003_ (.A1(_02896_),
    .A2(_02897_),
    .Y(_02898_),
    .B1(net2104));
 sg13g2_a22oi_1 _08004_ (.Y(_02899_),
    .B1(net2165),
    .B2(\rf_ram.RAM[26][3] ),
    .A2(net2209),
    .A1(\rf_ram.RAM[25][3] ));
 sg13g2_a22oi_1 _08005_ (.Y(_02900_),
    .B1(net2250),
    .B2(\rf_ram.RAM[24][3] ),
    .A2(net2297),
    .A1(\rf_ram.RAM[27][3] ));
 sg13g2_a21oi_1 _08006_ (.A1(_02899_),
    .A2(_02900_),
    .Y(_02901_),
    .B1(net2085));
 sg13g2_a22oi_1 _08007_ (.Y(_02902_),
    .B1(net2169),
    .B2(net2808),
    .A2(net2213),
    .A1(net2659));
 sg13g2_a22oi_1 _08008_ (.Y(_02903_),
    .B1(net2255),
    .B2(net1634),
    .A2(net2301),
    .A1(net2893));
 sg13g2_a21oi_1 _08009_ (.A1(_02902_),
    .A2(_02903_),
    .Y(_02904_),
    .B1(net2262));
 sg13g2_a22oi_1 _08010_ (.Y(_02905_),
    .B1(net2171),
    .B2(net3184),
    .A2(net2215),
    .A1(net3152));
 sg13g2_a22oi_1 _08011_ (.Y(_02906_),
    .B1(net2257),
    .B2(net3133),
    .A2(net2303),
    .A1(net2750));
 sg13g2_a21oi_1 _08012_ (.A1(_02905_),
    .A2(_02906_),
    .Y(_02907_),
    .B1(net2069));
 sg13g2_a22oi_1 _08013_ (.Y(_02908_),
    .B1(net2169),
    .B2(net1714),
    .A2(net2213),
    .A1(net3080));
 sg13g2_a22oi_1 _08014_ (.Y(_02909_),
    .B1(net2255),
    .B2(net2687),
    .A2(net2301),
    .A1(net3153));
 sg13g2_a21oi_1 _08015_ (.A1(_02908_),
    .A2(_02909_),
    .Y(_02910_),
    .B1(net2080));
 sg13g2_nor4_1 _08016_ (.A(_02889_),
    .B(_02895_),
    .C(_02901_),
    .D(_02907_),
    .Y(_02911_));
 sg13g2_nor4_1 _08017_ (.A(_02892_),
    .B(_02898_),
    .C(_02904_),
    .D(_02910_),
    .Y(_02912_));
 sg13g2_a21oi_1 _08018_ (.A1(_02911_),
    .A2(_02912_),
    .Y(_00436_),
    .B1(net2386));
 sg13g2_a22oi_1 _08019_ (.Y(_02913_),
    .B1(net2165),
    .B2(\rf_ram.RAM[22][4] ),
    .A2(net2209),
    .A1(\rf_ram.RAM[21][4] ));
 sg13g2_a22oi_1 _08020_ (.Y(_02914_),
    .B1(net2250),
    .B2(\rf_ram.RAM[20][4] ),
    .A2(net2297),
    .A1(\rf_ram.RAM[23][4] ));
 sg13g2_a21oi_1 _08021_ (.A1(_02913_),
    .A2(_02914_),
    .Y(_02915_),
    .B1(net2069));
 sg13g2_a22oi_1 _08022_ (.Y(_02916_),
    .B1(net2169),
    .B2(net2627),
    .A2(net2213),
    .A1(net2777));
 sg13g2_a22oi_1 _08023_ (.Y(_02917_),
    .B1(net2255),
    .B2(net1639),
    .A2(net2301),
    .A1(\rf_ram.RAM[15][4] ));
 sg13g2_a21oi_1 _08024_ (.A1(_02916_),
    .A2(_02917_),
    .Y(_02918_),
    .B1(net2104));
 sg13g2_a22oi_1 _08025_ (.Y(_02919_),
    .B1(net2171),
    .B2(\rf_ram.RAM[26][4] ),
    .A2(net2215),
    .A1(\rf_ram.RAM[25][4] ));
 sg13g2_a22oi_1 _08026_ (.Y(_02920_),
    .B1(net2257),
    .B2(net2658),
    .A2(net2303),
    .A1(net2961));
 sg13g2_a21oi_1 _08027_ (.A1(_02919_),
    .A2(_02920_),
    .Y(_02921_),
    .B1(net2085));
 sg13g2_a22oi_1 _08028_ (.Y(_02922_),
    .B1(net2169),
    .B2(net2836),
    .A2(net2213),
    .A1(net2663));
 sg13g2_a22oi_1 _08029_ (.Y(_02923_),
    .B1(net2255),
    .B2(net1482),
    .A2(net2297),
    .A1(net3785));
 sg13g2_a21oi_1 _08030_ (.A1(_02922_),
    .A2(_02923_),
    .Y(_02924_),
    .B1(net2310));
 sg13g2_a22oi_1 _08031_ (.Y(_02925_),
    .B1(net2170),
    .B2(net2742),
    .A2(net2214),
    .A1(net2772));
 sg13g2_a22oi_1 _08032_ (.Y(_02926_),
    .B1(net2256),
    .B2(net2969),
    .A2(net2302),
    .A1(net1551));
 sg13g2_a21oi_1 _08033_ (.A1(_02925_),
    .A2(_02926_),
    .Y(_02927_),
    .B1(net2075));
 sg13g2_a22oi_1 _08034_ (.Y(_02928_),
    .B1(net2170),
    .B2(net2770),
    .A2(net2214),
    .A1(net1479));
 sg13g2_a22oi_1 _08035_ (.Y(_02929_),
    .B1(net2257),
    .B2(net2936),
    .A2(net2303),
    .A1(net2766));
 sg13g2_a21oi_1 _08036_ (.A1(_02928_),
    .A2(_02929_),
    .Y(_02930_),
    .B1(net2080));
 sg13g2_a22oi_1 _08037_ (.Y(_02931_),
    .B1(net2171),
    .B2(net2613),
    .A2(net2215),
    .A1(net1480));
 sg13g2_a22oi_1 _08038_ (.Y(_02932_),
    .B1(net2256),
    .B2(net1428),
    .A2(net2302),
    .A1(net2672));
 sg13g2_a21oi_1 _08039_ (.A1(_02931_),
    .A2(_02932_),
    .Y(_02933_),
    .B1(net2262));
 sg13g2_a22oi_1 _08040_ (.Y(_02934_),
    .B1(net2169),
    .B2(net1600),
    .A2(net2213),
    .A1(net2739));
 sg13g2_a22oi_1 _08041_ (.Y(_02935_),
    .B1(net2255),
    .B2(net1718),
    .A2(net2301),
    .A1(net2888));
 sg13g2_a21oi_1 _08042_ (.A1(_02934_),
    .A2(_02935_),
    .Y(_02936_),
    .B1(net2099));
 sg13g2_nor4_1 _08043_ (.A(_02921_),
    .B(_02927_),
    .C(_02930_),
    .D(_02933_),
    .Y(_02937_));
 sg13g2_nor4_1 _08044_ (.A(_02915_),
    .B(_02918_),
    .C(_02924_),
    .D(_02936_),
    .Y(_02938_));
 sg13g2_a21oi_1 _08045_ (.A1(_02937_),
    .A2(net3786),
    .Y(_00437_),
    .B1(net2386));
 sg13g2_a22oi_1 _08046_ (.Y(_02939_),
    .B1(net2170),
    .B2(\rf_ram.RAM[18][5] ),
    .A2(net2214),
    .A1(\rf_ram.RAM[17][5] ));
 sg13g2_a22oi_1 _08047_ (.Y(_02940_),
    .B1(net2256),
    .B2(\rf_ram.RAM[16][5] ),
    .A2(net2302),
    .A1(\rf_ram.RAM[19][5] ));
 sg13g2_a21oi_1 _08048_ (.A1(_02939_),
    .A2(_02940_),
    .Y(_02941_),
    .B1(net2075));
 sg13g2_a22oi_1 _08049_ (.Y(_02942_),
    .B1(net2170),
    .B2(net1658),
    .A2(net2214),
    .A1(net3028));
 sg13g2_a22oi_1 _08050_ (.Y(_02943_),
    .B1(net2256),
    .B2(net2861),
    .A2(net2302),
    .A1(net3798));
 sg13g2_a21oi_1 _08051_ (.A1(_02942_),
    .A2(_02943_),
    .Y(_02944_),
    .B1(net2104));
 sg13g2_a22oi_1 _08052_ (.Y(_02945_),
    .B1(net2169),
    .B2(net2642),
    .A2(net2213),
    .A1(net1546));
 sg13g2_a22oi_1 _08053_ (.Y(_02946_),
    .B1(net2255),
    .B2(net1649),
    .A2(net2301),
    .A1(net1591));
 sg13g2_a21oi_1 _08054_ (.A1(_02945_),
    .A2(_02946_),
    .Y(_02947_),
    .B1(net2099));
 sg13g2_a22oi_1 _08055_ (.Y(_02948_),
    .B1(net2170),
    .B2(net3329),
    .A2(net2214),
    .A1(\rf_ram.RAM[25][5] ));
 sg13g2_a22oi_1 _08056_ (.Y(_02949_),
    .B1(net2256),
    .B2(net2992),
    .A2(net2302),
    .A1(\rf_ram.RAM[27][5] ));
 sg13g2_a21oi_1 _08057_ (.A1(_02948_),
    .A2(_02949_),
    .Y(_02950_),
    .B1(net2085));
 sg13g2_a22oi_1 _08058_ (.Y(_02951_),
    .B1(net2171),
    .B2(net2610),
    .A2(net2215),
    .A1(net1713));
 sg13g2_a22oi_1 _08059_ (.Y(_02952_),
    .B1(net2257),
    .B2(net2625),
    .A2(net2301),
    .A1(net2667));
 sg13g2_a21oi_1 _08060_ (.A1(_02951_),
    .A2(_02952_),
    .Y(_02953_),
    .B1(net2310));
 sg13g2_a22oi_1 _08061_ (.Y(_02954_),
    .B1(net2170),
    .B2(\rf_ram.RAM[30][5] ),
    .A2(net2214),
    .A1(\rf_ram.RAM[29][5] ));
 sg13g2_a22oi_1 _08062_ (.Y(_02955_),
    .B1(net2256),
    .B2(\rf_ram.RAM[28][5] ),
    .A2(net2302),
    .A1(\rf_ram.RAM[31][5] ));
 sg13g2_a21oi_1 _08063_ (.A1(_02954_),
    .A2(_02955_),
    .Y(_02956_),
    .B1(net2080));
 sg13g2_a22oi_1 _08064_ (.Y(_02957_),
    .B1(net2170),
    .B2(net2877),
    .A2(net2214),
    .A1(net1515));
 sg13g2_a22oi_1 _08065_ (.Y(_02958_),
    .B1(net2256),
    .B2(net1651),
    .A2(net2302),
    .A1(net2781));
 sg13g2_a21oi_1 _08066_ (.A1(_02957_),
    .A2(_02958_),
    .Y(_02959_),
    .B1(net2262));
 sg13g2_a22oi_1 _08067_ (.Y(_02960_),
    .B1(net2170),
    .B2(net1726),
    .A2(net2214),
    .A1(net3067));
 sg13g2_a22oi_1 _08068_ (.Y(_02961_),
    .B1(net2256),
    .B2(net2788),
    .A2(net2302),
    .A1(\rf_ram.RAM[23][5] ));
 sg13g2_a21oi_1 _08069_ (.A1(_02960_),
    .A2(_02961_),
    .Y(_02962_),
    .B1(net2069));
 sg13g2_nor4_1 _08070_ (.A(_02941_),
    .B(_02947_),
    .C(_02953_),
    .D(_02959_),
    .Y(_02963_));
 sg13g2_nor4_1 _08071_ (.A(_02944_),
    .B(_02950_),
    .C(_02956_),
    .D(_02962_),
    .Y(_02964_));
 sg13g2_a21oi_1 _08072_ (.A1(_02963_),
    .A2(net3799),
    .Y(_00438_),
    .B1(net2388));
 sg13g2_a22oi_1 _08073_ (.Y(_02965_),
    .B1(net2172),
    .B2(net1430),
    .A2(net2216),
    .A1(net2812));
 sg13g2_a22oi_1 _08074_ (.Y(_02966_),
    .B1(net2254),
    .B2(net3054),
    .A2(net2300),
    .A1(net2851));
 sg13g2_a21oi_1 _08075_ (.A1(_02965_),
    .A2(_02966_),
    .Y(_02967_),
    .B1(net2069));
 sg13g2_a22oi_1 _08076_ (.Y(_02968_),
    .B1(net2167),
    .B2(net1504),
    .A2(net2211),
    .A1(net1601));
 sg13g2_a22oi_1 _08077_ (.Y(_02969_),
    .B1(net2253),
    .B2(net1739),
    .A2(net2299),
    .A1(net2699));
 sg13g2_a21oi_1 _08078_ (.A1(_02968_),
    .A2(_02969_),
    .Y(_02970_),
    .B1(net2080));
 sg13g2_a22oi_1 _08079_ (.Y(_02971_),
    .B1(net2168),
    .B2(net1661),
    .A2(net2212),
    .A1(net2682));
 sg13g2_a22oi_1 _08080_ (.Y(_02972_),
    .B1(net2254),
    .B2(net1463),
    .A2(net2300),
    .A1(net1719));
 sg13g2_a21oi_1 _08081_ (.A1(_02971_),
    .A2(_02972_),
    .Y(_02973_),
    .B1(net2310));
 sg13g2_a22oi_1 _08082_ (.Y(_02974_),
    .B1(net2172),
    .B2(net3226),
    .A2(net2216),
    .A1(net2890));
 sg13g2_a22oi_1 _08083_ (.Y(_02975_),
    .B1(net2253),
    .B2(net2697),
    .A2(net2304),
    .A1(net3770));
 sg13g2_a21oi_1 _08084_ (.A1(_02974_),
    .A2(_02975_),
    .Y(_02976_),
    .B1(net2075));
 sg13g2_a22oi_1 _08085_ (.Y(_02977_),
    .B1(net2168),
    .B2(net1519),
    .A2(net2212),
    .A1(net1529));
 sg13g2_a22oi_1 _08086_ (.Y(_02978_),
    .B1(net2254),
    .B2(net1684),
    .A2(net2300),
    .A1(net1506));
 sg13g2_a21oi_1 _08087_ (.A1(_02977_),
    .A2(_02978_),
    .Y(_02979_),
    .B1(net2099));
 sg13g2_a22oi_1 _08088_ (.Y(_02980_),
    .B1(net2168),
    .B2(net2693),
    .A2(net2212),
    .A1(net1637));
 sg13g2_a22oi_1 _08089_ (.Y(_02981_),
    .B1(net2254),
    .B2(net2874),
    .A2(net2300),
    .A1(net2988));
 sg13g2_a21oi_1 _08090_ (.A1(_02980_),
    .A2(_02981_),
    .Y(_02982_),
    .B1(net2085));
 sg13g2_a22oi_1 _08091_ (.Y(_02983_),
    .B1(net2167),
    .B2(net2762),
    .A2(net2211),
    .A1(net2717));
 sg13g2_a22oi_1 _08092_ (.Y(_02984_),
    .B1(net2253),
    .B2(net3169),
    .A2(net2299),
    .A1(net1513));
 sg13g2_a21oi_1 _08093_ (.A1(_02983_),
    .A2(_02984_),
    .Y(_02985_),
    .B1(net2262));
 sg13g2_a22oi_1 _08094_ (.Y(_02986_),
    .B1(net2167),
    .B2(net2696),
    .A2(net2211),
    .A1(net1681));
 sg13g2_a22oi_1 _08095_ (.Y(_02987_),
    .B1(net2258),
    .B2(net2605),
    .A2(net2299),
    .A1(net3221));
 sg13g2_a21oi_1 _08096_ (.A1(_02986_),
    .A2(_02987_),
    .Y(_02988_),
    .B1(net2104));
 sg13g2_nor4_1 _08097_ (.A(_02967_),
    .B(_02973_),
    .C(_02979_),
    .D(_02982_),
    .Y(_02989_));
 sg13g2_nor4_1 _08098_ (.A(_02970_),
    .B(_02976_),
    .C(_02985_),
    .D(_02988_),
    .Y(_02990_));
 sg13g2_a21oi_1 _08099_ (.A1(_02989_),
    .A2(_02990_),
    .Y(_00439_),
    .B1(net2388));
 sg13g2_a22oi_1 _08100_ (.Y(_02991_),
    .B1(net2168),
    .B2(net3132),
    .A2(net2212),
    .A1(net2965));
 sg13g2_a22oi_1 _08101_ (.Y(_02992_),
    .B1(net2254),
    .B2(net3146),
    .A2(net2300),
    .A1(net2982));
 sg13g2_a21oi_1 _08102_ (.A1(_02991_),
    .A2(_02992_),
    .Y(_02993_),
    .B1(net2264));
 sg13g2_a22oi_1 _08103_ (.Y(_02994_),
    .B1(net2167),
    .B2(\rf_ram.RAM[18][7] ),
    .A2(net2211),
    .A1(\rf_ram.RAM[17][7] ));
 sg13g2_a22oi_1 _08104_ (.Y(_02995_),
    .B1(net2253),
    .B2(\rf_ram.RAM[16][7] ),
    .A2(net2299),
    .A1(\rf_ram.RAM[19][7] ));
 sg13g2_a21oi_1 _08105_ (.A1(_02994_),
    .A2(_02995_),
    .Y(_02996_),
    .B1(net2075));
 sg13g2_a22oi_1 _08106_ (.Y(_02997_),
    .B1(net2167),
    .B2(net3274),
    .A2(net2211),
    .A1(net2622));
 sg13g2_a22oi_1 _08107_ (.Y(_02998_),
    .B1(net2253),
    .B2(net3075),
    .A2(net2299),
    .A1(net2686));
 sg13g2_a21oi_1 _08108_ (.A1(_02997_),
    .A2(_02998_),
    .Y(_02999_),
    .B1(net2106));
 sg13g2_a22oi_1 _08109_ (.Y(_03000_),
    .B1(net2167),
    .B2(net1621),
    .A2(net2211),
    .A1(net1646));
 sg13g2_a22oi_1 _08110_ (.Y(_03001_),
    .B1(net2253),
    .B2(net2666),
    .A2(net2299),
    .A1(net3779));
 sg13g2_a21oi_1 _08111_ (.A1(_03000_),
    .A2(_03001_),
    .Y(_03002_),
    .B1(net2086));
 sg13g2_a22oi_1 _08112_ (.Y(_03003_),
    .B1(net2168),
    .B2(net3293),
    .A2(net2212),
    .A1(net3180));
 sg13g2_a22oi_1 _08113_ (.Y(_03004_),
    .B1(net2254),
    .B2(net2845),
    .A2(net2300),
    .A1(net1502));
 sg13g2_a21oi_1 _08114_ (.A1(_03003_),
    .A2(_03004_),
    .Y(_03005_),
    .B1(net2311));
 sg13g2_a22oi_1 _08115_ (.Y(_03006_),
    .B1(net2167),
    .B2(net2795),
    .A2(net2211),
    .A1(\rf_ram.RAM[29][7] ));
 sg13g2_a22oi_1 _08116_ (.Y(_03007_),
    .B1(net2253),
    .B2(net1424),
    .A2(net2299),
    .A1(\rf_ram.RAM[31][7] ));
 sg13g2_a21oi_1 _08117_ (.A1(_03006_),
    .A2(_03007_),
    .Y(_03008_),
    .B1(net2080));
 sg13g2_a22oi_1 _08118_ (.Y(_03009_),
    .B1(net2168),
    .B2(net2837),
    .A2(net2212),
    .A1(net2819));
 sg13g2_a22oi_1 _08119_ (.Y(_03010_),
    .B1(net2254),
    .B2(net2867),
    .A2(net2300),
    .A1(net1525));
 sg13g2_a21oi_1 _08120_ (.A1(_03009_),
    .A2(_03010_),
    .Y(_03011_),
    .B1(net2099));
 sg13g2_a22oi_1 _08121_ (.Y(_03012_),
    .B1(net2167),
    .B2(net2763),
    .A2(net2211),
    .A1(net2704));
 sg13g2_a22oi_1 _08122_ (.Y(_03013_),
    .B1(net2253),
    .B2(net2822),
    .A2(net2299),
    .A1(net3257));
 sg13g2_a21oi_1 _08123_ (.A1(_03012_),
    .A2(_03013_),
    .Y(_03014_),
    .B1(net2071));
 sg13g2_nor4_1 _08124_ (.A(_02993_),
    .B(_02996_),
    .C(_03005_),
    .D(_03011_),
    .Y(_03015_));
 sg13g2_nor4_1 _08125_ (.A(_02999_),
    .B(_03002_),
    .C(_03008_),
    .D(_03014_),
    .Y(_03016_));
 sg13g2_a21oi_1 _08126_ (.A1(_03015_),
    .A2(net3780),
    .Y(_00440_),
    .B1(net2388));
 sg13g2_a22oi_1 _08127_ (.Y(_03017_),
    .B1(net2159),
    .B2(net3344),
    .A2(net2203),
    .A1(net3387));
 sg13g2_a22oi_1 _08128_ (.Y(_03018_),
    .B1(net2245),
    .B2(net1488),
    .A2(net2291),
    .A1(net3187));
 sg13g2_a21oi_1 _08129_ (.A1(_03017_),
    .A2(_03018_),
    .Y(_03019_),
    .B1(net2070));
 sg13g2_a22oi_1 _08130_ (.Y(_03020_),
    .B1(net2159),
    .B2(net2846),
    .A2(net2203),
    .A1(net3069));
 sg13g2_a22oi_1 _08131_ (.Y(_03021_),
    .B1(net2245),
    .B2(net2953),
    .A2(net2291),
    .A1(net3774));
 sg13g2_a21oi_1 _08132_ (.A1(_03020_),
    .A2(_03021_),
    .Y(_03022_),
    .B1(net2263));
 sg13g2_a22oi_1 _08133_ (.Y(_03023_),
    .B1(net2159),
    .B2(net1433),
    .A2(net2203),
    .A1(net1657));
 sg13g2_a22oi_1 _08134_ (.Y(_03024_),
    .B1(net2246),
    .B2(net1746),
    .A2(net2292),
    .A1(net2930));
 sg13g2_a21oi_1 _08135_ (.A1(_03023_),
    .A2(_03024_),
    .Y(_03025_),
    .B1(net2074));
 sg13g2_a22oi_1 _08136_ (.Y(_03026_),
    .B1(net2160),
    .B2(net3043),
    .A2(net2204),
    .A1(net2881));
 sg13g2_a22oi_1 _08137_ (.Y(_03027_),
    .B1(net2246),
    .B2(net2794),
    .A2(net2292),
    .A1(net2775));
 sg13g2_a21oi_1 _08138_ (.A1(_03026_),
    .A2(_03027_),
    .Y(_03028_),
    .B1(net2100));
 sg13g2_a22oi_1 _08139_ (.Y(_03029_),
    .B1(net2160),
    .B2(net1612),
    .A2(net2204),
    .A1(net2644));
 sg13g2_a22oi_1 _08140_ (.Y(_03030_),
    .B1(net2246),
    .B2(net1656),
    .A2(net2292),
    .A1(net2949));
 sg13g2_a21oi_1 _08141_ (.A1(_03029_),
    .A2(_03030_),
    .Y(_03031_),
    .B1(net2309));
 sg13g2_a22oi_1 _08142_ (.Y(_03032_),
    .B1(net2159),
    .B2(net1484),
    .A2(net2203),
    .A1(net2853));
 sg13g2_a22oi_1 _08143_ (.Y(_03033_),
    .B1(net2245),
    .B2(net3203),
    .A2(net2291),
    .A1(net2880));
 sg13g2_a21oi_1 _08144_ (.A1(_03032_),
    .A2(_03033_),
    .Y(_03034_),
    .B1(net2079));
 sg13g2_a22oi_1 _08145_ (.Y(_03035_),
    .B1(net2160),
    .B2(net2955),
    .A2(net2204),
    .A1(net2866));
 sg13g2_a22oi_1 _08146_ (.Y(_03036_),
    .B1(net2246),
    .B2(net1495),
    .A2(net2292),
    .A1(net3099));
 sg13g2_a21oi_1 _08147_ (.A1(_03035_),
    .A2(_03036_),
    .Y(_03037_),
    .B1(net2105));
 sg13g2_a22oi_1 _08148_ (.Y(_03038_),
    .B1(net2160),
    .B2(net3061),
    .A2(net2204),
    .A1(net1453));
 sg13g2_a22oi_1 _08149_ (.Y(_03039_),
    .B1(net2246),
    .B2(net2637),
    .A2(net2292),
    .A1(net3122));
 sg13g2_a21oi_1 _08150_ (.A1(_03038_),
    .A2(_03039_),
    .Y(_03040_),
    .B1(net2085));
 sg13g2_nor4_1 _08151_ (.A(_03019_),
    .B(_03025_),
    .C(_03031_),
    .D(_03034_),
    .Y(_03041_));
 sg13g2_nor4_1 _08152_ (.A(_03022_),
    .B(_03028_),
    .C(_03037_),
    .D(_03040_),
    .Y(_03042_));
 sg13g2_a21oi_1 _08153_ (.A1(_03041_),
    .A2(_03042_),
    .Y(_00441_),
    .B1(net2386));
 sg13g2_a22oi_1 _08154_ (.Y(_03043_),
    .B1(net2156),
    .B2(\rf_ram.RAM[6][9] ),
    .A2(net2200),
    .A1(\rf_ram.RAM[5][9] ));
 sg13g2_a22oi_1 _08155_ (.Y(_03044_),
    .B1(net2243),
    .B2(\rf_ram.RAM[4][9] ),
    .A2(net2289),
    .A1(\rf_ram.RAM[7][9] ));
 sg13g2_a21oi_1 _08156_ (.A1(_03043_),
    .A2(_03044_),
    .Y(_03045_),
    .B1(net2263));
 sg13g2_a22oi_1 _08157_ (.Y(_03046_),
    .B1(net2157),
    .B2(net2960),
    .A2(net2201),
    .A1(\rf_ram.RAM[25][9] ));
 sg13g2_a22oi_1 _08158_ (.Y(_03047_),
    .B1(net2244),
    .B2(net3042),
    .A2(net2290),
    .A1(\rf_ram.RAM[27][9] ));
 sg13g2_a21oi_1 _08159_ (.A1(_03046_),
    .A2(_03047_),
    .Y(_03048_),
    .B1(net2084));
 sg13g2_a22oi_1 _08160_ (.Y(_03049_),
    .B1(net2156),
    .B2(\rf_ram.RAM[30][9] ),
    .A2(net2200),
    .A1(\rf_ram.RAM[29][9] ));
 sg13g2_a22oi_1 _08161_ (.Y(_03050_),
    .B1(net2243),
    .B2(\rf_ram.RAM[28][9] ),
    .A2(net2289),
    .A1(\rf_ram.RAM[31][9] ));
 sg13g2_a21oi_1 _08162_ (.A1(_03049_),
    .A2(_03050_),
    .Y(_03051_),
    .B1(net2079));
 sg13g2_a22oi_1 _08163_ (.Y(_03052_),
    .B1(net2157),
    .B2(net1490),
    .A2(net2201),
    .A1(net3800));
 sg13g2_a22oi_1 _08164_ (.Y(_03053_),
    .B1(net2244),
    .B2(net2998),
    .A2(net2290),
    .A1(\rf_ram.RAM[11][9] ));
 sg13g2_a21oi_1 _08165_ (.A1(_03052_),
    .A2(_03053_),
    .Y(_03054_),
    .B1(net2100));
 sg13g2_a22oi_1 _08166_ (.Y(_03055_),
    .B1(net2156),
    .B2(\rf_ram.RAM[18][9] ),
    .A2(net2200),
    .A1(\rf_ram.RAM[17][9] ));
 sg13g2_a22oi_1 _08167_ (.Y(_03056_),
    .B1(net2243),
    .B2(\rf_ram.RAM[16][9] ),
    .A2(net2289),
    .A1(\rf_ram.RAM[19][9] ));
 sg13g2_a21oi_1 _08168_ (.A1(_03055_),
    .A2(_03056_),
    .Y(_03057_),
    .B1(net2074));
 sg13g2_a22oi_1 _08169_ (.Y(_03058_),
    .B1(net2157),
    .B2(net2629),
    .A2(net2201),
    .A1(\rf_ram.RAM[1][9] ));
 sg13g2_a22oi_1 _08170_ (.Y(_03059_),
    .B1(net2244),
    .B2(\rf_ram.RAM[0][9] ),
    .A2(net2290),
    .A1(\rf_ram.RAM[3][9] ));
 sg13g2_a21oi_1 _08171_ (.A1(_03058_),
    .A2(_03059_),
    .Y(_03060_),
    .B1(net2309));
 sg13g2_a22oi_1 _08172_ (.Y(_03061_),
    .B1(net2156),
    .B2(\rf_ram.RAM[14][9] ),
    .A2(net2200),
    .A1(\rf_ram.RAM[13][9] ));
 sg13g2_a22oi_1 _08173_ (.Y(_03062_),
    .B1(net2243),
    .B2(\rf_ram.RAM[12][9] ),
    .A2(net2289),
    .A1(\rf_ram.RAM[15][9] ));
 sg13g2_a21oi_1 _08174_ (.A1(_03061_),
    .A2(_03062_),
    .Y(_03063_),
    .B1(net2105));
 sg13g2_a22oi_1 _08175_ (.Y(_03064_),
    .B1(net2157),
    .B2(net1692),
    .A2(net2201),
    .A1(net3108));
 sg13g2_a22oi_1 _08176_ (.Y(_03065_),
    .B1(net2244),
    .B2(net1472),
    .A2(net2290),
    .A1(\rf_ram.RAM[23][9] ));
 sg13g2_a21oi_1 _08177_ (.A1(_03064_),
    .A2(_03065_),
    .Y(_03066_),
    .B1(net2070));
 sg13g2_nor4_1 _08178_ (.A(_03045_),
    .B(_03051_),
    .C(_03057_),
    .D(_03063_),
    .Y(_03067_));
 sg13g2_nor4_1 _08179_ (.A(_03048_),
    .B(_03054_),
    .C(_03060_),
    .D(_03066_),
    .Y(_03068_));
 sg13g2_a21oi_1 _08180_ (.A1(_03067_),
    .A2(net3801),
    .Y(_00442_),
    .B1(net2386));
 sg13g2_a22oi_1 _08181_ (.Y(_03069_),
    .B1(net2159),
    .B2(net2714),
    .A2(net2203),
    .A1(net3215));
 sg13g2_a22oi_1 _08182_ (.Y(_03070_),
    .B1(net2245),
    .B2(net1733),
    .A2(net2291),
    .A1(net1633));
 sg13g2_a21oi_1 _08183_ (.A1(_03069_),
    .A2(_03070_),
    .Y(_03071_),
    .B1(net2105));
 sg13g2_a22oi_1 _08184_ (.Y(_03072_),
    .B1(net2159),
    .B2(net2973),
    .A2(net2203),
    .A1(net2677));
 sg13g2_a22oi_1 _08185_ (.Y(_03073_),
    .B1(net2245),
    .B2(net3285),
    .A2(net2291),
    .A1(net3320));
 sg13g2_a21oi_1 _08186_ (.A1(_03072_),
    .A2(_03073_),
    .Y(_03074_),
    .B1(net2084));
 sg13g2_a22oi_1 _08187_ (.Y(_03075_),
    .B1(net2159),
    .B2(net2945),
    .A2(net2203),
    .A1(net3149));
 sg13g2_a22oi_1 _08188_ (.Y(_03076_),
    .B1(net2245),
    .B2(net3256),
    .A2(net2291),
    .A1(net1682));
 sg13g2_a21oi_1 _08189_ (.A1(_03075_),
    .A2(_03076_),
    .Y(_03077_),
    .B1(net2070));
 sg13g2_a22oi_1 _08190_ (.Y(_03078_),
    .B1(net2160),
    .B2(net1441),
    .A2(net2204),
    .A1(\rf_ram.RAM[9][10] ));
 sg13g2_a22oi_1 _08191_ (.Y(_03079_),
    .B1(net2246),
    .B2(\rf_ram.RAM[8][10] ),
    .A2(net2292),
    .A1(\rf_ram.RAM[11][10] ));
 sg13g2_a21oi_1 _08192_ (.A1(_03078_),
    .A2(_03079_),
    .Y(_03080_),
    .B1(net2100));
 sg13g2_a22oi_1 _08193_ (.Y(_03081_),
    .B1(net2159),
    .B2(net1462),
    .A2(net2203),
    .A1(net1687));
 sg13g2_a22oi_1 _08194_ (.Y(_03082_),
    .B1(net2245),
    .B2(net2896),
    .A2(net2291),
    .A1(net1647));
 sg13g2_a21oi_1 _08195_ (.A1(_03081_),
    .A2(_03082_),
    .Y(_03083_),
    .B1(net2074));
 sg13g2_a22oi_1 _08196_ (.Y(_03084_),
    .B1(net2156),
    .B2(net2751),
    .A2(net2200),
    .A1(net2991));
 sg13g2_a22oi_1 _08197_ (.Y(_03085_),
    .B1(net2245),
    .B2(net2959),
    .A2(net2291),
    .A1(\rf_ram.RAM[31][10] ));
 sg13g2_a21oi_1 _08198_ (.A1(_03084_),
    .A2(_03085_),
    .Y(_03086_),
    .B1(net2079));
 sg13g2_a22oi_1 _08199_ (.Y(_03087_),
    .B1(net2157),
    .B2(net1501),
    .A2(net2201),
    .A1(net3196));
 sg13g2_a22oi_1 _08200_ (.Y(_03088_),
    .B1(net2244),
    .B2(net1550),
    .A2(net2290),
    .A1(net1468));
 sg13g2_a21oi_1 _08201_ (.A1(_03087_),
    .A2(_03088_),
    .Y(_03089_),
    .B1(net2309));
 sg13g2_a22oi_1 _08202_ (.Y(_03090_),
    .B1(net2158),
    .B2(net2701),
    .A2(net2202),
    .A1(net1560));
 sg13g2_a22oi_1 _08203_ (.Y(_03091_),
    .B1(net2243),
    .B2(net2942),
    .A2(net2289),
    .A1(net3777));
 sg13g2_a21oi_1 _08204_ (.A1(_03090_),
    .A2(_03091_),
    .Y(_03092_),
    .B1(net2263));
 sg13g2_nor4_1 _08205_ (.A(_03071_),
    .B(_03077_),
    .C(_03083_),
    .D(_03089_),
    .Y(_03093_));
 sg13g2_nor4_1 _08206_ (.A(_03074_),
    .B(_03080_),
    .C(_03086_),
    .D(_03092_),
    .Y(_03094_));
 sg13g2_a21oi_1 _08207_ (.A1(_03093_),
    .A2(net3778),
    .Y(_00443_),
    .B1(net2386));
 sg13g2_a22oi_1 _08208_ (.Y(_03095_),
    .B1(net2155),
    .B2(net3267),
    .A2(net2199),
    .A1(net2987));
 sg13g2_a22oi_1 _08209_ (.Y(_03096_),
    .B1(net2242),
    .B2(net1660),
    .A2(net2285),
    .A1(net2635));
 sg13g2_a21oi_1 _08210_ (.A1(_03095_),
    .A2(_03096_),
    .Y(_03097_),
    .B1(net2084));
 sg13g2_a22oi_1 _08211_ (.Y(_03098_),
    .B1(net2152),
    .B2(net2878),
    .A2(net2196),
    .A1(net1492));
 sg13g2_a22oi_1 _08212_ (.Y(_03099_),
    .B1(net2239),
    .B2(net1635),
    .A2(net2285),
    .A1(net1712));
 sg13g2_a21oi_1 _08213_ (.A1(_03098_),
    .A2(_03099_),
    .Y(_03100_),
    .B1(net2079));
 sg13g2_a22oi_1 _08214_ (.Y(_03101_),
    .B1(net2152),
    .B2(net3250),
    .A2(net2196),
    .A1(net3109));
 sg13g2_a22oi_1 _08215_ (.Y(_03102_),
    .B1(net2239),
    .B2(net3170),
    .A2(net2285),
    .A1(net2744));
 sg13g2_a21oi_1 _08216_ (.A1(_03101_),
    .A2(_03102_),
    .Y(_03103_),
    .B1(net2309));
 sg13g2_a22oi_1 _08217_ (.Y(_03104_),
    .B1(net2152),
    .B2(net3040),
    .A2(net2196),
    .A1(net3063));
 sg13g2_a22oi_1 _08218_ (.Y(_03105_),
    .B1(net2239),
    .B2(net1485),
    .A2(net2285),
    .A1(net2747));
 sg13g2_a21oi_1 _08219_ (.A1(_03104_),
    .A2(_03105_),
    .Y(_03106_),
    .B1(net2070));
 sg13g2_a22oi_1 _08220_ (.Y(_03107_),
    .B1(net2152),
    .B2(net1645),
    .A2(net2196),
    .A1(net3290));
 sg13g2_a22oi_1 _08221_ (.Y(_03108_),
    .B1(net2239),
    .B2(net1483),
    .A2(net2288),
    .A1(net3047));
 sg13g2_a21oi_1 _08222_ (.A1(_03107_),
    .A2(_03108_),
    .Y(_03109_),
    .B1(net2105));
 sg13g2_a22oi_1 _08223_ (.Y(_03110_),
    .B1(net2152),
    .B2(net2647),
    .A2(net2196),
    .A1(net2927));
 sg13g2_a22oi_1 _08224_ (.Y(_03111_),
    .B1(net2239),
    .B2(net3044),
    .A2(net2285),
    .A1(net2858));
 sg13g2_a21oi_1 _08225_ (.A1(_03110_),
    .A2(_03111_),
    .Y(_03112_),
    .B1(net2263));
 sg13g2_a22oi_1 _08226_ (.Y(_03113_),
    .B1(net2152),
    .B2(net1454),
    .A2(net2196),
    .A1(net2948));
 sg13g2_a22oi_1 _08227_ (.Y(_03114_),
    .B1(net2239),
    .B2(net2947),
    .A2(net2285),
    .A1(net1693));
 sg13g2_a21oi_1 _08228_ (.A1(_03113_),
    .A2(_03114_),
    .Y(_03115_),
    .B1(net2074));
 sg13g2_a22oi_1 _08229_ (.Y(_03116_),
    .B1(net2152),
    .B2(net3056),
    .A2(net2196),
    .A1(net3276));
 sg13g2_a22oi_1 _08230_ (.Y(_03117_),
    .B1(net2239),
    .B2(net1486),
    .A2(net2285),
    .A1(net3174));
 sg13g2_a21oi_1 _08231_ (.A1(_03116_),
    .A2(_03117_),
    .Y(_03118_),
    .B1(net2100));
 sg13g2_nor4_1 _08232_ (.A(_03097_),
    .B(_03103_),
    .C(_03109_),
    .D(_03115_),
    .Y(_03119_));
 sg13g2_nor4_1 _08233_ (.A(_03100_),
    .B(_03106_),
    .C(_03112_),
    .D(_03118_),
    .Y(_03120_));
 sg13g2_a21oi_1 _08234_ (.A1(_03119_),
    .A2(_03120_),
    .Y(_00444_),
    .B1(net2386));
 sg13g2_a22oi_1 _08235_ (.Y(_03121_),
    .B1(net2157),
    .B2(net3160),
    .A2(net2201),
    .A1(net1734));
 sg13g2_a22oi_1 _08236_ (.Y(_03122_),
    .B1(net2244),
    .B2(net2844),
    .A2(net2290),
    .A1(net3165));
 sg13g2_a21oi_1 _08237_ (.A1(_03121_),
    .A2(_03122_),
    .Y(_03123_),
    .B1(net2309));
 sg13g2_a22oi_1 _08238_ (.Y(_03124_),
    .B1(net2156),
    .B2(net1467),
    .A2(net2200),
    .A1(\rf_ram.RAM[17][12] ));
 sg13g2_a22oi_1 _08239_ (.Y(_03125_),
    .B1(net2243),
    .B2(\rf_ram.RAM[16][12] ),
    .A2(net2289),
    .A1(\rf_ram.RAM[19][12] ));
 sg13g2_a21oi_1 _08240_ (.A1(_03124_),
    .A2(_03125_),
    .Y(_03126_),
    .B1(net2074));
 sg13g2_a22oi_1 _08241_ (.Y(_03127_),
    .B1(net2158),
    .B2(net2833),
    .A2(net2202),
    .A1(net2761));
 sg13g2_a22oi_1 _08242_ (.Y(_03128_),
    .B1(net2247),
    .B2(net1680),
    .A2(net2293),
    .A1(net1475));
 sg13g2_a21oi_1 _08243_ (.A1(_03127_),
    .A2(_03128_),
    .Y(_03129_),
    .B1(net2105));
 sg13g2_a22oi_1 _08244_ (.Y(_03130_),
    .B1(net2157),
    .B2(net3186),
    .A2(net2201),
    .A1(net3318));
 sg13g2_a22oi_1 _08245_ (.Y(_03131_),
    .B1(net2244),
    .B2(net3308),
    .A2(net2290),
    .A1(net3377));
 sg13g2_a21oi_1 _08246_ (.A1(_03130_),
    .A2(_03131_),
    .Y(_03132_),
    .B1(net2263));
 sg13g2_a22oi_1 _08247_ (.Y(_03133_),
    .B1(net2158),
    .B2(net2671),
    .A2(net2202),
    .A1(net2924));
 sg13g2_a22oi_1 _08248_ (.Y(_03134_),
    .B1(net2247),
    .B2(net1427),
    .A2(net2293),
    .A1(net3233));
 sg13g2_a21oi_1 _08249_ (.A1(_03133_),
    .A2(_03134_),
    .Y(_03135_),
    .B1(net2070));
 sg13g2_a22oi_1 _08250_ (.Y(_03136_),
    .B1(net2156),
    .B2(net3192),
    .A2(net2200),
    .A1(net2809));
 sg13g2_a22oi_1 _08251_ (.Y(_03137_),
    .B1(net2243),
    .B2(net2798),
    .A2(net2289),
    .A1(net3139));
 sg13g2_a21oi_1 _08252_ (.A1(_03136_),
    .A2(_03137_),
    .Y(_03138_),
    .B1(net2079));
 sg13g2_a22oi_1 _08253_ (.Y(_03139_),
    .B1(net2156),
    .B2(net1528),
    .A2(net2200),
    .A1(net1717));
 sg13g2_a22oi_1 _08254_ (.Y(_03140_),
    .B1(net2243),
    .B2(net2954),
    .A2(net2289),
    .A1(net1474));
 sg13g2_a21oi_1 _08255_ (.A1(_03139_),
    .A2(_03140_),
    .Y(_03141_),
    .B1(net2084));
 sg13g2_a22oi_1 _08256_ (.Y(_03142_),
    .B1(net2157),
    .B2(net1559),
    .A2(net2201),
    .A1(net3168));
 sg13g2_a22oi_1 _08257_ (.Y(_03143_),
    .B1(net2244),
    .B2(net1420),
    .A2(net2290),
    .A1(net3771));
 sg13g2_a21oi_1 _08258_ (.A1(_03142_),
    .A2(_03143_),
    .Y(_03144_),
    .B1(net2100));
 sg13g2_nor4_1 _08259_ (.A(_03129_),
    .B(_03135_),
    .C(_03138_),
    .D(_03141_),
    .Y(_03145_));
 sg13g2_nor4_1 _08260_ (.A(_03123_),
    .B(_03126_),
    .C(_03132_),
    .D(_03144_),
    .Y(_03146_));
 sg13g2_a21oi_1 _08261_ (.A1(_03145_),
    .A2(net3772),
    .Y(_00445_),
    .B1(net2386));
 sg13g2_a22oi_1 _08262_ (.Y(_03147_),
    .B1(net2163),
    .B2(net3085),
    .A2(net2207),
    .A1(net1641));
 sg13g2_a22oi_1 _08263_ (.Y(_03148_),
    .B1(net2249),
    .B2(net3119),
    .A2(net2295),
    .A1(net2911));
 sg13g2_a21oi_1 _08264_ (.A1(_03147_),
    .A2(_03148_),
    .Y(_03149_),
    .B1(net2101));
 sg13g2_a22oi_1 _08265_ (.Y(_03150_),
    .B1(net2168),
    .B2(\rf_ram.RAM[30][13] ),
    .A2(net2212),
    .A1(\rf_ram.RAM[29][13] ));
 sg13g2_a22oi_1 _08266_ (.Y(_03151_),
    .B1(net2254),
    .B2(\rf_ram.RAM[28][13] ),
    .A2(net2300),
    .A1(\rf_ram.RAM[31][13] ));
 sg13g2_a21oi_1 _08267_ (.A1(_03150_),
    .A2(_03151_),
    .Y(_03152_),
    .B1(net2080));
 sg13g2_a22oi_1 _08268_ (.Y(_03153_),
    .B1(net2163),
    .B2(net1650),
    .A2(net2207),
    .A1(net2956));
 sg13g2_a22oi_1 _08269_ (.Y(_03154_),
    .B1(net2249),
    .B2(net3150),
    .A2(net2295),
    .A1(net3070));
 sg13g2_a21oi_1 _08270_ (.A1(_03153_),
    .A2(_03154_),
    .Y(_03155_),
    .B1(net2104));
 sg13g2_a22oi_1 _08271_ (.Y(_03156_),
    .B1(net2154),
    .B2(net2619),
    .A2(net2198),
    .A1(net3245));
 sg13g2_a22oi_1 _08272_ (.Y(_03157_),
    .B1(net2241),
    .B2(net3200),
    .A2(net2287),
    .A1(net3103));
 sg13g2_a21oi_1 _08273_ (.A1(_03156_),
    .A2(_03157_),
    .Y(_03158_),
    .B1(net2070));
 sg13g2_a22oi_1 _08274_ (.Y(_03159_),
    .B1(net2155),
    .B2(net3294),
    .A2(net2199),
    .A1(net1701));
 sg13g2_a22oi_1 _08275_ (.Y(_03160_),
    .B1(net2242),
    .B2(net1481),
    .A2(net2288),
    .A1(net2854));
 sg13g2_a21oi_1 _08276_ (.A1(_03159_),
    .A2(_03160_),
    .Y(_03161_),
    .B1(net2074));
 sg13g2_a22oi_1 _08277_ (.Y(_03162_),
    .B1(net2155),
    .B2(net1642),
    .A2(net2199),
    .A1(net3213));
 sg13g2_a22oi_1 _08278_ (.Y(_03163_),
    .B1(net2242),
    .B2(net3240),
    .A2(net2288),
    .A1(net3018));
 sg13g2_a21oi_1 _08279_ (.A1(_03162_),
    .A2(_03163_),
    .Y(_03164_),
    .B1(net2263));
 sg13g2_a22oi_1 _08280_ (.Y(_03165_),
    .B1(net2163),
    .B2(net1703),
    .A2(net2207),
    .A1(net3148));
 sg13g2_a22oi_1 _08281_ (.Y(_03166_),
    .B1(net2249),
    .B2(net3094),
    .A2(net2295),
    .A1(net3117));
 sg13g2_a21oi_1 _08282_ (.A1(_03165_),
    .A2(_03166_),
    .Y(_03167_),
    .B1(net2084));
 sg13g2_a22oi_1 _08283_ (.Y(_03168_),
    .B1(net2155),
    .B2(net1516),
    .A2(net2199),
    .A1(net2727));
 sg13g2_a22oi_1 _08284_ (.Y(_03169_),
    .B1(net2242),
    .B2(net2859),
    .A2(net2288),
    .A1(net1564));
 sg13g2_a21oi_1 _08285_ (.A1(_03168_),
    .A2(_03169_),
    .Y(_03170_),
    .B1(net2311));
 sg13g2_nor4_1 _08286_ (.A(_03149_),
    .B(_03152_),
    .C(_03155_),
    .D(_03167_),
    .Y(_03171_));
 sg13g2_nor4_1 _08287_ (.A(_03158_),
    .B(_03161_),
    .C(_03164_),
    .D(_03170_),
    .Y(_03172_));
 sg13g2_a21oi_1 _08288_ (.A1(_03171_),
    .A2(_03172_),
    .Y(_00446_),
    .B1(net2386));
 sg13g2_a22oi_1 _08289_ (.Y(_03173_),
    .B1(net2136),
    .B2(\rf_ram.RAM[10][14] ),
    .A2(net2180),
    .A1(\rf_ram.RAM[9][14] ));
 sg13g2_a22oi_1 _08290_ (.Y(_03174_),
    .B1(net2224),
    .B2(\rf_ram.RAM[8][14] ),
    .A2(net2271),
    .A1(\rf_ram.RAM[11][14] ));
 sg13g2_a21oi_1 _08291_ (.A1(_03173_),
    .A2(_03174_),
    .Y(_03175_),
    .B1(net2097));
 sg13g2_a22oi_1 _08292_ (.Y(_03176_),
    .B1(net2136),
    .B2(\rf_ram.RAM[14][14] ),
    .A2(net2180),
    .A1(\rf_ram.RAM[13][14] ));
 sg13g2_a22oi_1 _08293_ (.Y(_03177_),
    .B1(net2224),
    .B2(\rf_ram.RAM[12][14] ),
    .A2(net2272),
    .A1(\rf_ram.RAM[15][14] ));
 sg13g2_a21oi_1 _08294_ (.A1(_03176_),
    .A2(_03177_),
    .Y(_03178_),
    .B1(net2103));
 sg13g2_a22oi_1 _08295_ (.Y(_03179_),
    .B1(net2137),
    .B2(net3816),
    .A2(net2181),
    .A1(\rf_ram.RAM[21][14] ));
 sg13g2_a22oi_1 _08296_ (.Y(_03180_),
    .B1(net2225),
    .B2(\rf_ram.RAM[20][14] ),
    .A2(net2272),
    .A1(\rf_ram.RAM[23][14] ));
 sg13g2_a21oi_1 _08297_ (.A1(_03179_),
    .A2(_03180_),
    .Y(_03181_),
    .B1(net2067));
 sg13g2_a22oi_1 _08298_ (.Y(_03182_),
    .B1(net2137),
    .B2(\rf_ram.RAM[30][14] ),
    .A2(net2181),
    .A1(\rf_ram.RAM[29][14] ));
 sg13g2_a22oi_1 _08299_ (.Y(_03183_),
    .B1(net2224),
    .B2(\rf_ram.RAM[28][14] ),
    .A2(net2271),
    .A1(\rf_ram.RAM[31][14] ));
 sg13g2_a21oi_1 _08300_ (.A1(_03182_),
    .A2(_03183_),
    .Y(_03184_),
    .B1(net2077));
 sg13g2_a22oi_1 _08301_ (.Y(_03185_),
    .B1(net2137),
    .B2(\rf_ram.RAM[6][14] ),
    .A2(net2181),
    .A1(\rf_ram.RAM[5][14] ));
 sg13g2_a22oi_1 _08302_ (.Y(_03186_),
    .B1(net2225),
    .B2(\rf_ram.RAM[4][14] ),
    .A2(net2272),
    .A1(\rf_ram.RAM[7][14] ));
 sg13g2_a21oi_1 _08303_ (.A1(_03185_),
    .A2(_03186_),
    .Y(_03187_),
    .B1(net2261));
 sg13g2_a22oi_1 _08304_ (.Y(_03188_),
    .B1(net2136),
    .B2(\rf_ram.RAM[2][14] ),
    .A2(net2180),
    .A1(\rf_ram.RAM[1][14] ));
 sg13g2_a22oi_1 _08305_ (.Y(_03189_),
    .B1(net2224),
    .B2(\rf_ram.RAM[0][14] ),
    .A2(net2271),
    .A1(\rf_ram.RAM[3][14] ));
 sg13g2_a21oi_1 _08306_ (.A1(_03188_),
    .A2(_03189_),
    .Y(_03190_),
    .B1(net2308));
 sg13g2_a22oi_1 _08307_ (.Y(_03191_),
    .B1(net2136),
    .B2(\rf_ram.RAM[18][14] ),
    .A2(net2180),
    .A1(\rf_ram.RAM[17][14] ));
 sg13g2_a22oi_1 _08308_ (.Y(_03192_),
    .B1(net2224),
    .B2(\rf_ram.RAM[16][14] ),
    .A2(net2271),
    .A1(\rf_ram.RAM[19][14] ));
 sg13g2_a21oi_1 _08309_ (.A1(_03191_),
    .A2(_03192_),
    .Y(_03193_),
    .B1(net2072));
 sg13g2_a22oi_1 _08310_ (.Y(_03194_),
    .B1(net2136),
    .B2(\rf_ram.RAM[26][14] ),
    .A2(net2180),
    .A1(\rf_ram.RAM[25][14] ));
 sg13g2_a22oi_1 _08311_ (.Y(_03195_),
    .B1(net2224),
    .B2(\rf_ram.RAM[24][14] ),
    .A2(net2271),
    .A1(\rf_ram.RAM[27][14] ));
 sg13g2_a21oi_1 _08312_ (.A1(_03194_),
    .A2(_03195_),
    .Y(_03196_),
    .B1(net2082));
 sg13g2_nor4_1 _08313_ (.A(_03175_),
    .B(_03181_),
    .C(_03187_),
    .D(_03193_),
    .Y(_03197_));
 sg13g2_nor4_1 _08314_ (.A(_03178_),
    .B(_03184_),
    .C(_03190_),
    .D(_03196_),
    .Y(_03198_));
 sg13g2_a21oi_1 _08315_ (.A1(net3817),
    .A2(_03198_),
    .Y(_00447_),
    .B1(net2385));
 sg13g2_a22oi_1 _08316_ (.Y(_03199_),
    .B1(net2154),
    .B2(net1449),
    .A2(net2198),
    .A1(net1620));
 sg13g2_a22oi_1 _08317_ (.Y(_03200_),
    .B1(net2241),
    .B2(net3091),
    .A2(net2287),
    .A1(net2823));
 sg13g2_a21oi_1 _08318_ (.A1(_03199_),
    .A2(_03200_),
    .Y(_03201_),
    .B1(net2079));
 sg13g2_a22oi_1 _08319_ (.Y(_03202_),
    .B1(net2139),
    .B2(net3059),
    .A2(net2183),
    .A1(net3191));
 sg13g2_a22oi_1 _08320_ (.Y(_03203_),
    .B1(net2227),
    .B2(net3141),
    .A2(net2274),
    .A1(net2868));
 sg13g2_a21oi_1 _08321_ (.A1(_03202_),
    .A2(_03203_),
    .Y(_03204_),
    .B1(net2309));
 sg13g2_a22oi_1 _08322_ (.Y(_03205_),
    .B1(net2139),
    .B2(net2737),
    .A2(net2183),
    .A1(net2923));
 sg13g2_a22oi_1 _08323_ (.Y(_03206_),
    .B1(net2227),
    .B2(net3275),
    .A2(net2274),
    .A1(net3270));
 sg13g2_a21oi_1 _08324_ (.A1(_03205_),
    .A2(_03206_),
    .Y(_03207_),
    .B1(net2084));
 sg13g2_a22oi_1 _08325_ (.Y(_03208_),
    .B1(net2139),
    .B2(net1588),
    .A2(net2183),
    .A1(net1624));
 sg13g2_a22oi_1 _08326_ (.Y(_03209_),
    .B1(net2227),
    .B2(net1672),
    .A2(net2274),
    .A1(net3182));
 sg13g2_a21oi_1 _08327_ (.A1(_03208_),
    .A2(_03209_),
    .Y(_03210_),
    .B1(net2102));
 sg13g2_a22oi_1 _08328_ (.Y(_03211_),
    .B1(net2154),
    .B2(net1618),
    .A2(net2198),
    .A1(net3135));
 sg13g2_a22oi_1 _08329_ (.Y(_03212_),
    .B1(net2241),
    .B2(net2631),
    .A2(net2287),
    .A1(net1445));
 sg13g2_a21oi_1 _08330_ (.A1(_03211_),
    .A2(_03212_),
    .Y(_03213_),
    .B1(net2263));
 sg13g2_a22oi_1 _08331_ (.Y(_03214_),
    .B1(net2154),
    .B2(net2722),
    .A2(net2198),
    .A1(net2706));
 sg13g2_a22oi_1 _08332_ (.Y(_03215_),
    .B1(net2241),
    .B2(net3171),
    .A2(net2287),
    .A1(net2734));
 sg13g2_a21oi_1 _08333_ (.A1(_03214_),
    .A2(_03215_),
    .Y(_03216_),
    .B1(net2100));
 sg13g2_a22oi_1 _08334_ (.Y(_03217_),
    .B1(net2154),
    .B2(net2645),
    .A2(net2198),
    .A1(net3307));
 sg13g2_a22oi_1 _08335_ (.Y(_03218_),
    .B1(net2241),
    .B2(net1530),
    .A2(net2287),
    .A1(net2962));
 sg13g2_a21oi_1 _08336_ (.A1(_03217_),
    .A2(_03218_),
    .Y(_03219_),
    .B1(net2074));
 sg13g2_a22oi_1 _08337_ (.Y(_03220_),
    .B1(net2139),
    .B2(net1640),
    .A2(net2183),
    .A1(net1503));
 sg13g2_a22oi_1 _08338_ (.Y(_03221_),
    .B1(net2227),
    .B2(net1431),
    .A2(net2274),
    .A1(net1451));
 sg13g2_a21oi_1 _08339_ (.A1(_03220_),
    .A2(_03221_),
    .Y(_03222_),
    .B1(net2067));
 sg13g2_nor4_1 _08340_ (.A(_03201_),
    .B(_03213_),
    .C(_03216_),
    .D(_03219_),
    .Y(_03223_));
 sg13g2_nor4_1 _08341_ (.A(_03204_),
    .B(_03207_),
    .C(_03210_),
    .D(_03222_),
    .Y(_03224_));
 sg13g2_a21oi_1 _08342_ (.A1(_03223_),
    .A2(_03224_),
    .Y(_00448_),
    .B1(net2387));
 sg13g2_a22oi_1 _08343_ (.Y(_03225_),
    .B1(net2162),
    .B2(\rf_ram.RAM[6][16] ),
    .A2(net2206),
    .A1(\rf_ram.RAM[5][16] ));
 sg13g2_a22oi_1 _08344_ (.Y(_03226_),
    .B1(net2248),
    .B2(\rf_ram.RAM[4][16] ),
    .A2(net2294),
    .A1(\rf_ram.RAM[7][16] ));
 sg13g2_a21oi_1 _08345_ (.A1(_03225_),
    .A2(_03226_),
    .Y(_03227_),
    .B1(net2262));
 sg13g2_a22oi_1 _08346_ (.Y(_03228_),
    .B1(net2154),
    .B2(net1706),
    .A2(net2198),
    .A1(net3166));
 sg13g2_a22oi_1 _08347_ (.Y(_03229_),
    .B1(net2241),
    .B2(net3129),
    .A2(net2287),
    .A1(net2783));
 sg13g2_a21oi_1 _08348_ (.A1(_03228_),
    .A2(_03229_),
    .Y(_03230_),
    .B1(net2079));
 sg13g2_a22oi_1 _08349_ (.Y(_03231_),
    .B1(net2163),
    .B2(net1688),
    .A2(net2207),
    .A1(\rf_ram.RAM[21][16] ));
 sg13g2_a22oi_1 _08350_ (.Y(_03232_),
    .B1(net2249),
    .B2(\rf_ram.RAM[20][16] ),
    .A2(net2295),
    .A1(\rf_ram.RAM[23][16] ));
 sg13g2_a21oi_1 _08351_ (.A1(_03231_),
    .A2(_03232_),
    .Y(_03233_),
    .B1(net2069));
 sg13g2_a22oi_1 _08352_ (.Y(_03234_),
    .B1(net2162),
    .B2(net1493),
    .A2(net2206),
    .A1(net3218));
 sg13g2_a22oi_1 _08353_ (.Y(_03235_),
    .B1(net2248),
    .B2(net2632),
    .A2(net2294),
    .A1(\rf_ram.RAM[19][16] ));
 sg13g2_a21oi_1 _08354_ (.A1(_03234_),
    .A2(_03235_),
    .Y(_03236_),
    .B1(net2075));
 sg13g2_a22oi_1 _08355_ (.Y(_03237_),
    .B1(net2163),
    .B2(net3190),
    .A2(net2207),
    .A1(net2745));
 sg13g2_a22oi_1 _08356_ (.Y(_03238_),
    .B1(net2249),
    .B2(net2653),
    .A2(net2305),
    .A1(net1565));
 sg13g2_a21oi_1 _08357_ (.A1(_03237_),
    .A2(_03238_),
    .Y(_03239_),
    .B1(net2310));
 sg13g2_a22oi_1 _08358_ (.Y(_03240_),
    .B1(net2154),
    .B2(net2814),
    .A2(net2198),
    .A1(net2652));
 sg13g2_a22oi_1 _08359_ (.Y(_03241_),
    .B1(net2241),
    .B2(net1665),
    .A2(net2287),
    .A1(net2661));
 sg13g2_a21oi_1 _08360_ (.A1(_03240_),
    .A2(_03241_),
    .Y(_03242_),
    .B1(net2105));
 sg13g2_a22oi_1 _08361_ (.Y(_03243_),
    .B1(net2166),
    .B2(net3140),
    .A2(net2210),
    .A1(net3134));
 sg13g2_a22oi_1 _08362_ (.Y(_03244_),
    .B1(net2252),
    .B2(net2828),
    .A2(net2295),
    .A1(net3782));
 sg13g2_a21oi_1 _08363_ (.A1(_03243_),
    .A2(_03244_),
    .Y(_03245_),
    .B1(net2101));
 sg13g2_a22oi_1 _08364_ (.Y(_03246_),
    .B1(net2154),
    .B2(net3050),
    .A2(net2198),
    .A1(net2997));
 sg13g2_a22oi_1 _08365_ (.Y(_03247_),
    .B1(net2241),
    .B2(net2758),
    .A2(net2287),
    .A1(net3079));
 sg13g2_a21oi_1 _08366_ (.A1(_03246_),
    .A2(_03247_),
    .Y(_03248_),
    .B1(net2084));
 sg13g2_nor4_1 _08367_ (.A(_03227_),
    .B(_03233_),
    .C(_03239_),
    .D(_03245_),
    .Y(_03249_));
 sg13g2_nor4_1 _08368_ (.A(_03230_),
    .B(_03236_),
    .C(_03242_),
    .D(_03248_),
    .Y(_03250_));
 sg13g2_a21oi_1 _08369_ (.A1(net3783),
    .A2(_03250_),
    .Y(_00449_),
    .B1(net2387));
 sg13g2_a22oi_1 _08370_ (.Y(_03251_),
    .B1(net2137),
    .B2(net2726),
    .A2(net2181),
    .A1(net2980));
 sg13g2_a22oi_1 _08371_ (.Y(_03252_),
    .B1(net2228),
    .B2(net3003),
    .A2(net2275),
    .A1(net1720));
 sg13g2_a21oi_1 _08372_ (.A1(_03251_),
    .A2(_03252_),
    .Y(_03253_),
    .B1(net2082));
 sg13g2_a22oi_1 _08373_ (.Y(_03254_),
    .B1(net2137),
    .B2(net1491),
    .A2(net2181),
    .A1(net3242));
 sg13g2_a22oi_1 _08374_ (.Y(_03255_),
    .B1(net2228),
    .B2(net1444),
    .A2(net2275),
    .A1(net3298));
 sg13g2_a21oi_1 _08375_ (.A1(_03254_),
    .A2(_03255_),
    .Y(_03256_),
    .B1(net2309));
 sg13g2_a22oi_1 _08376_ (.Y(_03257_),
    .B1(net2137),
    .B2(net1497),
    .A2(net2181),
    .A1(net3236));
 sg13g2_a22oi_1 _08377_ (.Y(_03258_),
    .B1(net2225),
    .B2(net2970),
    .A2(net2272),
    .A1(net2989));
 sg13g2_a21oi_1 _08378_ (.A1(_03257_),
    .A2(_03258_),
    .Y(_03259_),
    .B1(net2100));
 sg13g2_a22oi_1 _08379_ (.Y(_03260_),
    .B1(net2137),
    .B2(net2694),
    .A2(net2181),
    .A1(net2723));
 sg13g2_a22oi_1 _08380_ (.Y(_03261_),
    .B1(net2225),
    .B2(net2895),
    .A2(net2272),
    .A1(net3776));
 sg13g2_a21oi_1 _08381_ (.A1(_03260_),
    .A2(_03261_),
    .Y(_03262_),
    .B1(net2260));
 sg13g2_a22oi_1 _08382_ (.Y(_03263_),
    .B1(net2138),
    .B2(net2643),
    .A2(net2182),
    .A1(net3038));
 sg13g2_a22oi_1 _08383_ (.Y(_03264_),
    .B1(net2228),
    .B2(net2756),
    .A2(net2275),
    .A1(net3336));
 sg13g2_a21oi_1 _08384_ (.A1(_03263_),
    .A2(_03264_),
    .Y(_03265_),
    .B1(net2070));
 sg13g2_a22oi_1 _08385_ (.Y(_03266_),
    .B1(net2153),
    .B2(net1510),
    .A2(net2197),
    .A1(net2817));
 sg13g2_a22oi_1 _08386_ (.Y(_03267_),
    .B1(net2240),
    .B2(net2676),
    .A2(net2286),
    .A1(net3216));
 sg13g2_a21oi_1 _08387_ (.A1(_03266_),
    .A2(_03267_),
    .Y(_03268_),
    .B1(net2077));
 sg13g2_a22oi_1 _08388_ (.Y(_03269_),
    .B1(net2137),
    .B2(net3179),
    .A2(net2181),
    .A1(net1452));
 sg13g2_a22oi_1 _08389_ (.Y(_03270_),
    .B1(net2225),
    .B2(net1729),
    .A2(net2272),
    .A1(net1460));
 sg13g2_a21oi_1 _08390_ (.A1(_03269_),
    .A2(_03270_),
    .Y(_03271_),
    .B1(net2102));
 sg13g2_a22oi_1 _08391_ (.Y(_03272_),
    .B1(net2153),
    .B2(net3107),
    .A2(net2197),
    .A1(net2771));
 sg13g2_a22oi_1 _08392_ (.Y(_03273_),
    .B1(net2240),
    .B2(net3002),
    .A2(net2286),
    .A1(net2909));
 sg13g2_a21oi_1 _08393_ (.A1(_03272_),
    .A2(_03273_),
    .Y(_03274_),
    .B1(net2072));
 sg13g2_nor4_1 _08394_ (.A(_03253_),
    .B(_03256_),
    .C(_03265_),
    .D(_03271_),
    .Y(_03275_));
 sg13g2_nor4_1 _08395_ (.A(_03259_),
    .B(_03262_),
    .C(_03268_),
    .D(_03274_),
    .Y(_03276_));
 sg13g2_a21oi_1 _08396_ (.A1(_03275_),
    .A2(_03276_),
    .Y(_00450_),
    .B1(net2387));
 sg13g2_a22oi_1 _08397_ (.Y(_03277_),
    .B1(net2153),
    .B2(net2897),
    .A2(net2197),
    .A1(net3178));
 sg13g2_a22oi_1 _08398_ (.Y(_03278_),
    .B1(net2240),
    .B2(net2780),
    .A2(net2286),
    .A1(\rf_ram.RAM[3][18] ));
 sg13g2_a21oi_1 _08399_ (.A1(_03277_),
    .A2(_03278_),
    .Y(_03279_),
    .B1(net2309));
 sg13g2_a22oi_1 _08400_ (.Y(_03280_),
    .B1(net2153),
    .B2(net2884),
    .A2(net2197),
    .A1(\rf_ram.RAM[17][18] ));
 sg13g2_a22oi_1 _08401_ (.Y(_03281_),
    .B1(net2240),
    .B2(net1514),
    .A2(net2286),
    .A1(net3248));
 sg13g2_a21oi_1 _08402_ (.A1(_03280_),
    .A2(_03281_),
    .Y(_03282_),
    .B1(net2074));
 sg13g2_a22oi_1 _08403_ (.Y(_03283_),
    .B1(net2153),
    .B2(net1745),
    .A2(net2199),
    .A1(net1549));
 sg13g2_a22oi_1 _08404_ (.Y(_03284_),
    .B1(net2242),
    .B2(net2983),
    .A2(net2288),
    .A1(\rf_ram.RAM[15][18] ));
 sg13g2_a21oi_1 _08405_ (.A1(_03283_),
    .A2(_03284_),
    .Y(_03285_),
    .B1(net2105));
 sg13g2_a22oi_1 _08406_ (.Y(_03286_),
    .B1(net2153),
    .B2(net1435),
    .A2(net2197),
    .A1(net2615));
 sg13g2_a22oi_1 _08407_ (.Y(_03287_),
    .B1(net2240),
    .B2(net1437),
    .A2(net2286),
    .A1(net3790));
 sg13g2_a21oi_1 _08408_ (.A1(_03286_),
    .A2(_03287_),
    .Y(_03288_),
    .B1(net2070));
 sg13g2_a22oi_1 _08409_ (.Y(_03289_),
    .B1(net2152),
    .B2(net1500),
    .A2(net2196),
    .A1(net2796));
 sg13g2_a22oi_1 _08410_ (.Y(_03290_),
    .B1(net2239),
    .B2(net1527),
    .A2(net2285),
    .A1(net1748));
 sg13g2_a21oi_1 _08411_ (.A1(_03289_),
    .A2(_03290_),
    .Y(_03291_),
    .B1(net2084));
 sg13g2_a22oi_1 _08412_ (.Y(_03292_),
    .B1(net2153),
    .B2(net2832),
    .A2(net2197),
    .A1(net1610));
 sg13g2_a22oi_1 _08413_ (.Y(_03293_),
    .B1(net2240),
    .B2(net1715),
    .A2(net2286),
    .A1(net1691));
 sg13g2_a21oi_1 _08414_ (.A1(_03292_),
    .A2(_03293_),
    .Y(_03294_),
    .B1(net2079));
 sg13g2_a22oi_1 _08415_ (.Y(_03295_),
    .B1(net2155),
    .B2(net1512),
    .A2(net2199),
    .A1(net1708));
 sg13g2_a22oi_1 _08416_ (.Y(_03296_),
    .B1(net2240),
    .B2(net1648),
    .A2(net2286),
    .A1(\rf_ram.RAM[7][18] ));
 sg13g2_a21oi_1 _08417_ (.A1(_03295_),
    .A2(_03296_),
    .Y(_03297_),
    .B1(net2263));
 sg13g2_a22oi_1 _08418_ (.Y(_03298_),
    .B1(net2153),
    .B2(net2856),
    .A2(net2197),
    .A1(net1489));
 sg13g2_a22oi_1 _08419_ (.Y(_03299_),
    .B1(net2240),
    .B2(net2835),
    .A2(net2286),
    .A1(net2760));
 sg13g2_a21oi_1 _08420_ (.A1(_03298_),
    .A2(_03299_),
    .Y(_03300_),
    .B1(net2100));
 sg13g2_nor4_1 _08421_ (.A(_03279_),
    .B(_03285_),
    .C(_03291_),
    .D(_03294_),
    .Y(_03301_));
 sg13g2_nor4_1 _08422_ (.A(_03282_),
    .B(_03288_),
    .C(_03297_),
    .D(_03300_),
    .Y(_03302_));
 sg13g2_a21oi_1 _08423_ (.A1(_03301_),
    .A2(net3791),
    .Y(_00451_),
    .B1(net2387));
 sg13g2_a22oi_1 _08424_ (.Y(_03303_),
    .B1(net2136),
    .B2(\rf_ram.RAM[6][19] ),
    .A2(net2180),
    .A1(\rf_ram.RAM[5][19] ));
 sg13g2_a22oi_1 _08425_ (.Y(_03304_),
    .B1(net2225),
    .B2(\rf_ram.RAM[4][19] ),
    .A2(net2271),
    .A1(\rf_ram.RAM[7][19] ));
 sg13g2_a21oi_1 _08426_ (.A1(_03303_),
    .A2(_03304_),
    .Y(_03305_),
    .B1(net2260));
 sg13g2_a22oi_1 _08427_ (.Y(_03306_),
    .B1(net2140),
    .B2(net1508),
    .A2(net2184),
    .A1(net2801));
 sg13g2_a22oi_1 _08428_ (.Y(_03307_),
    .B1(net2226),
    .B2(net1526),
    .A2(net2273),
    .A1(\rf_ram.RAM[23][19] ));
 sg13g2_a21oi_1 _08429_ (.A1(_03306_),
    .A2(_03307_),
    .Y(_03308_),
    .B1(net2067));
 sg13g2_a22oi_1 _08430_ (.Y(_03309_),
    .B1(net2136),
    .B2(\rf_ram.RAM[10][19] ),
    .A2(net2180),
    .A1(\rf_ram.RAM[9][19] ));
 sg13g2_a22oi_1 _08431_ (.Y(_03310_),
    .B1(net2224),
    .B2(\rf_ram.RAM[8][19] ),
    .A2(net2271),
    .A1(\rf_ram.RAM[11][19] ));
 sg13g2_a21oi_1 _08432_ (.A1(_03309_),
    .A2(_03310_),
    .Y(_03311_),
    .B1(net2097));
 sg13g2_a22oi_1 _08433_ (.Y(_03312_),
    .B1(net2140),
    .B2(net1434),
    .A2(net2184),
    .A1(\rf_ram.RAM[1][19] ));
 sg13g2_a22oi_1 _08434_ (.Y(_03313_),
    .B1(net2226),
    .B2(net1566),
    .A2(net2273),
    .A1(\rf_ram.RAM[3][19] ));
 sg13g2_a21oi_1 _08435_ (.A1(_03312_),
    .A2(_03313_),
    .Y(_03314_),
    .B1(net2308));
 sg13g2_a22oi_1 _08436_ (.Y(_03315_),
    .B1(net2138),
    .B2(net1471),
    .A2(net2182),
    .A1(\rf_ram.RAM[13][19] ));
 sg13g2_a22oi_1 _08437_ (.Y(_03316_),
    .B1(net2225),
    .B2(\rf_ram.RAM[12][19] ),
    .A2(net2272),
    .A1(\rf_ram.RAM[15][19] ));
 sg13g2_a21oi_1 _08438_ (.A1(_03315_),
    .A2(_03316_),
    .Y(_03317_),
    .B1(net2102));
 sg13g2_a22oi_1 _08439_ (.Y(_03318_),
    .B1(net2133),
    .B2(net3807),
    .A2(net2177),
    .A1(\rf_ram.RAM[29][19] ));
 sg13g2_a22oi_1 _08440_ (.Y(_03319_),
    .B1(net2222),
    .B2(\rf_ram.RAM[28][19] ),
    .A2(net2269),
    .A1(\rf_ram.RAM[31][19] ));
 sg13g2_a21oi_1 _08441_ (.A1(_03318_),
    .A2(_03319_),
    .Y(_03320_),
    .B1(net2077));
 sg13g2_a22oi_1 _08442_ (.Y(_03321_),
    .B1(net2136),
    .B2(\rf_ram.RAM[18][19] ),
    .A2(net2180),
    .A1(\rf_ram.RAM[17][19] ));
 sg13g2_a22oi_1 _08443_ (.Y(_03322_),
    .B1(net2224),
    .B2(\rf_ram.RAM[16][19] ),
    .A2(net2271),
    .A1(\rf_ram.RAM[19][19] ));
 sg13g2_a21oi_1 _08444_ (.A1(_03321_),
    .A2(_03322_),
    .Y(_03323_),
    .B1(net2072));
 sg13g2_a22oi_1 _08445_ (.Y(_03324_),
    .B1(net2140),
    .B2(\rf_ram.RAM[26][19] ),
    .A2(net2184),
    .A1(\rf_ram.RAM[25][19] ));
 sg13g2_a22oi_1 _08446_ (.Y(_03325_),
    .B1(net2226),
    .B2(\rf_ram.RAM[24][19] ),
    .A2(net2273),
    .A1(\rf_ram.RAM[27][19] ));
 sg13g2_a21oi_1 _08447_ (.A1(_03324_),
    .A2(_03325_),
    .Y(_03326_),
    .B1(net2082));
 sg13g2_nor4_1 _08448_ (.A(_03305_),
    .B(_03311_),
    .C(_03317_),
    .D(_03320_),
    .Y(_03327_));
 sg13g2_nor4_1 _08449_ (.A(_03308_),
    .B(_03314_),
    .C(_03323_),
    .D(_03326_),
    .Y(_03328_));
 sg13g2_a21oi_1 _08450_ (.A1(net3808),
    .A2(_03328_),
    .Y(_00452_),
    .B1(net2385));
 sg13g2_a22oi_1 _08451_ (.Y(_03329_),
    .B1(net2140),
    .B2(net1554),
    .A2(net2184),
    .A1(net1567));
 sg13g2_a22oi_1 _08452_ (.Y(_03330_),
    .B1(net2226),
    .B2(net3074),
    .A2(net2273),
    .A1(net3154));
 sg13g2_a21oi_1 _08453_ (.A1(_03329_),
    .A2(_03330_),
    .Y(_03331_),
    .B1(net2102));
 sg13g2_a22oi_1 _08454_ (.Y(_03332_),
    .B1(net2139),
    .B2(net2670),
    .A2(net2183),
    .A1(net2636));
 sg13g2_a22oi_1 _08455_ (.Y(_03333_),
    .B1(net2227),
    .B2(net2935),
    .A2(net2274),
    .A1(net3013));
 sg13g2_a21oi_1 _08456_ (.A1(_03332_),
    .A2(_03333_),
    .Y(_03334_),
    .B1(net2077));
 sg13g2_a22oi_1 _08457_ (.Y(_03335_),
    .B1(net2139),
    .B2(net2976),
    .A2(net2183),
    .A1(net1592));
 sg13g2_a22oi_1 _08458_ (.Y(_03336_),
    .B1(net2226),
    .B2(net1602),
    .A2(net2273),
    .A1(net2905));
 sg13g2_a21oi_1 _08459_ (.A1(_03335_),
    .A2(_03336_),
    .Y(_03337_),
    .B1(net2097));
 sg13g2_a22oi_1 _08460_ (.Y(_03338_),
    .B1(net2139),
    .B2(net3001),
    .A2(net2183),
    .A1(net1616));
 sg13g2_a22oi_1 _08461_ (.Y(_03339_),
    .B1(net2227),
    .B2(net2692),
    .A2(net2274),
    .A1(net2609));
 sg13g2_a21oi_1 _08462_ (.A1(_03338_),
    .A2(_03339_),
    .Y(_03340_),
    .B1(net2260));
 sg13g2_a22oi_1 _08463_ (.Y(_03341_),
    .B1(net2140),
    .B2(net2606),
    .A2(net2184),
    .A1(net1732));
 sg13g2_a22oi_1 _08464_ (.Y(_03342_),
    .B1(net2226),
    .B2(net2786),
    .A2(net2273),
    .A1(net1683));
 sg13g2_a21oi_1 _08465_ (.A1(_03341_),
    .A2(_03342_),
    .Y(_03343_),
    .B1(net2308));
 sg13g2_a22oi_1 _08466_ (.Y(_03344_),
    .B1(net2141),
    .B2(net1663),
    .A2(net2185),
    .A1(net3300));
 sg13g2_a22oi_1 _08467_ (.Y(_03345_),
    .B1(net2227),
    .B2(net3283),
    .A2(net2274),
    .A1(net3239));
 sg13g2_a21oi_1 _08468_ (.A1(_03344_),
    .A2(_03345_),
    .Y(_03346_),
    .B1(net2082));
 sg13g2_a22oi_1 _08469_ (.Y(_03347_),
    .B1(net2140),
    .B2(net3082),
    .A2(net2184),
    .A1(net3244));
 sg13g2_a22oi_1 _08470_ (.Y(_03348_),
    .B1(net2226),
    .B2(net2979),
    .A2(net2273),
    .A1(net3306));
 sg13g2_a21oi_1 _08471_ (.A1(_03347_),
    .A2(_03348_),
    .Y(_03349_),
    .B1(net2067));
 sg13g2_a22oi_1 _08472_ (.Y(_03350_),
    .B1(net2139),
    .B2(net3118),
    .A2(net2183),
    .A1(net3231));
 sg13g2_a22oi_1 _08473_ (.Y(_03351_),
    .B1(net2227),
    .B2(net2813),
    .A2(net2274),
    .A1(net1659));
 sg13g2_a21oi_1 _08474_ (.A1(_03350_),
    .A2(_03351_),
    .Y(_03352_),
    .B1(net2072));
 sg13g2_nor4_1 _08475_ (.A(_03331_),
    .B(_03337_),
    .C(_03343_),
    .D(_03349_),
    .Y(_03353_));
 sg13g2_nor4_1 _08476_ (.A(_03334_),
    .B(_03340_),
    .C(_03346_),
    .D(_03352_),
    .Y(_03354_));
 sg13g2_a21oi_1 _08477_ (.A1(_03353_),
    .A2(_03354_),
    .Y(_00453_),
    .B1(net2385));
 sg13g2_a22oi_1 _08478_ (.Y(_03355_),
    .B1(net2150),
    .B2(net1535),
    .A2(net2194),
    .A1(net3167));
 sg13g2_a22oi_1 _08479_ (.Y(_03356_),
    .B1(net2237),
    .B2(net3194),
    .A2(net2283),
    .A1(net2802));
 sg13g2_a21oi_1 _08480_ (.A1(_03355_),
    .A2(_03356_),
    .Y(_03357_),
    .B1(net2098));
 sg13g2_a22oi_1 _08481_ (.Y(_03358_),
    .B1(net2147),
    .B2(net1689),
    .A2(net2191),
    .A1(net1711));
 sg13g2_a22oi_1 _08482_ (.Y(_03359_),
    .B1(net2233),
    .B2(net1443),
    .A2(net2280),
    .A1(net1614));
 sg13g2_a21oi_1 _08483_ (.A1(_03358_),
    .A2(_03359_),
    .Y(_03360_),
    .B1(net2312));
 sg13g2_a22oi_1 _08484_ (.Y(_03361_),
    .B1(net2147),
    .B2(net3068),
    .A2(net2191),
    .A1(net3177));
 sg13g2_a22oi_1 _08485_ (.Y(_03362_),
    .B1(net2233),
    .B2(net1541),
    .A2(net2280),
    .A1(net3025));
 sg13g2_a21oi_1 _08486_ (.A1(_03361_),
    .A2(_03362_),
    .Y(_03363_),
    .B1(net2068));
 sg13g2_a22oi_1 _08487_ (.Y(_03364_),
    .B1(net2147),
    .B2(net2774),
    .A2(net2191),
    .A1(net2951));
 sg13g2_a22oi_1 _08488_ (.Y(_03365_),
    .B1(net2233),
    .B2(net2847),
    .A2(net2280),
    .A1(net2623));
 sg13g2_a21oi_1 _08489_ (.A1(_03364_),
    .A2(_03365_),
    .Y(_03366_),
    .B1(net2261));
 sg13g2_a22oi_1 _08490_ (.Y(_03367_),
    .B1(net2150),
    .B2(net2633),
    .A2(net2194),
    .A1(net3030));
 sg13g2_a22oi_1 _08491_ (.Y(_03368_),
    .B1(net2237),
    .B2(net3259),
    .A2(net2283),
    .A1(net3278));
 sg13g2_a21oi_1 _08492_ (.A1(_03367_),
    .A2(_03368_),
    .Y(_03369_),
    .B1(net2103));
 sg13g2_a22oi_1 _08493_ (.Y(_03370_),
    .B1(net2150),
    .B2(net1568),
    .A2(net2194),
    .A1(net3296));
 sg13g2_a22oi_1 _08494_ (.Y(_03371_),
    .B1(net2235),
    .B2(net1742),
    .A2(net2283),
    .A1(net1625));
 sg13g2_a21oi_1 _08495_ (.A1(_03370_),
    .A2(_03371_),
    .Y(_03372_),
    .B1(net2083));
 sg13g2_a22oi_1 _08496_ (.Y(_03373_),
    .B1(net2147),
    .B2(net3017),
    .A2(net2191),
    .A1(net2871));
 sg13g2_a22oi_1 _08497_ (.Y(_03374_),
    .B1(net2233),
    .B2(net3324),
    .A2(net2283),
    .A1(net3252));
 sg13g2_a21oi_1 _08498_ (.A1(_03373_),
    .A2(_03374_),
    .Y(_03375_),
    .B1(net2078));
 sg13g2_a22oi_1 _08499_ (.Y(_03376_),
    .B1(net2150),
    .B2(net1583),
    .A2(net2194),
    .A1(net2797));
 sg13g2_a22oi_1 _08500_ (.Y(_03377_),
    .B1(net2237),
    .B2(net2769),
    .A2(net2280),
    .A1(net2870));
 sg13g2_a21oi_1 _08501_ (.A1(_03376_),
    .A2(_03377_),
    .Y(_03378_),
    .B1(net2073));
 sg13g2_nor4_1 _08502_ (.A(_03363_),
    .B(_03369_),
    .C(_03372_),
    .D(_03375_),
    .Y(_03379_));
 sg13g2_nor4_1 _08503_ (.A(_03357_),
    .B(_03360_),
    .C(_03366_),
    .D(_03378_),
    .Y(_03380_));
 sg13g2_a21oi_1 _08504_ (.A1(_03379_),
    .A2(_03380_),
    .Y(_00454_),
    .B1(net2385));
 sg13g2_a22oi_1 _08505_ (.Y(_03381_),
    .B1(net2162),
    .B2(net1604),
    .A2(net2206),
    .A1(net2821));
 sg13g2_a22oi_1 _08506_ (.Y(_03382_),
    .B1(net2248),
    .B2(net3238),
    .A2(net2294),
    .A1(net1629));
 sg13g2_a21oi_1 _08507_ (.A1(_03381_),
    .A2(_03382_),
    .Y(_03383_),
    .B1(net2262));
 sg13g2_a22oi_1 _08508_ (.Y(_03384_),
    .B1(net2163),
    .B2(net1643),
    .A2(net2207),
    .A1(net2648));
 sg13g2_a22oi_1 _08509_ (.Y(_03385_),
    .B1(net2248),
    .B2(net3295),
    .A2(net2294),
    .A1(net3302));
 sg13g2_a21oi_1 _08510_ (.A1(_03384_),
    .A2(_03385_),
    .Y(_03386_),
    .B1(net2086));
 sg13g2_a22oi_1 _08511_ (.Y(_03387_),
    .B1(net2162),
    .B2(net3297),
    .A2(net2206),
    .A1(net3260));
 sg13g2_a22oi_1 _08512_ (.Y(_03388_),
    .B1(net2248),
    .B2(net2972),
    .A2(net2294),
    .A1(net3789));
 sg13g2_a21oi_1 _08513_ (.A1(_03387_),
    .A2(_03388_),
    .Y(_03389_),
    .B1(net2075));
 sg13g2_a22oi_1 _08514_ (.Y(_03390_),
    .B1(net2163),
    .B2(net2641),
    .A2(net2207),
    .A1(net2805));
 sg13g2_a22oi_1 _08515_ (.Y(_03391_),
    .B1(net2249),
    .B2(net3027),
    .A2(net2295),
    .A1(net1727));
 sg13g2_a21oi_1 _08516_ (.A1(_03390_),
    .A2(_03391_),
    .Y(_03392_),
    .B1(net2069));
 sg13g2_a22oi_1 _08517_ (.Y(_03393_),
    .B1(net2162),
    .B2(net2674),
    .A2(net2206),
    .A1(net2886));
 sg13g2_a22oi_1 _08518_ (.Y(_03394_),
    .B1(net2248),
    .B2(net3219),
    .A2(net2294),
    .A1(net2604));
 sg13g2_a21oi_1 _08519_ (.A1(_03393_),
    .A2(_03394_),
    .Y(_03395_),
    .B1(net2099));
 sg13g2_a22oi_1 _08520_ (.Y(_03396_),
    .B1(net2162),
    .B2(net2915),
    .A2(net2206),
    .A1(net3322));
 sg13g2_a22oi_1 _08521_ (.Y(_03397_),
    .B1(net2248),
    .B2(net2931),
    .A2(net2295),
    .A1(net3123));
 sg13g2_a21oi_1 _08522_ (.A1(_03396_),
    .A2(_03397_),
    .Y(_03398_),
    .B1(net2310));
 sg13g2_a22oi_1 _08523_ (.Y(_03399_),
    .B1(net2162),
    .B2(net3210),
    .A2(net2206),
    .A1(net2792));
 sg13g2_a22oi_1 _08524_ (.Y(_03400_),
    .B1(net2248),
    .B2(net1664),
    .A2(net2294),
    .A1(net1543));
 sg13g2_a21oi_1 _08525_ (.A1(_03399_),
    .A2(_03400_),
    .Y(_03401_),
    .B1(net2080));
 sg13g2_a22oi_1 _08526_ (.Y(_03402_),
    .B1(net2162),
    .B2(net1476),
    .A2(net2206),
    .A1(net2892));
 sg13g2_a22oi_1 _08527_ (.Y(_03403_),
    .B1(net2249),
    .B2(net3024),
    .A2(net2294),
    .A1(net1710));
 sg13g2_a21oi_1 _08528_ (.A1(_03402_),
    .A2(_03403_),
    .Y(_03404_),
    .B1(net2104));
 sg13g2_nor4_1 _08529_ (.A(_03383_),
    .B(_03389_),
    .C(_03401_),
    .D(_03404_),
    .Y(_03405_));
 sg13g2_nor4_1 _08530_ (.A(_03386_),
    .B(_03392_),
    .C(_03395_),
    .D(_03398_),
    .Y(_03406_));
 sg13g2_a21oi_1 _08531_ (.A1(_03405_),
    .A2(_03406_),
    .Y(_00455_),
    .B1(net2387));
 sg13g2_a22oi_1 _08532_ (.Y(_03407_),
    .B1(net2147),
    .B2(net3247),
    .A2(net2191),
    .A1(net3241));
 sg13g2_a22oi_1 _08533_ (.Y(_03408_),
    .B1(net2233),
    .B2(net1694),
    .A2(net2280),
    .A1(net2725));
 sg13g2_a21oi_1 _08534_ (.A1(_03407_),
    .A2(_03408_),
    .Y(_03409_),
    .B1(net2103));
 sg13g2_a22oi_1 _08535_ (.Y(_03410_),
    .B1(net2133),
    .B2(net3229),
    .A2(net2177),
    .A1(net3052));
 sg13g2_a22oi_1 _08536_ (.Y(_03411_),
    .B1(net2221),
    .B2(net1606),
    .A2(net2268),
    .A1(net3037));
 sg13g2_a21oi_1 _08537_ (.A1(_03410_),
    .A2(_03411_),
    .Y(_03412_),
    .B1(net2308));
 sg13g2_a22oi_1 _08538_ (.Y(_03413_),
    .B1(net2147),
    .B2(net1487),
    .A2(net2191),
    .A1(net1608));
 sg13g2_a22oi_1 _08539_ (.Y(_03414_),
    .B1(net2233),
    .B2(net1499),
    .A2(net2280),
    .A1(net2864));
 sg13g2_a21oi_1 _08540_ (.A1(_03413_),
    .A2(_03414_),
    .Y(_03415_),
    .B1(net2078));
 sg13g2_a22oi_1 _08541_ (.Y(_03416_),
    .B1(net2140),
    .B2(net3035),
    .A2(net2184),
    .A1(net1743));
 sg13g2_a22oi_1 _08542_ (.Y(_03417_),
    .B1(net2222),
    .B2(net3224),
    .A2(net2269),
    .A1(net2883));
 sg13g2_a21oi_1 _08543_ (.A1(_03416_),
    .A2(_03417_),
    .Y(_03418_),
    .B1(net2097));
 sg13g2_a22oi_1 _08544_ (.Y(_03419_),
    .B1(net2143),
    .B2(net2912),
    .A2(net2187),
    .A1(net3781));
 sg13g2_a22oi_1 _08545_ (.Y(_03420_),
    .B1(net2229),
    .B2(net1458),
    .A2(net2279),
    .A1(\rf_ram.RAM[27][23] ));
 sg13g2_a21oi_1 _08546_ (.A1(_03419_),
    .A2(_03420_),
    .Y(_03421_),
    .B1(net2083));
 sg13g2_a22oi_1 _08547_ (.Y(_03422_),
    .B1(net2143),
    .B2(net1741),
    .A2(net2187),
    .A1(net2863));
 sg13g2_a22oi_1 _08548_ (.Y(_03423_),
    .B1(net2229),
    .B2(net3124),
    .A2(net2279),
    .A1(net1577));
 sg13g2_a21oi_1 _08549_ (.A1(_03422_),
    .A2(_03423_),
    .Y(_03424_),
    .B1(net2068));
 sg13g2_a22oi_1 _08550_ (.Y(_03425_),
    .B1(net2140),
    .B2(net2736),
    .A2(net2184),
    .A1(net3006));
 sg13g2_a22oi_1 _08551_ (.Y(_03426_),
    .B1(net2226),
    .B2(net3113),
    .A2(net2273),
    .A1(net1669));
 sg13g2_a21oi_1 _08552_ (.A1(_03425_),
    .A2(_03426_),
    .Y(_03427_),
    .B1(net2260));
 sg13g2_a22oi_1 _08553_ (.Y(_03428_),
    .B1(net2147),
    .B2(net3105),
    .A2(net2191),
    .A1(net2630));
 sg13g2_a22oi_1 _08554_ (.Y(_03429_),
    .B1(net2233),
    .B2(net2921),
    .A2(net2280),
    .A1(net1558));
 sg13g2_a21oi_1 _08555_ (.A1(_03428_),
    .A2(_03429_),
    .Y(_03430_),
    .B1(net2073));
 sg13g2_nor4_1 _08556_ (.A(_03409_),
    .B(_03415_),
    .C(_03421_),
    .D(_03424_),
    .Y(_03431_));
 sg13g2_nor4_1 _08557_ (.A(_03412_),
    .B(_03418_),
    .C(_03427_),
    .D(_03430_),
    .Y(_03432_));
 sg13g2_a21oi_1 _08558_ (.A1(_03431_),
    .A2(_03432_),
    .Y(_00456_),
    .B1(net2385));
 sg13g2_a22oi_1 _08559_ (.Y(_03433_),
    .B1(net2149),
    .B2(net2790),
    .A2(net2193),
    .A1(net2624));
 sg13g2_a22oi_1 _08560_ (.Y(_03434_),
    .B1(net2235),
    .B2(net3204),
    .A2(net2282),
    .A1(net1667));
 sg13g2_a21oi_1 _08561_ (.A1(_03433_),
    .A2(_03434_),
    .Y(_03435_),
    .B1(net2078));
 sg13g2_a22oi_1 _08562_ (.Y(_03436_),
    .B1(net2164),
    .B2(net3176),
    .A2(net2208),
    .A1(net3220));
 sg13g2_a22oi_1 _08563_ (.Y(_03437_),
    .B1(net2251),
    .B2(net3291),
    .A2(net2296),
    .A1(net1699));
 sg13g2_a21oi_1 _08564_ (.A1(_03436_),
    .A2(_03437_),
    .Y(_03438_),
    .B1(net2085));
 sg13g2_a22oi_1 _08565_ (.Y(_03439_),
    .B1(net2165),
    .B2(net2675),
    .A2(net2208),
    .A1(net1603));
 sg13g2_a22oi_1 _08566_ (.Y(_03440_),
    .B1(net2235),
    .B2(net2746),
    .A2(net2282),
    .A1(net3159));
 sg13g2_a21oi_1 _08567_ (.A1(_03439_),
    .A2(_03440_),
    .Y(_03441_),
    .B1(net2069));
 sg13g2_a22oi_1 _08568_ (.Y(_03442_),
    .B1(net2164),
    .B2(net3227),
    .A2(net2208),
    .A1(net2838));
 sg13g2_a22oi_1 _08569_ (.Y(_03443_),
    .B1(net2251),
    .B2(net2724),
    .A2(net2296),
    .A1(net1695));
 sg13g2_a21oi_1 _08570_ (.A1(_03442_),
    .A2(_03443_),
    .Y(_03444_),
    .B1(net2262));
 sg13g2_a22oi_1 _08571_ (.Y(_03445_),
    .B1(net2149),
    .B2(net1662),
    .A2(net2193),
    .A1(net2755));
 sg13g2_a22oi_1 _08572_ (.Y(_03446_),
    .B1(net2235),
    .B2(net2656),
    .A2(net2282),
    .A1(net2655));
 sg13g2_a21oi_1 _08573_ (.A1(_03445_),
    .A2(_03446_),
    .Y(_03447_),
    .B1(net2073));
 sg13g2_a22oi_1 _08574_ (.Y(_03448_),
    .B1(net2164),
    .B2(net1722),
    .A2(net2209),
    .A1(net3106));
 sg13g2_a22oi_1 _08575_ (.Y(_03449_),
    .B1(net2251),
    .B2(net2940),
    .A2(net2296),
    .A1(net3249));
 sg13g2_a21oi_1 _08576_ (.A1(_03448_),
    .A2(_03449_),
    .Y(_03450_),
    .B1(net2104));
 sg13g2_a22oi_1 _08577_ (.Y(_03451_),
    .B1(net2165),
    .B2(net3057),
    .A2(net2209),
    .A1(net2733));
 sg13g2_a22oi_1 _08578_ (.Y(_03452_),
    .B1(net2251),
    .B2(net1556),
    .A2(net2296),
    .A1(net2857));
 sg13g2_a21oi_1 _08579_ (.A1(_03451_),
    .A2(_03452_),
    .Y(_03453_),
    .B1(net2310));
 sg13g2_a22oi_1 _08580_ (.Y(_03454_),
    .B1(net2164),
    .B2(net2759),
    .A2(net2208),
    .A1(net1548));
 sg13g2_a22oi_1 _08581_ (.Y(_03455_),
    .B1(net2251),
    .B2(net2879),
    .A2(net2296),
    .A1(net2787));
 sg13g2_a21oi_1 _08582_ (.A1(_03454_),
    .A2(_03455_),
    .Y(_03456_),
    .B1(net2099));
 sg13g2_nor4_1 _08583_ (.A(_03435_),
    .B(_03441_),
    .C(_03447_),
    .D(_03453_),
    .Y(_03457_));
 sg13g2_nor4_1 _08584_ (.A(_03438_),
    .B(_03444_),
    .C(_03450_),
    .D(_03456_),
    .Y(_03458_));
 sg13g2_a21oi_1 _08585_ (.A1(_03457_),
    .A2(_03458_),
    .Y(_00457_),
    .B1(net2387));
 sg13g2_a22oi_1 _08586_ (.Y(_03459_),
    .B1(net2148),
    .B2(net2986),
    .A2(net2192),
    .A1(net2743));
 sg13g2_a22oi_1 _08587_ (.Y(_03460_),
    .B1(net2234),
    .B2(net1678),
    .A2(net2277),
    .A1(net1698));
 sg13g2_a21oi_1 _08588_ (.A1(_03459_),
    .A2(_03460_),
    .Y(_03461_),
    .B1(net2073));
 sg13g2_a22oi_1 _08589_ (.Y(_03462_),
    .B1(net2148),
    .B2(net1653),
    .A2(net2192),
    .A1(net2908));
 sg13g2_a22oi_1 _08590_ (.Y(_03463_),
    .B1(net2234),
    .B2(net2827),
    .A2(net2281),
    .A1(net2705));
 sg13g2_a21oi_1 _08591_ (.A1(_03462_),
    .A2(_03463_),
    .Y(_03464_),
    .B1(net2078));
 sg13g2_a22oi_1 _08592_ (.Y(_03465_),
    .B1(net2149),
    .B2(net2872),
    .A2(net2193),
    .A1(net3072));
 sg13g2_a22oi_1 _08593_ (.Y(_03466_),
    .B1(net2236),
    .B2(net2752),
    .A2(net2282),
    .A1(net3023));
 sg13g2_a21oi_1 _08594_ (.A1(_03465_),
    .A2(_03466_),
    .Y(_03467_),
    .B1(net2103));
 sg13g2_a22oi_1 _08595_ (.Y(_03468_),
    .B1(net2145),
    .B2(net1544),
    .A2(net2189),
    .A1(net2873));
 sg13g2_a22oi_1 _08596_ (.Y(_03469_),
    .B1(net2231),
    .B2(net3078),
    .A2(net2277),
    .A1(net1652));
 sg13g2_a21oi_1 _08597_ (.A1(_03468_),
    .A2(_03469_),
    .Y(_03470_),
    .B1(net2068));
 sg13g2_a22oi_1 _08598_ (.Y(_03471_),
    .B1(net2145),
    .B2(net1464),
    .A2(net2189),
    .A1(net1626));
 sg13g2_a22oi_1 _08599_ (.Y(_03472_),
    .B1(net2231),
    .B2(net2950),
    .A2(net2279),
    .A1(net1627));
 sg13g2_a21oi_1 _08600_ (.A1(_03471_),
    .A2(_03472_),
    .Y(_03473_),
    .B1(net2307));
 sg13g2_a22oi_1 _08601_ (.Y(_03474_),
    .B1(net2145),
    .B2(net1536),
    .A2(net2189),
    .A1(net3208));
 sg13g2_a22oi_1 _08602_ (.Y(_03475_),
    .B1(net2231),
    .B2(net1425),
    .A2(net2277),
    .A1(net2875));
 sg13g2_a21oi_1 _08603_ (.A1(_03474_),
    .A2(_03475_),
    .Y(_03476_),
    .B1(net2098));
 sg13g2_a22oi_1 _08604_ (.Y(_03477_),
    .B1(net2142),
    .B2(net1679),
    .A2(net2186),
    .A1(net1674));
 sg13g2_a22oi_1 _08605_ (.Y(_03478_),
    .B1(net2229),
    .B2(net1465),
    .A2(net2276),
    .A1(net3775));
 sg13g2_a21oi_1 _08606_ (.A1(_03477_),
    .A2(_03478_),
    .Y(_03479_),
    .B1(net2261));
 sg13g2_a22oi_1 _08607_ (.Y(_03480_),
    .B1(net2145),
    .B2(net2974),
    .A2(net2189),
    .A1(net3026));
 sg13g2_a22oi_1 _08608_ (.Y(_03481_),
    .B1(net2231),
    .B2(net3193),
    .A2(net2277),
    .A1(net2616));
 sg13g2_a21oi_1 _08609_ (.A1(_03480_),
    .A2(_03481_),
    .Y(_03482_),
    .B1(net2083));
 sg13g2_nor4_1 _08610_ (.A(_03461_),
    .B(_03464_),
    .C(_03467_),
    .D(_03479_),
    .Y(_03483_));
 sg13g2_nor4_1 _08611_ (.A(_03470_),
    .B(_03473_),
    .C(_03476_),
    .D(_03482_),
    .Y(_03484_));
 sg13g2_a21oi_1 _08612_ (.A1(_03483_),
    .A2(_03484_),
    .Y(_00458_),
    .B1(net2384));
 sg13g2_a22oi_1 _08613_ (.Y(_03485_),
    .B1(net2145),
    .B2(\rf_ram.RAM[22][26] ),
    .A2(net2189),
    .A1(\rf_ram.RAM[21][26] ));
 sg13g2_a22oi_1 _08614_ (.Y(_03486_),
    .B1(net2231),
    .B2(\rf_ram.RAM[20][26] ),
    .A2(net2277),
    .A1(\rf_ram.RAM[23][26] ));
 sg13g2_a21oi_1 _08615_ (.A1(_03485_),
    .A2(_03486_),
    .Y(_03487_),
    .B1(net2068));
 sg13g2_a22oi_1 _08616_ (.Y(_03488_),
    .B1(net2145),
    .B2(net3205),
    .A2(net2189),
    .A1(net3098));
 sg13g2_a22oi_1 _08617_ (.Y(_03489_),
    .B1(net2231),
    .B2(net3031),
    .A2(net2277),
    .A1(\rf_ram.RAM[3][26] ));
 sg13g2_a21oi_1 _08618_ (.A1(_03488_),
    .A2(_03489_),
    .Y(_03490_),
    .B1(net2312));
 sg13g2_a22oi_1 _08619_ (.Y(_03491_),
    .B1(net2145),
    .B2(net1517),
    .A2(net2189),
    .A1(net1584));
 sg13g2_a22oi_1 _08620_ (.Y(_03492_),
    .B1(net2231),
    .B2(net1520),
    .A2(net2277),
    .A1(net2984));
 sg13g2_a21oi_1 _08621_ (.A1(_03491_),
    .A2(_03492_),
    .Y(_03493_),
    .B1(net2073));
 sg13g2_a22oi_1 _08622_ (.Y(_03494_),
    .B1(net2147),
    .B2(\rf_ram.RAM[10][26] ),
    .A2(net2191),
    .A1(\rf_ram.RAM[9][26] ));
 sg13g2_a22oi_1 _08623_ (.Y(_03495_),
    .B1(net2233),
    .B2(\rf_ram.RAM[8][26] ),
    .A2(net2280),
    .A1(\rf_ram.RAM[11][26] ));
 sg13g2_a21oi_1 _08624_ (.A1(_03494_),
    .A2(_03495_),
    .Y(_03496_),
    .B1(net2098));
 sg13g2_a22oi_1 _08625_ (.Y(_03497_),
    .B1(net2148),
    .B2(\rf_ram.RAM[26][26] ),
    .A2(net2192),
    .A1(\rf_ram.RAM[25][26] ));
 sg13g2_a22oi_1 _08626_ (.Y(_03498_),
    .B1(net2234),
    .B2(\rf_ram.RAM[24][26] ),
    .A2(net2281),
    .A1(\rf_ram.RAM[27][26] ));
 sg13g2_a21oi_1 _08627_ (.A1(_03497_),
    .A2(_03498_),
    .Y(_03499_),
    .B1(net2083));
 sg13g2_a22oi_1 _08628_ (.Y(_03500_),
    .B1(net2148),
    .B2(\rf_ram.RAM[30][26] ),
    .A2(net2192),
    .A1(\rf_ram.RAM[29][26] ));
 sg13g2_a22oi_1 _08629_ (.Y(_03501_),
    .B1(net2234),
    .B2(\rf_ram.RAM[28][26] ),
    .A2(net2281),
    .A1(\rf_ram.RAM[31][26] ));
 sg13g2_a21oi_1 _08630_ (.A1(_03500_),
    .A2(_03501_),
    .Y(_03502_),
    .B1(net2078));
 sg13g2_a22oi_1 _08631_ (.Y(_03503_),
    .B1(net2145),
    .B2(net3086),
    .A2(net2189),
    .A1(net2964));
 sg13g2_a22oi_1 _08632_ (.Y(_03504_),
    .B1(net2231),
    .B2(net2937),
    .A2(net2277),
    .A1(net2668));
 sg13g2_a21oi_1 _08633_ (.A1(_03503_),
    .A2(_03504_),
    .Y(_03505_),
    .B1(net2106));
 sg13g2_a22oi_1 _08634_ (.Y(_03506_),
    .B1(net2148),
    .B2(net1725),
    .A2(net2192),
    .A1(net2804));
 sg13g2_a22oi_1 _08635_ (.Y(_03507_),
    .B1(net2234),
    .B2(net1623),
    .A2(net2281),
    .A1(net3794));
 sg13g2_a21oi_1 _08636_ (.A1(_03506_),
    .A2(_03507_),
    .Y(_03508_),
    .B1(net2261));
 sg13g2_nor4_1 _08637_ (.A(_03487_),
    .B(_03490_),
    .C(_03493_),
    .D(_03505_),
    .Y(_03509_));
 sg13g2_nor4_1 _08638_ (.A(_03496_),
    .B(_03499_),
    .C(_03502_),
    .D(_03508_),
    .Y(_03510_));
 sg13g2_a21oi_2 _08639_ (.B1(net2384),
    .Y(_00459_),
    .A2(_03510_),
    .A1(_03509_));
 sg13g2_a22oi_1 _08640_ (.Y(_03511_),
    .B1(net2144),
    .B2(net1496),
    .A2(net2188),
    .A1(net2735));
 sg13g2_a22oi_1 _08641_ (.Y(_03512_),
    .B1(net2230),
    .B2(net2779),
    .A2(net2278),
    .A1(net2910));
 sg13g2_a21oi_1 _08642_ (.A1(_03511_),
    .A2(_03512_),
    .Y(_03513_),
    .B1(net2307));
 sg13g2_a22oi_1 _08643_ (.Y(_03514_),
    .B1(net2144),
    .B2(net2685),
    .A2(net2188),
    .A1(net2818));
 sg13g2_a22oi_1 _08644_ (.Y(_03515_),
    .B1(net2230),
    .B2(net3120),
    .A2(net2278),
    .A1(net3313));
 sg13g2_a21oi_1 _08645_ (.A1(_03514_),
    .A2(_03515_),
    .Y(_03516_),
    .B1(net2068));
 sg13g2_a22oi_1 _08646_ (.Y(_03517_),
    .B1(net2144),
    .B2(net2731),
    .A2(net2188),
    .A1(net2721));
 sg13g2_a22oi_1 _08647_ (.Y(_03518_),
    .B1(net2230),
    .B2(net1563),
    .A2(net2278),
    .A1(net3089));
 sg13g2_a21oi_1 _08648_ (.A1(_03517_),
    .A2(_03518_),
    .Y(_03519_),
    .B1(net2103));
 sg13g2_a22oi_1 _08649_ (.Y(_03520_),
    .B1(net2144),
    .B2(net1579),
    .A2(net2188),
    .A1(net3214));
 sg13g2_a22oi_1 _08650_ (.Y(_03521_),
    .B1(net2230),
    .B2(net3228),
    .A2(net2278),
    .A1(net2688));
 sg13g2_a21oi_1 _08651_ (.A1(_03520_),
    .A2(_03521_),
    .Y(_03522_),
    .B1(net2098));
 sg13g2_a22oi_1 _08652_ (.Y(_03523_),
    .B1(net2144),
    .B2(net3016),
    .A2(net2188),
    .A1(net3189));
 sg13g2_a22oi_1 _08653_ (.Y(_03524_),
    .B1(net2230),
    .B2(net3323),
    .A2(net2278),
    .A1(net3048));
 sg13g2_a21oi_1 _08654_ (.A1(_03523_),
    .A2(_03524_),
    .Y(_03525_),
    .B1(net2083));
 sg13g2_a22oi_1 _08655_ (.Y(_03526_),
    .B1(net2144),
    .B2(net2730),
    .A2(net2188),
    .A1(net2764));
 sg13g2_a22oi_1 _08656_ (.Y(_03527_),
    .B1(net2230),
    .B2(net1738),
    .A2(net2278),
    .A1(net1574));
 sg13g2_a21oi_1 _08657_ (.A1(_03526_),
    .A2(_03527_),
    .Y(_03528_),
    .B1(net2073));
 sg13g2_a22oi_1 _08658_ (.Y(_03529_),
    .B1(net2144),
    .B2(net2767),
    .A2(net2188),
    .A1(net2967));
 sg13g2_a22oi_1 _08659_ (.Y(_03530_),
    .B1(net2230),
    .B2(net2815),
    .A2(net2278),
    .A1(net2784));
 sg13g2_a21oi_1 _08660_ (.A1(_03529_),
    .A2(_03530_),
    .Y(_03531_),
    .B1(net2078));
 sg13g2_a22oi_1 _08661_ (.Y(_03532_),
    .B1(net2144),
    .B2(net2754),
    .A2(net2188),
    .A1(net2900));
 sg13g2_a22oi_1 _08662_ (.Y(_03533_),
    .B1(net2230),
    .B2(net3280),
    .A2(net2278),
    .A1(net3014));
 sg13g2_a21oi_1 _08663_ (.A1(_03532_),
    .A2(_03533_),
    .Y(_03534_),
    .B1(net2261));
 sg13g2_nor4_1 _08664_ (.A(_03513_),
    .B(_03519_),
    .C(_03525_),
    .D(_03528_),
    .Y(_03535_));
 sg13g2_nor4_1 _08665_ (.A(_03516_),
    .B(_03522_),
    .C(_03531_),
    .D(_03534_),
    .Y(_03536_));
 sg13g2_a21oi_1 _08666_ (.A1(_03535_),
    .A2(_03536_),
    .Y(_00460_),
    .B1(net2384));
 sg13g2_a22oi_1 _08667_ (.Y(_03537_),
    .B1(net2142),
    .B2(net1628),
    .A2(net2186),
    .A1(net3097));
 sg13g2_a22oi_1 _08668_ (.Y(_03538_),
    .B1(net2229),
    .B2(net2977),
    .A2(net2276),
    .A1(net2679));
 sg13g2_a21oi_1 _08669_ (.A1(_03537_),
    .A2(_03538_),
    .Y(_03539_),
    .B1(net2083));
 sg13g2_a22oi_1 _08670_ (.Y(_03540_),
    .B1(net2142),
    .B2(net1613),
    .A2(net2186),
    .A1(net1609));
 sg13g2_a22oi_1 _08671_ (.Y(_03541_),
    .B1(net2232),
    .B2(net3077),
    .A2(net2279),
    .A1(\rf_ram.RAM[19][28] ));
 sg13g2_a21oi_1 _08672_ (.A1(_03540_),
    .A2(_03541_),
    .Y(_03542_),
    .B1(net2073));
 sg13g2_a22oi_1 _08673_ (.Y(_03543_),
    .B1(net2142),
    .B2(net2782),
    .A2(net2186),
    .A1(net2966));
 sg13g2_a22oi_1 _08674_ (.Y(_03544_),
    .B1(net2229),
    .B2(net1505),
    .A2(net2276),
    .A1(net1705));
 sg13g2_a21oi_1 _08675_ (.A1(_03543_),
    .A2(_03544_),
    .Y(_03545_),
    .B1(net2068));
 sg13g2_a22oi_1 _08676_ (.Y(_03546_),
    .B1(net2142),
    .B2(net1538),
    .A2(net2186),
    .A1(net1523));
 sg13g2_a22oi_1 _08677_ (.Y(_03547_),
    .B1(net2229),
    .B2(net2920),
    .A2(net2276),
    .A1(net3183));
 sg13g2_a21oi_1 _08678_ (.A1(_03546_),
    .A2(_03547_),
    .Y(_03548_),
    .B1(net2098));
 sg13g2_a22oi_1 _08679_ (.Y(_03549_),
    .B1(net2142),
    .B2(net1521),
    .A2(net2187),
    .A1(net2891));
 sg13g2_a22oi_1 _08680_ (.Y(_03550_),
    .B1(net2232),
    .B2(net1704),
    .A2(net2276),
    .A1(net3788));
 sg13g2_a21oi_1 _08681_ (.A1(_03549_),
    .A2(_03550_),
    .Y(_03551_),
    .B1(net2103));
 sg13g2_a22oi_1 _08682_ (.Y(_03552_),
    .B1(net2143),
    .B2(net1673),
    .A2(net2187),
    .A1(net3100));
 sg13g2_a22oi_1 _08683_ (.Y(_03553_),
    .B1(net2232),
    .B2(net2614),
    .A2(net2276),
    .A1(net2842));
 sg13g2_a21oi_1 _08684_ (.A1(_03552_),
    .A2(_03553_),
    .Y(_03554_),
    .B1(net2261));
 sg13g2_a22oi_1 _08685_ (.Y(_03555_),
    .B1(net2143),
    .B2(net2715),
    .A2(net2186),
    .A1(net1533));
 sg13g2_a22oi_1 _08686_ (.Y(_03556_),
    .B1(net2229),
    .B2(net2902),
    .A2(net2276),
    .A1(net1607));
 sg13g2_a21oi_1 _08687_ (.A1(_03555_),
    .A2(_03556_),
    .Y(_03557_),
    .B1(net2078));
 sg13g2_a22oi_1 _08688_ (.Y(_03558_),
    .B1(net2142),
    .B2(net1671),
    .A2(net2186),
    .A1(net2985));
 sg13g2_a22oi_1 _08689_ (.Y(_03559_),
    .B1(net2229),
    .B2(net2689),
    .A2(net2276),
    .A1(net2617));
 sg13g2_a21oi_1 _08690_ (.A1(_03558_),
    .A2(_03559_),
    .Y(_03560_),
    .B1(net2307));
 sg13g2_nor4_1 _08691_ (.A(_03539_),
    .B(_03545_),
    .C(_03551_),
    .D(_03557_),
    .Y(_03561_));
 sg13g2_nor4_1 _08692_ (.A(_03542_),
    .B(_03548_),
    .C(_03554_),
    .D(_03560_),
    .Y(_03562_));
 sg13g2_a21oi_1 _08693_ (.A1(_03561_),
    .A2(_03562_),
    .Y(_00461_),
    .B1(net2384));
 sg13g2_a22oi_1 _08694_ (.Y(_03563_),
    .B1(net2131),
    .B2(net3034),
    .A2(net2175),
    .A1(net3114));
 sg13g2_a22oi_1 _08695_ (.Y(_03564_),
    .B1(net2219),
    .B2(net2957),
    .A2(net2266),
    .A1(net2709));
 sg13g2_a21oi_1 _08696_ (.A1(_03563_),
    .A2(_03564_),
    .Y(_03565_),
    .B1(net2260));
 sg13g2_a22oi_1 _08697_ (.Y(_03566_),
    .B1(net2131),
    .B2(net3065),
    .A2(net2175),
    .A1(net3288));
 sg13g2_a22oi_1 _08698_ (.Y(_03567_),
    .B1(net2219),
    .B2(net1455),
    .A2(net2266),
    .A1(net2925));
 sg13g2_a21oi_1 _08699_ (.A1(_03566_),
    .A2(_03567_),
    .Y(_03568_),
    .B1(net2097));
 sg13g2_a22oi_1 _08700_ (.Y(_03569_),
    .B1(net2130),
    .B2(net2876),
    .A2(net2174),
    .A1(net2748));
 sg13g2_a22oi_1 _08701_ (.Y(_03570_),
    .B1(net2218),
    .B2(net2887),
    .A2(net2265),
    .A1(net3053));
 sg13g2_a21oi_1 _08702_ (.A1(_03569_),
    .A2(_03570_),
    .Y(_03571_),
    .B1(net2072));
 sg13g2_a22oi_1 _08703_ (.Y(_03572_),
    .B1(net2133),
    .B2(net1581),
    .A2(net2177),
    .A1(net1586));
 sg13g2_a22oi_1 _08704_ (.Y(_03573_),
    .B1(net2221),
    .B2(net1438),
    .A2(net2268),
    .A1(net2907));
 sg13g2_a21oi_1 _08705_ (.A1(_03572_),
    .A2(_03573_),
    .Y(_03574_),
    .B1(net2102));
 sg13g2_a22oi_1 _08706_ (.Y(_03575_),
    .B1(net2131),
    .B2(net1457),
    .A2(net2175),
    .A1(net3066));
 sg13g2_a22oi_1 _08707_ (.Y(_03576_),
    .B1(net2219),
    .B2(net3232),
    .A2(net2266),
    .A1(net3407));
 sg13g2_a21oi_1 _08708_ (.A1(_03575_),
    .A2(_03576_),
    .Y(_03577_),
    .B1(net2067));
 sg13g2_a22oi_1 _08709_ (.Y(_03578_),
    .B1(net2133),
    .B2(net1632),
    .A2(net2177),
    .A1(net2971));
 sg13g2_a22oi_1 _08710_ (.Y(_03579_),
    .B1(net2221),
    .B2(net2906),
    .A2(net2268),
    .A1(net1448));
 sg13g2_a21oi_1 _08711_ (.A1(_03578_),
    .A2(_03579_),
    .Y(_03580_),
    .B1(net2082));
 sg13g2_a22oi_1 _08712_ (.Y(_03581_),
    .B1(net2130),
    .B2(net2869),
    .A2(net2174),
    .A1(net1595));
 sg13g2_a22oi_1 _08713_ (.Y(_03582_),
    .B1(net2218),
    .B2(net2611),
    .A2(net2265),
    .A1(net3265));
 sg13g2_a21oi_1 _08714_ (.A1(_03581_),
    .A2(_03582_),
    .Y(_03583_),
    .B1(net2308));
 sg13g2_a22oi_1 _08715_ (.Y(_03584_),
    .B1(net2134),
    .B2(net3104),
    .A2(net2178),
    .A1(net3234));
 sg13g2_a22oi_1 _08716_ (.Y(_03585_),
    .B1(net2222),
    .B2(net1466),
    .A2(net2268),
    .A1(net2939));
 sg13g2_a21oi_1 _08717_ (.A1(_03584_),
    .A2(_03585_),
    .Y(_03586_),
    .B1(net2077));
 sg13g2_nor4_1 _08718_ (.A(_03565_),
    .B(_03571_),
    .C(_03577_),
    .D(_03583_),
    .Y(_03587_));
 sg13g2_nor4_1 _08719_ (.A(_03568_),
    .B(_03574_),
    .C(_03580_),
    .D(_03586_),
    .Y(_03588_));
 sg13g2_a21oi_1 _08720_ (.A1(_03587_),
    .A2(_03588_),
    .Y(_00462_),
    .B1(net2384));
 sg13g2_a22oi_1 _08721_ (.Y(_03589_),
    .B1(net2132),
    .B2(\rf_ram.RAM[30][30] ),
    .A2(net2176),
    .A1(\rf_ram.RAM[29][30] ));
 sg13g2_a22oi_1 _08722_ (.Y(_03590_),
    .B1(net2220),
    .B2(\rf_ram.RAM[28][30] ),
    .A2(net2267),
    .A1(\rf_ram.RAM[31][30] ));
 sg13g2_a21oi_1 _08723_ (.A1(_03589_),
    .A2(_03590_),
    .Y(_03591_),
    .B1(net2077));
 sg13g2_a22oi_1 _08724_ (.Y(_03592_),
    .B1(net2132),
    .B2(\rf_ram.RAM[10][30] ),
    .A2(net2179),
    .A1(\rf_ram.RAM[9][30] ));
 sg13g2_a22oi_1 _08725_ (.Y(_03593_),
    .B1(net2223),
    .B2(\rf_ram.RAM[8][30] ),
    .A2(net2270),
    .A1(\rf_ram.RAM[11][30] ));
 sg13g2_a21oi_1 _08726_ (.A1(_03592_),
    .A2(_03593_),
    .Y(_03594_),
    .B1(net2097));
 sg13g2_a22oi_1 _08727_ (.Y(_03595_),
    .B1(net2132),
    .B2(\rf_ram.RAM[2][30] ),
    .A2(net2176),
    .A1(\rf_ram.RAM[1][30] ));
 sg13g2_a22oi_1 _08728_ (.Y(_03596_),
    .B1(net2220),
    .B2(\rf_ram.RAM[0][30] ),
    .A2(net2267),
    .A1(\rf_ram.RAM[3][30] ));
 sg13g2_a21oi_1 _08729_ (.A1(_03595_),
    .A2(_03596_),
    .Y(_03597_),
    .B1(net2308));
 sg13g2_a22oi_1 _08730_ (.Y(_03598_),
    .B1(net2132),
    .B2(\rf_ram.RAM[22][30] ),
    .A2(net2176),
    .A1(\rf_ram.RAM[21][30] ));
 sg13g2_a22oi_1 _08731_ (.Y(_03599_),
    .B1(net2220),
    .B2(\rf_ram.RAM[20][30] ),
    .A2(net2267),
    .A1(\rf_ram.RAM[23][30] ));
 sg13g2_a21oi_1 _08732_ (.A1(_03598_),
    .A2(_03599_),
    .Y(_03600_),
    .B1(net2067));
 sg13g2_a22oi_1 _08733_ (.Y(_03601_),
    .B1(net2132),
    .B2(\rf_ram.RAM[14][30] ),
    .A2(net2176),
    .A1(\rf_ram.RAM[13][30] ));
 sg13g2_a22oi_1 _08734_ (.Y(_03602_),
    .B1(net2220),
    .B2(\rf_ram.RAM[12][30] ),
    .A2(net2267),
    .A1(\rf_ram.RAM[15][30] ));
 sg13g2_a21oi_1 _08735_ (.A1(_03601_),
    .A2(_03602_),
    .Y(_03603_),
    .B1(net2102));
 sg13g2_a22oi_1 _08736_ (.Y(_03604_),
    .B1(net2135),
    .B2(\rf_ram.RAM[18][30] ),
    .A2(net2176),
    .A1(\rf_ram.RAM[17][30] ));
 sg13g2_a22oi_1 _08737_ (.Y(_03605_),
    .B1(net2220),
    .B2(\rf_ram.RAM[16][30] ),
    .A2(net2267),
    .A1(\rf_ram.RAM[19][30] ));
 sg13g2_a21oi_1 _08738_ (.A1(_03604_),
    .A2(_03605_),
    .Y(_03606_),
    .B1(net2072));
 sg13g2_a22oi_1 _08739_ (.Y(_03607_),
    .B1(net2132),
    .B2(net1507),
    .A2(net2176),
    .A1(net3813));
 sg13g2_a22oi_1 _08740_ (.Y(_03608_),
    .B1(net2220),
    .B2(\rf_ram.RAM[24][30] ),
    .A2(net2267),
    .A1(\rf_ram.RAM[27][30] ));
 sg13g2_a21oi_1 _08741_ (.A1(_03607_),
    .A2(_03608_),
    .Y(_03609_),
    .B1(net2082));
 sg13g2_a22oi_1 _08742_ (.Y(_03610_),
    .B1(net2135),
    .B2(\rf_ram.RAM[6][30] ),
    .A2(net2179),
    .A1(\rf_ram.RAM[5][30] ));
 sg13g2_a22oi_1 _08743_ (.Y(_03611_),
    .B1(net2223),
    .B2(\rf_ram.RAM[4][30] ),
    .A2(net2270),
    .A1(\rf_ram.RAM[7][30] ));
 sg13g2_a21oi_1 _08744_ (.A1(_03610_),
    .A2(_03611_),
    .Y(_03612_),
    .B1(net2260));
 sg13g2_nor4_1 _08745_ (.A(_03591_),
    .B(_03597_),
    .C(_03603_),
    .D(net3814),
    .Y(_03613_));
 sg13g2_nor4_1 _08746_ (.A(_03594_),
    .B(_03600_),
    .C(_03606_),
    .D(_03612_),
    .Y(_03614_));
 sg13g2_a21oi_1 _08747_ (.A1(net3815),
    .A2(_03614_),
    .Y(_00463_),
    .B1(net2384));
 sg13g2_a22oi_1 _08748_ (.Y(_03615_),
    .B1(net2131),
    .B2(net3051),
    .A2(net2175),
    .A1(\rf_ram.RAM[21][31] ));
 sg13g2_a22oi_1 _08749_ (.Y(_03616_),
    .B1(net2219),
    .B2(net1470),
    .A2(net2266),
    .A1(\rf_ram.RAM[23][31] ));
 sg13g2_a21oi_1 _08750_ (.A1(_03615_),
    .A2(_03616_),
    .Y(_03617_),
    .B1(net2067));
 sg13g2_a22oi_1 _08751_ (.Y(_03618_),
    .B1(net2130),
    .B2(net2698),
    .A2(net2174),
    .A1(\rf_ram.RAM[25][31] ));
 sg13g2_a22oi_1 _08752_ (.Y(_03619_),
    .B1(net2218),
    .B2(net3209),
    .A2(net2265),
    .A1(\rf_ram.RAM[27][31] ));
 sg13g2_a21oi_1 _08753_ (.A1(_03618_),
    .A2(_03619_),
    .Y(_03620_),
    .B1(net2082));
 sg13g2_a22oi_1 _08754_ (.Y(_03621_),
    .B1(net2130),
    .B2(\rf_ram.RAM[6][31] ),
    .A2(net2174),
    .A1(\rf_ram.RAM[5][31] ));
 sg13g2_a22oi_1 _08755_ (.Y(_03622_),
    .B1(net2218),
    .B2(\rf_ram.RAM[4][31] ),
    .A2(net2265),
    .A1(\rf_ram.RAM[7][31] ));
 sg13g2_a21oi_1 _08756_ (.A1(_03621_),
    .A2(_03622_),
    .Y(_03623_),
    .B1(net2260));
 sg13g2_a22oi_1 _08757_ (.Y(_03624_),
    .B1(net2130),
    .B2(\rf_ram.RAM[10][31] ),
    .A2(net2174),
    .A1(\rf_ram.RAM[9][31] ));
 sg13g2_a22oi_1 _08758_ (.Y(_03625_),
    .B1(net2218),
    .B2(\rf_ram.RAM[8][31] ),
    .A2(net2265),
    .A1(\rf_ram.RAM[11][31] ));
 sg13g2_a21oi_1 _08759_ (.A1(_03624_),
    .A2(_03625_),
    .Y(_03626_),
    .B1(net2097));
 sg13g2_a22oi_1 _08760_ (.Y(_03627_),
    .B1(net2130),
    .B2(net2703),
    .A2(net2174),
    .A1(\rf_ram.RAM[1][31] ));
 sg13g2_a22oi_1 _08761_ (.Y(_03628_),
    .B1(net2218),
    .B2(net1478),
    .A2(net2265),
    .A1(net3803));
 sg13g2_a21oi_1 _08762_ (.A1(_03627_),
    .A2(_03628_),
    .Y(_03629_),
    .B1(net2308));
 sg13g2_a22oi_1 _08763_ (.Y(_03630_),
    .B1(net2130),
    .B2(\rf_ram.RAM[30][31] ),
    .A2(net2174),
    .A1(\rf_ram.RAM[29][31] ));
 sg13g2_a22oi_1 _08764_ (.Y(_03631_),
    .B1(net2218),
    .B2(\rf_ram.RAM[28][31] ),
    .A2(net2265),
    .A1(\rf_ram.RAM[31][31] ));
 sg13g2_a21oi_1 _08765_ (.A1(_03630_),
    .A2(_03631_),
    .Y(_03632_),
    .B1(net2077));
 sg13g2_a22oi_1 _08766_ (.Y(_03633_),
    .B1(net2131),
    .B2(net2639),
    .A2(net2175),
    .A1(net3126));
 sg13g2_a22oi_1 _08767_ (.Y(_03634_),
    .B1(net2219),
    .B2(net1668),
    .A2(net2266),
    .A1(\rf_ram.RAM[15][31] ));
 sg13g2_a21oi_1 _08768_ (.A1(_03633_),
    .A2(_03634_),
    .Y(_03635_),
    .B1(net2102));
 sg13g2_a22oi_1 _08769_ (.Y(_03636_),
    .B1(net2130),
    .B2(\rf_ram.RAM[18][31] ),
    .A2(net2174),
    .A1(\rf_ram.RAM[17][31] ));
 sg13g2_a22oi_1 _08770_ (.Y(_03637_),
    .B1(net2218),
    .B2(\rf_ram.RAM[16][31] ),
    .A2(net2265),
    .A1(\rf_ram.RAM[19][31] ));
 sg13g2_a21oi_1 _08771_ (.A1(_03636_),
    .A2(_03637_),
    .Y(_03638_),
    .B1(net2072));
 sg13g2_nor4_1 _08772_ (.A(_03617_),
    .B(_03620_),
    .C(net3804),
    .D(_03635_),
    .Y(_03639_));
 sg13g2_nor4_1 _08773_ (.A(_03623_),
    .B(_03626_),
    .C(_03632_),
    .D(_03638_),
    .Y(_03640_));
 sg13g2_a21oi_1 _08774_ (.A1(net3805),
    .A2(_03640_),
    .Y(_00464_),
    .B1(net2384));
 sg13g2_nor2_1 _08775_ (.A(_01334_),
    .B(_01484_),
    .Y(_03641_));
 sg13g2_nand3_1 _08776_ (.B(_01428_),
    .C(net2365),
    .A(net2598),
    .Y(_03642_));
 sg13g2_nand2_1 _08777_ (.Y(_03643_),
    .A(net2597),
    .B(_01428_));
 sg13g2_nor2_1 _08778_ (.A(net3609),
    .B(_03643_),
    .Y(_03644_));
 sg13g2_a21oi_1 _08779_ (.A1(net2342),
    .A2(_03642_),
    .Y(_00465_),
    .B1(_03644_));
 sg13g2_and2_1 _08780_ (.A(net2581),
    .B(net1415),
    .X(_00466_));
 sg13g2_and2_1 _08781_ (.A(net1415),
    .B(\cpu.rf_ram_if.rtrig0 ),
    .X(_00467_));
 sg13g2_and2_1 _08782_ (.A(net2597),
    .B(net1414),
    .X(_00468_));
 sg13g2_nand2_1 _08783_ (.Y(_03645_),
    .A(net2602),
    .B(net3755));
 sg13g2_a21oi_1 _08784_ (.A1(net3723),
    .A2(_02687_),
    .Y(_03646_),
    .B1(_03645_));
 sg13g2_or2_1 _08785_ (.X(_00469_),
    .B(_03646_),
    .A(net2348));
 sg13g2_a21oi_1 _08786_ (.A1(net3340),
    .A2(net3759),
    .Y(_03647_),
    .B1(net2349));
 sg13g2_o21ai_1 _08787_ (.B1(_03647_),
    .Y(_03648_),
    .A1(net3340),
    .A2(net3759));
 sg13g2_a21oi_1 _08788_ (.A1(_02682_),
    .A2(_03648_),
    .Y(_00470_),
    .B1(_01334_));
 sg13g2_nor4_1 _08789_ (.A(\cpu.cpu.immdec.gen_immdec_w_eq_1.imm11_7[0] ),
    .B(\cpu.cpu.immdec.gen_immdec_w_eq_1.imm11_7[1] ),
    .C(\cpu.cpu.immdec.gen_immdec_w_eq_1.imm11_7[2] ),
    .D(\cpu.cpu.immdec.gen_immdec_w_eq_1.imm11_7[4] ),
    .Y(_03649_));
 sg13g2_a21oi_2 _08790_ (.B1(net2578),
    .Y(_03650_),
    .A2(_01492_),
    .A1(_01423_));
 sg13g2_a21oi_1 _08791_ (.A1(_01367_),
    .A2(_03649_),
    .Y(_03651_),
    .B1(_03650_));
 sg13g2_nand3_1 _08792_ (.B(_01484_),
    .C(_03651_),
    .A(net3340),
    .Y(_03652_));
 sg13g2_o21ai_1 _08793_ (.B1(_03652_),
    .Y(_00472_),
    .A1(net3340),
    .A2(_01363_));
 sg13g2_nand2_1 _08794_ (.Y(_00473_),
    .A(net2994),
    .B(_01519_));
 sg13g2_o21ai_1 _08795_ (.B1(net2597),
    .Y(_03653_),
    .A1(net3492),
    .A2(\cpu.cpu.state.o_cnt[2] ));
 sg13g2_a21oi_1 _08796_ (.A1(net3492),
    .A2(\cpu.cpu.state.o_cnt[2] ),
    .Y(_00474_),
    .B1(_03653_));
 sg13g2_a21oi_1 _08797_ (.A1(net3492),
    .A2(\cpu.cpu.state.o_cnt[2] ),
    .Y(_03654_),
    .B1(net3697));
 sg13g2_nand2_1 _08798_ (.Y(_03655_),
    .A(net2597),
    .B(_01425_));
 sg13g2_nor2_1 _08799_ (.A(net3698),
    .B(_03655_),
    .Y(_00475_));
 sg13g2_a21oi_1 _08800_ (.A1(_01347_),
    .A2(_01425_),
    .Y(_00476_),
    .B1(_03643_));
 sg13g2_nand3_1 _08801_ (.B(net3489),
    .C(_01428_),
    .A(net2601),
    .Y(_03656_));
 sg13g2_or2_1 _08802_ (.X(_03657_),
    .B(_01478_),
    .A(net3571));
 sg13g2_or2_1 _08803_ (.X(_03658_),
    .B(net2568),
    .A(net2569));
 sg13g2_nand3b_1 _08804_ (.B(_03657_),
    .C(_01507_),
    .Y(_03659_),
    .A_N(_03658_));
 sg13g2_o21ai_1 _08805_ (.B1(net2569),
    .Y(_03660_),
    .A1(\cpu.cpu.bne_or_bge ),
    .A2(net2568));
 sg13g2_nand3_1 _08806_ (.B(_01510_),
    .C(_03660_),
    .A(_01509_),
    .Y(_03661_));
 sg13g2_o21ai_1 _08807_ (.B1(_03661_),
    .Y(_03662_),
    .A1(_01421_),
    .A2(_01445_));
 sg13g2_or3_1 _08808_ (.A(_01421_),
    .B(_01445_),
    .C(_03661_),
    .X(_03663_));
 sg13g2_nand3_1 _08809_ (.B(_03662_),
    .C(_03663_),
    .A(_03658_),
    .Y(_03664_));
 sg13g2_and3_1 _08810_ (.X(_03665_),
    .A(\cpu.cpu.bne_or_bge ),
    .B(_03659_),
    .C(_03664_));
 sg13g2_a21oi_1 _08811_ (.A1(_03659_),
    .A2(_03664_),
    .Y(_03666_),
    .B1(net3660));
 sg13g2_nor3_1 _08812_ (.A(net2580),
    .B(_03665_),
    .C(_03666_),
    .Y(_03667_));
 sg13g2_nand2_1 _08813_ (.Y(_03668_),
    .A(net2597),
    .B(_02675_));
 sg13g2_nand3_1 _08814_ (.B(net2572),
    .C(_02675_),
    .A(net2601),
    .Y(_03669_));
 sg13g2_o21ai_1 _08815_ (.B1(_03656_),
    .Y(_00477_),
    .A1(net3661),
    .A2(_03669_));
 sg13g2_o21ai_1 _08816_ (.B1(_03668_),
    .Y(_00478_),
    .A1(_01335_),
    .A2(_03643_));
 sg13g2_a21oi_1 _08817_ (.A1(net3492),
    .A2(_01426_),
    .Y(_03670_),
    .B1(net3532));
 sg13g2_a21oi_1 _08818_ (.A1(_02682_),
    .A2(net3533),
    .Y(_00479_),
    .B1(_01334_));
 sg13g2_and2_1 _08819_ (.A(net2597),
    .B(net3439),
    .X(_00480_));
 sg13g2_and2_1 _08820_ (.A(net2597),
    .B(net3364),
    .X(_00481_));
 sg13g2_and2_1 _08821_ (.A(net2597),
    .B(net3334),
    .X(_00482_));
 sg13g2_nor3_1 _08822_ (.A(\cpu.cpu.bufreg2.i_bytecnt[1] ),
    .B(\cpu.cpu.bufreg2.i_bytecnt[0] ),
    .C(_01458_),
    .Y(_03671_));
 sg13g2_nand2_1 _08823_ (.Y(_03672_),
    .A(_01457_),
    .B(_03671_));
 sg13g2_or2_1 _08824_ (.X(_03673_),
    .B(\cpu.cpu.bufreg2.i_bytecnt[1] ),
    .A(\cpu.cpu.bufreg.data[1] ));
 sg13g2_nand3_1 _08825_ (.B(\cpu.cpu.bufreg2.i_bytecnt[0] ),
    .C(_03673_),
    .A(\cpu.cpu.bufreg.data[0] ),
    .Y(_03674_));
 sg13g2_nand2_1 _08826_ (.Y(_03675_),
    .A(\cpu.cpu.bufreg.data[1] ),
    .B(\cpu.cpu.bufreg2.i_bytecnt[1] ));
 sg13g2_nand4_1 _08827_ (.B(_01458_),
    .C(_03674_),
    .A(_01418_),
    .Y(_03676_),
    .D(_03675_));
 sg13g2_nand3_1 _08828_ (.B(_03672_),
    .C(_03676_),
    .A(net2357),
    .Y(_03677_));
 sg13g2_nor2_1 _08829_ (.A(net3594),
    .B(net2395),
    .Y(_03678_));
 sg13g2_nor2_1 _08830_ (.A(net3721),
    .B(net2396),
    .Y(_03679_));
 sg13g2_nor3_1 _08831_ (.A(net2354),
    .B(_03678_),
    .C(_03679_),
    .Y(_03680_));
 sg13g2_a21oi_1 _08832_ (.A1(net3652),
    .A2(net2354),
    .Y(_03681_),
    .B1(_03680_));
 sg13g2_nor2_1 _08833_ (.A(net3612),
    .B(net2124),
    .Y(_03682_));
 sg13g2_a21oi_1 _08834_ (.A1(net2124),
    .A2(_03681_),
    .Y(_00483_),
    .B1(_03682_));
 sg13g2_nand2_1 _08835_ (.Y(_03683_),
    .A(net3658),
    .B(net2395));
 sg13g2_nand2_1 _08836_ (.Y(_03684_),
    .A(\cpu.arbiter.i_wb_mem_rdt[1] ),
    .B(_01653_));
 sg13g2_a21oi_1 _08837_ (.A1(_03683_),
    .A2(_03684_),
    .Y(_03685_),
    .B1(net2354));
 sg13g2_a21oi_1 _08838_ (.A1(net3576),
    .A2(net2355),
    .Y(_03686_),
    .B1(net3659));
 sg13g2_nor2_1 _08839_ (.A(net3652),
    .B(net2124),
    .Y(_03687_));
 sg13g2_a21oi_1 _08840_ (.A1(net2124),
    .A2(_03686_),
    .Y(_00484_),
    .B1(_03687_));
 sg13g2_nor2_1 _08841_ (.A(\cpu.arbiter.i_wb_mem_rdt[2] ),
    .B(net2395),
    .Y(_03688_));
 sg13g2_nor2_1 _08842_ (.A(\cpu.i_wb_ext_rdt[2] ),
    .B(net2396),
    .Y(_03689_));
 sg13g2_nor3_1 _08843_ (.A(net2355),
    .B(_03688_),
    .C(_03689_),
    .Y(_03690_));
 sg13g2_a21oi_1 _08844_ (.A1(\cpu.arbiter.i_wb_cpu_dbus_dat[3] ),
    .A2(net2355),
    .Y(_03691_),
    .B1(_03690_));
 sg13g2_nor2_1 _08845_ (.A(net3576),
    .B(net2124),
    .Y(_03692_));
 sg13g2_a21oi_1 _08846_ (.A1(net2124),
    .A2(_03691_),
    .Y(_00485_),
    .B1(_03692_));
 sg13g2_nor2_1 _08847_ (.A(\cpu.arbiter.i_wb_mem_rdt[3] ),
    .B(net2395),
    .Y(_03693_));
 sg13g2_nor2_1 _08848_ (.A(net3642),
    .B(net2396),
    .Y(_03694_));
 sg13g2_nor3_1 _08849_ (.A(net2354),
    .B(_03693_),
    .C(_03694_),
    .Y(_03695_));
 sg13g2_a21oi_1 _08850_ (.A1(net3635),
    .A2(net2354),
    .Y(_03696_),
    .B1(net3643));
 sg13g2_nor2_1 _08851_ (.A(net3621),
    .B(net2124),
    .Y(_03697_));
 sg13g2_a21oi_1 _08852_ (.A1(net2124),
    .A2(_03696_),
    .Y(_00486_),
    .B1(_03697_));
 sg13g2_nor2_1 _08853_ (.A(\cpu.arbiter.i_wb_mem_rdt[4] ),
    .B(net2395),
    .Y(_03698_));
 sg13g2_nor2_1 _08854_ (.A(\cpu.i_wb_ext_rdt[4] ),
    .B(net2396),
    .Y(_03699_));
 sg13g2_nor3_1 _08855_ (.A(net2354),
    .B(_03698_),
    .C(_03699_),
    .Y(_03700_));
 sg13g2_a21oi_1 _08856_ (.A1(\cpu.arbiter.i_wb_cpu_dbus_dat[5] ),
    .A2(net2356),
    .Y(_03701_),
    .B1(_03700_));
 sg13g2_nor2_1 _08857_ (.A(net3635),
    .B(net2123),
    .Y(_03702_));
 sg13g2_a21oi_1 _08858_ (.A1(net2123),
    .A2(_03701_),
    .Y(_00487_),
    .B1(_03702_));
 sg13g2_nor2_1 _08859_ (.A(net3678),
    .B(_01654_),
    .Y(_03703_));
 sg13g2_nor2_1 _08860_ (.A(\cpu.i_wb_ext_rdt[5] ),
    .B(net2396),
    .Y(_03704_));
 sg13g2_nor3_1 _08861_ (.A(net2354),
    .B(_03703_),
    .C(_03704_),
    .Y(_03705_));
 sg13g2_a21oi_1 _08862_ (.A1(net3632),
    .A2(net2356),
    .Y(_03706_),
    .B1(_03705_));
 sg13g2_nor2_1 _08863_ (.A(net3686),
    .B(net2123),
    .Y(_03707_));
 sg13g2_a21oi_1 _08864_ (.A1(net2123),
    .A2(_03706_),
    .Y(_00488_),
    .B1(_03707_));
 sg13g2_nor2_1 _08865_ (.A(\cpu.arbiter.i_wb_mem_rdt[6] ),
    .B(_01654_),
    .Y(_03708_));
 sg13g2_nor2_1 _08866_ (.A(\cpu.i_wb_ext_rdt[6] ),
    .B(net2396),
    .Y(_03709_));
 sg13g2_nor3_1 _08867_ (.A(net2354),
    .B(_03708_),
    .C(_03709_),
    .Y(_03710_));
 sg13g2_a21oi_1 _08868_ (.A1(\cpu.arbiter.i_wb_cpu_dbus_dat[7] ),
    .A2(net2356),
    .Y(_03711_),
    .B1(_03710_));
 sg13g2_nor2_1 _08869_ (.A(net3632),
    .B(net2123),
    .Y(_03712_));
 sg13g2_a21oi_1 _08870_ (.A1(net2123),
    .A2(_03711_),
    .Y(_00489_),
    .B1(_03712_));
 sg13g2_nor2_1 _08871_ (.A(\cpu.arbiter.i_wb_mem_rdt[7] ),
    .B(net2395),
    .Y(_03713_));
 sg13g2_nor2_1 _08872_ (.A(\cpu.i_wb_ext_rdt[7] ),
    .B(net2396),
    .Y(_03714_));
 sg13g2_nor3_1 _08873_ (.A(net2355),
    .B(_03713_),
    .C(_03714_),
    .Y(_03715_));
 sg13g2_a21oi_1 _08874_ (.A1(\cpu.arbiter.i_wb_cpu_dbus_dat[8] ),
    .A2(net2356),
    .Y(_03716_),
    .B1(_03715_));
 sg13g2_nor2_1 _08875_ (.A(net3648),
    .B(net2123),
    .Y(_03717_));
 sg13g2_a21oi_1 _08876_ (.A1(net2123),
    .A2(_03716_),
    .Y(_00490_),
    .B1(_03717_));
 sg13g2_nor3_2 _08877_ (.A(_01405_),
    .B(net2395),
    .C(net2393),
    .Y(_03718_));
 sg13g2_a22oi_1 _08878_ (.Y(_03719_),
    .B1(net2371),
    .B2(net3692),
    .A2(net2353),
    .A1(net3552));
 sg13g2_nor2_1 _08879_ (.A(net3738),
    .B(net2125),
    .Y(_03720_));
 sg13g2_a21oi_1 _08880_ (.A1(net2125),
    .A2(_03719_),
    .Y(_00491_),
    .B1(_03720_));
 sg13g2_a22oi_1 _08881_ (.Y(_03721_),
    .B1(net2371),
    .B2(\cpu.arbiter.i_wb_mem_rdt[9] ),
    .A2(net2353),
    .A1(net3546));
 sg13g2_nor2_1 _08882_ (.A(net3552),
    .B(net2122),
    .Y(_03722_));
 sg13g2_a21oi_1 _08883_ (.A1(net2122),
    .A2(_03721_),
    .Y(_00492_),
    .B1(_03722_));
 sg13g2_a22oi_1 _08884_ (.Y(_03723_),
    .B1(net2371),
    .B2(\cpu.arbiter.i_wb_mem_rdt[10] ),
    .A2(net2353),
    .A1(\cpu.arbiter.i_wb_cpu_dbus_dat[11] ));
 sg13g2_nor2_1 _08885_ (.A(net3546),
    .B(net2126),
    .Y(_03724_));
 sg13g2_a21oi_1 _08886_ (.A1(net2126),
    .A2(_03723_),
    .Y(_00493_),
    .B1(_03724_));
 sg13g2_a22oi_1 _08887_ (.Y(_03725_),
    .B1(net2370),
    .B2(\cpu.arbiter.i_wb_mem_rdt[11] ),
    .A2(net2351),
    .A1(net3548));
 sg13g2_nor2_1 _08888_ (.A(net3610),
    .B(net2118),
    .Y(_03726_));
 sg13g2_a21oi_1 _08889_ (.A1(net2118),
    .A2(_03725_),
    .Y(_00494_),
    .B1(_03726_));
 sg13g2_a22oi_1 _08890_ (.Y(_03727_),
    .B1(net2370),
    .B2(\cpu.arbiter.i_wb_mem_rdt[12] ),
    .A2(net2351),
    .A1(\cpu.arbiter.i_wb_cpu_dbus_dat[13] ));
 sg13g2_nor2_1 _08891_ (.A(net3548),
    .B(net2118),
    .Y(_03728_));
 sg13g2_a21oi_1 _08892_ (.A1(net2118),
    .A2(_03727_),
    .Y(_00495_),
    .B1(_03728_));
 sg13g2_a22oi_1 _08893_ (.Y(_03729_),
    .B1(net2370),
    .B2(\cpu.arbiter.i_wb_mem_rdt[13] ),
    .A2(net2351),
    .A1(\cpu.arbiter.i_wb_cpu_dbus_dat[14] ));
 sg13g2_nor2_1 _08894_ (.A(net3617),
    .B(net2118),
    .Y(_03730_));
 sg13g2_a21oi_1 _08895_ (.A1(net2118),
    .A2(_03729_),
    .Y(_00496_),
    .B1(_03730_));
 sg13g2_a22oi_1 _08896_ (.Y(_03731_),
    .B1(net2370),
    .B2(net3628),
    .A2(net2351),
    .A1(net3598));
 sg13g2_nor2_1 _08897_ (.A(net3639),
    .B(net2118),
    .Y(_03732_));
 sg13g2_a21oi_1 _08898_ (.A1(net2118),
    .A2(_03731_),
    .Y(_00497_),
    .B1(_03732_));
 sg13g2_a22oi_1 _08899_ (.Y(_03733_),
    .B1(_03718_),
    .B2(\cpu.arbiter.i_wb_mem_rdt[15] ),
    .A2(net2353),
    .A1(net3586));
 sg13g2_nor2_1 _08900_ (.A(net3598),
    .B(net2122),
    .Y(_03734_));
 sg13g2_a21oi_1 _08901_ (.A1(net2122),
    .A2(_03733_),
    .Y(_00498_),
    .B1(_03734_));
 sg13g2_a22oi_1 _08902_ (.Y(_03735_),
    .B1(net2370),
    .B2(net3494),
    .A2(net2352),
    .A1(net3588));
 sg13g2_nor2_1 _08903_ (.A(net3586),
    .B(net2122),
    .Y(_03736_));
 sg13g2_a21oi_1 _08904_ (.A1(net2121),
    .A2(_03735_),
    .Y(_00499_),
    .B1(_03736_));
 sg13g2_a22oi_1 _08905_ (.Y(_03737_),
    .B1(net2371),
    .B2(net3485),
    .A2(net2352),
    .A1(\cpu.arbiter.i_wb_cpu_dbus_dat[18] ));
 sg13g2_nor2_1 _08906_ (.A(net3588),
    .B(net2121),
    .Y(_03738_));
 sg13g2_a21oi_1 _08907_ (.A1(net2121),
    .A2(_03737_),
    .Y(_00500_),
    .B1(_03738_));
 sg13g2_a22oi_1 _08908_ (.Y(_03739_),
    .B1(net2370),
    .B2(net3565),
    .A2(net2352),
    .A1(net3580));
 sg13g2_nor2_1 _08909_ (.A(net3631),
    .B(net2120),
    .Y(_03740_));
 sg13g2_a21oi_1 _08910_ (.A1(net2120),
    .A2(_03739_),
    .Y(_00501_),
    .B1(_03740_));
 sg13g2_a22oi_1 _08911_ (.Y(_03741_),
    .B1(net2370),
    .B2(\cpu.arbiter.i_wb_mem_rdt[19] ),
    .A2(net2352),
    .A1(net3521));
 sg13g2_nor2_1 _08912_ (.A(net3580),
    .B(net2119),
    .Y(_03742_));
 sg13g2_a21oi_1 _08913_ (.A1(net2119),
    .A2(_03741_),
    .Y(_00502_),
    .B1(_03742_));
 sg13g2_a22oi_1 _08914_ (.Y(_03743_),
    .B1(net2369),
    .B2(\cpu.arbiter.i_wb_mem_rdt[20] ),
    .A2(net2353),
    .A1(net3519));
 sg13g2_nor2_1 _08915_ (.A(net3521),
    .B(net2119),
    .Y(_03744_));
 sg13g2_a21oi_1 _08916_ (.A1(net2119),
    .A2(_03743_),
    .Y(_00503_),
    .B1(_03744_));
 sg13g2_a22oi_1 _08917_ (.Y(_03745_),
    .B1(net2369),
    .B2(\cpu.arbiter.i_wb_mem_rdt[21] ),
    .A2(net2353),
    .A1(\cpu.arbiter.i_wb_cpu_dbus_dat[22] ));
 sg13g2_nor2_1 _08918_ (.A(net3519),
    .B(net2119),
    .Y(_03746_));
 sg13g2_a21oi_1 _08919_ (.A1(net2119),
    .A2(_03745_),
    .Y(_00504_),
    .B1(_03746_));
 sg13g2_a22oi_1 _08920_ (.Y(_03747_),
    .B1(net2369),
    .B2(\cpu.arbiter.i_wb_mem_rdt[22] ),
    .A2(net2352),
    .A1(\cpu.arbiter.i_wb_cpu_dbus_dat[23] ));
 sg13g2_nor2_1 _08921_ (.A(net3550),
    .B(net2120),
    .Y(_03748_));
 sg13g2_a21oi_1 _08922_ (.A1(net2120),
    .A2(_03747_),
    .Y(_00505_),
    .B1(_03748_));
 sg13g2_a22oi_1 _08923_ (.Y(_03749_),
    .B1(net2371),
    .B2(\cpu.arbiter.i_wb_mem_rdt[23] ),
    .A2(net2352),
    .A1(\cpu.arbiter.i_wb_cpu_dbus_dat[24] ));
 sg13g2_nor2_1 _08924_ (.A(net3650),
    .B(net2119),
    .Y(_03750_));
 sg13g2_a21oi_1 _08925_ (.A1(net2119),
    .A2(_03749_),
    .Y(_00506_),
    .B1(_03750_));
 sg13g2_mux2_1 _08926_ (.A0(net3716),
    .A1(net3637),
    .S(net2349),
    .X(_00507_));
 sg13g2_mux2_1 _08927_ (.A0(net3730),
    .A1(net3690),
    .S(net2349),
    .X(_00508_));
 sg13g2_nor2_1 _08928_ (.A(net3718),
    .B(net2365),
    .Y(_03751_));
 sg13g2_a21oi_1 _08929_ (.A1(_01345_),
    .A2(net2365),
    .Y(_00509_),
    .B1(_03751_));
 sg13g2_mux2_1 _08930_ (.A0(net2576),
    .A1(net3678),
    .S(net2349),
    .X(_00510_));
 sg13g2_mux2_1 _08931_ (.A0(net2574),
    .A1(net3683),
    .S(net2349),
    .X(_00511_));
 sg13g2_nand2_2 _08932_ (.Y(_03752_),
    .A(net3669),
    .B(net2345));
 sg13g2_o21ai_1 _08933_ (.B1(_03752_),
    .Y(_00512_),
    .A1(_01342_),
    .A2(net2350));
 sg13g2_and2_1 _08934_ (.A(net3694),
    .B(net2345),
    .X(_03753_));
 sg13g2_a21o_1 _08935_ (.A2(net2365),
    .A1(net2569),
    .B1(_03753_),
    .X(_00513_));
 sg13g2_and2_1 _08936_ (.A(net3628),
    .B(net2345),
    .X(_03754_));
 sg13g2_a21o_1 _08937_ (.A2(net2364),
    .A1(net2568),
    .B1(_03754_),
    .X(_00514_));
 sg13g2_and2_1 _08938_ (.A(net3558),
    .B(net2346),
    .X(_03755_));
 sg13g2_a21o_1 _08939_ (.A2(net2366),
    .A1(net3516),
    .B1(_03755_),
    .X(_00515_));
 sg13g2_a21oi_1 _08940_ (.A1(net2573),
    .A2(net2578),
    .Y(_03756_),
    .B1(_01423_));
 sg13g2_nor2_1 _08941_ (.A(net2566),
    .B(_03756_),
    .Y(_03757_));
 sg13g2_nor2_2 _08942_ (.A(net2346),
    .B(_03757_),
    .Y(_03758_));
 sg13g2_nor2b_2 _08943_ (.A(net2346),
    .B_N(_03757_),
    .Y(_03759_));
 sg13g2_a221oi_1 _08944_ (.B2(net3753),
    .C1(_03755_),
    .B1(_03759_),
    .A1(\cpu.cpu.immdec.gen_immdec_w_eq_1.imm24_20[0] ),
    .Y(_03760_),
    .A2(_03758_));
 sg13g2_inv_1 _08945_ (.Y(_00516_),
    .A(net3754));
 sg13g2_a22oi_1 _08946_ (.Y(_03761_),
    .B1(_03759_),
    .B2(\cpu.cpu.immdec.gen_immdec_w_eq_1.imm24_20[2] ),
    .A2(_03758_),
    .A1(\cpu.cpu.immdec.gen_immdec_w_eq_1.imm24_20[1] ));
 sg13g2_o21ai_1 _08947_ (.B1(_03761_),
    .Y(_00517_),
    .A1(_01359_),
    .A2(net2363));
 sg13g2_a22oi_1 _08948_ (.Y(_03762_),
    .B1(_03759_),
    .B2(net3701),
    .A2(_03758_),
    .A1(\cpu.cpu.immdec.gen_immdec_w_eq_1.imm24_20[2] ));
 sg13g2_o21ai_1 _08949_ (.B1(net3702),
    .Y(_00518_),
    .A1(_01360_),
    .A2(net2363));
 sg13g2_a22oi_1 _08950_ (.Y(_03763_),
    .B1(_03759_),
    .B2(net3719),
    .A2(_03758_),
    .A1(net3701));
 sg13g2_o21ai_1 _08951_ (.B1(_03763_),
    .Y(_00519_),
    .A1(_01353_),
    .A2(net2363));
 sg13g2_a22oi_1 _08952_ (.Y(_03764_),
    .B1(_03759_),
    .B2(net3696),
    .A2(_03758_),
    .A1(net3719));
 sg13g2_o21ai_1 _08953_ (.B1(_03764_),
    .Y(_00520_),
    .A1(_01361_),
    .A2(net2363));
 sg13g2_and4_1 _08954_ (.A(_01345_),
    .B(net2579),
    .C(_01487_),
    .D(net2365),
    .X(_03765_));
 sg13g2_a21oi_1 _08955_ (.A1(net2566),
    .A2(net2365),
    .Y(_03766_),
    .B1(_03765_));
 sg13g2_nor2b_1 _08956_ (.A(net2344),
    .B_N(net3398),
    .Y(_03767_));
 sg13g2_a21oi_1 _08957_ (.A1(net3556),
    .A2(net2344),
    .Y(_03768_),
    .B1(_03767_));
 sg13g2_nor2_1 _08958_ (.A(net3696),
    .B(net2315),
    .Y(_03769_));
 sg13g2_a21oi_1 _08959_ (.A1(net2315),
    .A2(_03768_),
    .Y(_00521_),
    .B1(_03769_));
 sg13g2_nor2b_1 _08960_ (.A(net2344),
    .B_N(net3362),
    .Y(_03770_));
 sg13g2_a21oi_1 _08961_ (.A1(\cpu.arbiter.i_wb_mem_rdt[26] ),
    .A2(net2344),
    .Y(_03771_),
    .B1(_03770_));
 sg13g2_nor2_1 _08962_ (.A(net3398),
    .B(net2314),
    .Y(_03772_));
 sg13g2_a21oi_1 _08963_ (.A1(net2314),
    .A2(_03771_),
    .Y(_00522_),
    .B1(_03772_));
 sg13g2_nor2b_1 _08964_ (.A(net2344),
    .B_N(\cpu.cpu.immdec.gen_immdec_w_eq_1.imm30_25[3] ),
    .Y(_03773_));
 sg13g2_a21oi_1 _08965_ (.A1(\cpu.arbiter.i_wb_mem_rdt[27] ),
    .A2(net2344),
    .Y(_03774_),
    .B1(_03773_));
 sg13g2_nor2_1 _08966_ (.A(net3362),
    .B(net2314),
    .Y(_03775_));
 sg13g2_a21oi_1 _08967_ (.A1(net2314),
    .A2(_03774_),
    .Y(_00523_),
    .B1(_03775_));
 sg13g2_nor2b_1 _08968_ (.A(net2344),
    .B_N(\cpu.cpu.immdec.gen_immdec_w_eq_1.imm30_25[4] ),
    .Y(_03776_));
 sg13g2_a21oi_1 _08969_ (.A1(\cpu.arbiter.i_wb_mem_rdt[28] ),
    .A2(net2344),
    .Y(_03777_),
    .B1(_03776_));
 sg13g2_nor2_1 _08970_ (.A(net3373),
    .B(net2314),
    .Y(_03778_));
 sg13g2_a21oi_1 _08971_ (.A1(net2314),
    .A2(_03777_),
    .Y(_00524_),
    .B1(_03778_));
 sg13g2_nor2b_1 _08972_ (.A(net2345),
    .B_N(net3420),
    .Y(_03779_));
 sg13g2_a21oi_1 _08973_ (.A1(\cpu.arbiter.i_wb_mem_rdt[29] ),
    .A2(net2345),
    .Y(_03780_),
    .B1(_03779_));
 sg13g2_nor2_1 _08974_ (.A(net3457),
    .B(net2314),
    .Y(_03781_));
 sg13g2_a21oi_1 _08975_ (.A1(net2314),
    .A2(_03780_),
    .Y(_00525_),
    .B1(_03781_));
 sg13g2_a21oi_1 _08976_ (.A1(net2577),
    .A2(net2579),
    .Y(_03782_),
    .B1(\cpu.cpu.decode.opcode[1] ));
 sg13g2_o21ai_1 _08977_ (.B1(_01474_),
    .Y(_03783_),
    .A1(\cpu.cpu.immdec.gen_immdec_w_eq_1.imm19_12_20[0] ),
    .A2(_03782_));
 sg13g2_a21oi_1 _08978_ (.A1(_01432_),
    .A2(_03782_),
    .Y(_03784_),
    .B1(_03783_));
 sg13g2_a21oi_1 _08979_ (.A1(net3254),
    .A2(_01473_),
    .Y(_03785_),
    .B1(_03784_));
 sg13g2_o21ai_1 _08980_ (.B1(net2315),
    .Y(_03786_),
    .A1(net2350),
    .A2(_03785_));
 sg13g2_a21oi_1 _08981_ (.A1(\cpu.arbiter.i_wb_mem_rdt[30] ),
    .A2(net2345),
    .Y(_03787_),
    .B1(_03786_));
 sg13g2_nor2_1 _08982_ (.A(net3420),
    .B(net2315),
    .Y(_03788_));
 sg13g2_nor2_1 _08983_ (.A(_03787_),
    .B(_03788_),
    .Y(_00526_));
 sg13g2_nor2_1 _08984_ (.A(_01432_),
    .B(net2348),
    .Y(_03789_));
 sg13g2_nand3_1 _08985_ (.B(net2566),
    .C(net2365),
    .A(net3254),
    .Y(_03790_));
 sg13g2_a22oi_1 _08986_ (.Y(_03791_),
    .B1(_03789_),
    .B2(_01418_),
    .A2(net2348),
    .A1(\cpu.arbiter.i_wb_mem_rdt[7] ));
 sg13g2_nand2_1 _08987_ (.Y(_00527_),
    .A(_03790_),
    .B(_03791_));
 sg13g2_o21ai_1 _08988_ (.B1(_01453_),
    .Y(_03792_),
    .A1(net2578),
    .A2(\cpu.cpu.decode.opcode[1] ));
 sg13g2_a21oi_1 _08989_ (.A1(_01431_),
    .A2(_03792_),
    .Y(_03793_),
    .B1(net2566));
 sg13g2_or2_1 _08990_ (.X(_03794_),
    .B(_03793_),
    .A(net2348));
 sg13g2_inv_1 _08991_ (.Y(_03795_),
    .A(net2313));
 sg13g2_a21oi_1 _08992_ (.A1(net3440),
    .A2(net2366),
    .Y(_03796_),
    .B1(_03755_));
 sg13g2_nor2_1 _08993_ (.A(net3510),
    .B(net2313),
    .Y(_03797_));
 sg13g2_a21oi_1 _08994_ (.A1(net2313),
    .A2(_03796_),
    .Y(_00528_),
    .B1(_03797_));
 sg13g2_a21oi_1 _08995_ (.A1(\cpu.cpu.immdec.gen_immdec_w_eq_1.imm19_12_20[2] ),
    .A2(net2363),
    .Y(_03798_),
    .B1(net2117));
 sg13g2_a22oi_1 _08996_ (.Y(_00529_),
    .B1(_03798_),
    .B2(_03752_),
    .A2(_03795_),
    .A1(_01369_));
 sg13g2_nor2_1 _08997_ (.A(net3487),
    .B(net2313),
    .Y(_03799_));
 sg13g2_a21oi_1 _08998_ (.A1(net3435),
    .A2(net2364),
    .Y(_03800_),
    .B1(_03753_));
 sg13g2_a21oi_1 _08999_ (.A1(net2313),
    .A2(_03800_),
    .Y(_00530_),
    .B1(_03799_));
 sg13g2_a21oi_1 _09000_ (.A1(net3418),
    .A2(net2363),
    .Y(_03801_),
    .B1(_03754_));
 sg13g2_nor2_1 _09001_ (.A(net3435),
    .B(net2313),
    .Y(_03802_));
 sg13g2_a21oi_1 _09002_ (.A1(_03794_),
    .A2(_03801_),
    .Y(_00531_),
    .B1(_03802_));
 sg13g2_nor2_1 _09003_ (.A(\cpu.cpu.immdec.gen_immdec_w_eq_1.imm19_12_20[5] ),
    .B(net2346),
    .Y(_03803_));
 sg13g2_o21ai_1 _09004_ (.B1(_03794_),
    .Y(_03804_),
    .A1(\cpu.arbiter.i_wb_mem_rdt[15] ),
    .A2(net2364));
 sg13g2_nand2_1 _09005_ (.Y(_03805_),
    .A(net3418),
    .B(net2117));
 sg13g2_o21ai_1 _09006_ (.B1(_03805_),
    .Y(_00532_),
    .A1(_03803_),
    .A2(_03804_));
 sg13g2_nand2_1 _09007_ (.Y(_03806_),
    .A(net3494),
    .B(net2347));
 sg13g2_a21oi_1 _09008_ (.A1(net3615),
    .A2(net2363),
    .Y(_03807_),
    .B1(net2117));
 sg13g2_a22oi_1 _09009_ (.Y(_00533_),
    .B1(_03806_),
    .B2(_03807_),
    .A2(net2117),
    .A1(_01364_));
 sg13g2_nand2_1 _09010_ (.Y(_03808_),
    .A(net3485),
    .B(net2346));
 sg13g2_a21oi_1 _09011_ (.A1(net3578),
    .A2(net2363),
    .Y(_03809_),
    .B1(net2117));
 sg13g2_a22oi_1 _09012_ (.Y(_00534_),
    .B1(_03808_),
    .B2(_03809_),
    .A2(net2117),
    .A1(_01366_));
 sg13g2_nor2_1 _09013_ (.A(net3578),
    .B(net2313),
    .Y(_03810_));
 sg13g2_nor2_1 _09014_ (.A(_01368_),
    .B(net2346),
    .Y(_03811_));
 sg13g2_a21oi_1 _09015_ (.A1(net3565),
    .A2(net2346),
    .Y(_03812_),
    .B1(_03811_));
 sg13g2_a21oi_1 _09016_ (.A1(net2313),
    .A2(_03812_),
    .Y(_00535_),
    .B1(_03810_));
 sg13g2_a21oi_1 _09017_ (.A1(net2573),
    .A2(_01432_),
    .Y(_03813_),
    .B1(net2348));
 sg13g2_o21ai_1 _09018_ (.B1(_03813_),
    .Y(_03814_),
    .A1(net2573),
    .A2(\cpu.cpu.immdec.gen_immdec_w_eq_1.imm24_20[0] ));
 sg13g2_a22oi_1 _09019_ (.Y(_03815_),
    .B1(net2117),
    .B2(net3623),
    .A2(net2346),
    .A1(\cpu.arbiter.i_wb_mem_rdt[19] ));
 sg13g2_o21ai_1 _09020_ (.B1(net3624),
    .Y(_00536_),
    .A1(net2117),
    .A2(_03814_));
 sg13g2_mux2_1 _09021_ (.A0(net3640),
    .A1(\cpu.arbiter.i_wb_mem_rdt[31] ),
    .S(net2348),
    .X(_00537_));
 sg13g2_mux2_1 _09022_ (.A0(\cpu.cpu.bufreg.i_sh_signed ),
    .A1(net3732),
    .S(net2350),
    .X(_00538_));
 sg13g2_a21oi_1 _09023_ (.A1(_03659_),
    .A2(_03664_),
    .Y(_03816_),
    .B1(net2566));
 sg13g2_a21o_1 _09024_ (.A2(net2567),
    .A1(net3571),
    .B1(_03816_),
    .X(_00539_));
 sg13g2_nor2_1 _09025_ (.A(net2368),
    .B(net2122),
    .Y(_03817_));
 sg13g2_nor2_1 _09026_ (.A(net3734),
    .B(net2367),
    .Y(_03818_));
 sg13g2_a21oi_1 _09027_ (.A1(net3751),
    .A2(net2367),
    .Y(_03819_),
    .B1(_03818_));
 sg13g2_a22oi_1 _09028_ (.Y(_03820_),
    .B1(_03819_),
    .B2(net2351),
    .A2(net2369),
    .A1(net3584));
 sg13g2_nand2_1 _09029_ (.Y(_03821_),
    .A(net3751),
    .B(net2065));
 sg13g2_o21ai_1 _09030_ (.B1(_03821_),
    .Y(_00540_),
    .A1(net2065),
    .A2(_03820_));
 sg13g2_xor2_1 _09031_ (.B(net3734),
    .A(\cpu.arbiter.i_wb_cpu_dbus_dat[24] ),
    .X(_03822_));
 sg13g2_o21ai_1 _09032_ (.B1(net2351),
    .Y(_03823_),
    .A1(\cpu.arbiter.i_wb_cpu_dbus_dat[26] ),
    .A2(net2367));
 sg13g2_a21o_1 _09033_ (.A2(_03822_),
    .A1(net2367),
    .B1(_03823_),
    .X(_03824_));
 sg13g2_a21oi_1 _09034_ (.A1(net3556),
    .A2(net2369),
    .Y(_03825_),
    .B1(net2065));
 sg13g2_a22oi_1 _09035_ (.Y(_00541_),
    .B1(_03824_),
    .B2(_03825_),
    .A2(net2065),
    .A1(_01350_));
 sg13g2_xnor2_1 _09036_ (.Y(_03826_),
    .A(_01348_),
    .B(_01462_));
 sg13g2_o21ai_1 _09037_ (.B1(net2351),
    .Y(_03827_),
    .A1(net3674),
    .A2(net2367));
 sg13g2_a21o_1 _09038_ (.A2(_03826_),
    .A1(net2367),
    .B1(_03827_),
    .X(_03828_));
 sg13g2_a21oi_1 _09039_ (.A1(net3536),
    .A2(net2369),
    .Y(_03829_),
    .B1(net2065));
 sg13g2_a22oi_1 _09040_ (.Y(_00542_),
    .B1(_03828_),
    .B2(_03829_),
    .A2(net2065),
    .A1(_01348_));
 sg13g2_o21ai_1 _09041_ (.B1(net3674),
    .Y(_03830_),
    .A1(\cpu.arbiter.i_wb_cpu_dbus_dat[26] ),
    .A2(_01462_));
 sg13g2_nor2b_1 _09042_ (.A(_01463_),
    .B_N(_03830_),
    .Y(_03831_));
 sg13g2_o21ai_1 _09043_ (.B1(net2351),
    .Y(_03832_),
    .A1(\cpu.arbiter.i_wb_cpu_dbus_dat[28] ),
    .A2(net2367));
 sg13g2_a21o_1 _09044_ (.A2(_03831_),
    .A1(net2367),
    .B1(_03832_),
    .X(_03833_));
 sg13g2_a21oi_1 _09045_ (.A1(net3602),
    .A2(net2369),
    .Y(_03834_),
    .B1(net2065));
 sg13g2_a22oi_1 _09046_ (.Y(_00543_),
    .B1(_03833_),
    .B2(_03834_),
    .A2(net2065),
    .A1(_01349_));
 sg13g2_xnor2_1 _09047_ (.Y(_03835_),
    .A(net3739),
    .B(_01463_));
 sg13g2_o21ai_1 _09048_ (.B1(net2352),
    .Y(_03836_),
    .A1(\cpu.arbiter.i_wb_cpu_dbus_dat[29] ),
    .A2(net2368));
 sg13g2_a21o_1 _09049_ (.A2(_03835_),
    .A1(net2368),
    .B1(_03836_),
    .X(_03837_));
 sg13g2_a21oi_1 _09050_ (.A1(net3613),
    .A2(net2369),
    .Y(_03838_),
    .B1(net2066));
 sg13g2_a22oi_1 _09051_ (.Y(_00544_),
    .B1(_03837_),
    .B2(_03838_),
    .A2(net2066),
    .A1(_01351_));
 sg13g2_nand4_1 _09052_ (.B(\cpu.cpu.state.o_cnt[2] ),
    .C(_01459_),
    .A(net3492),
    .Y(_03839_),
    .D(_03671_));
 sg13g2_nand3_1 _09053_ (.B(net2353),
    .C(_03839_),
    .A(_01467_),
    .Y(_03840_));
 sg13g2_a21oi_1 _09054_ (.A1(net3591),
    .A2(net2371),
    .Y(_03841_),
    .B1(net2066));
 sg13g2_a22oi_1 _09055_ (.Y(_00545_),
    .B1(_03840_),
    .B2(_03841_),
    .A2(net2066),
    .A1(_01352_));
 sg13g2_a22oi_1 _09056_ (.Y(_03842_),
    .B1(_03718_),
    .B2(\cpu.arbiter.i_wb_mem_rdt[30] ),
    .A2(_02680_),
    .A1(\cpu.arbiter.i_wb_cpu_dbus_dat[31] ));
 sg13g2_nand2_1 _09057_ (.Y(_03843_),
    .A(net3450),
    .B(net2066));
 sg13g2_o21ai_1 _09058_ (.B1(_03843_),
    .Y(_00546_),
    .A1(net2066),
    .A2(_03842_));
 sg13g2_a22oi_1 _09059_ (.Y(_03844_),
    .B1(net2371),
    .B2(\cpu.arbiter.i_wb_mem_rdt[31] ),
    .A2(net2357),
    .A1(_01441_));
 sg13g2_nand2_1 _09060_ (.Y(_03845_),
    .A(net3464),
    .B(net2066));
 sg13g2_o21ai_1 _09061_ (.B1(_03845_),
    .Y(_00547_),
    .A1(_03817_),
    .A2(_03844_));
 sg13g2_o21ai_1 _09062_ (.B1(_01477_),
    .Y(_03846_),
    .A1(\cpu.cpu.state.cnt_r[1] ),
    .A2(\cpu.cpu.state.cnt_r[0] ));
 sg13g2_nand2_1 _09063_ (.Y(_03847_),
    .A(net2376),
    .B(_03846_));
 sg13g2_o21ai_1 _09064_ (.B1(_03847_),
    .Y(_03848_),
    .A1(net2376),
    .A2(_01471_));
 sg13g2_nor2_1 _09065_ (.A(net3747),
    .B(_03848_),
    .Y(_03849_));
 sg13g2_a21oi_1 _09066_ (.A1(_01341_),
    .A2(_03848_),
    .Y(_00548_),
    .B1(_03849_));
 sg13g2_o21ai_1 _09067_ (.B1(_02804_),
    .Y(_03850_),
    .A1(_01355_),
    .A2(net2376));
 sg13g2_mux2_1 _09068_ (.A0(_03850_),
    .A1(net3747),
    .S(_03848_),
    .X(_00549_));
 sg13g2_nand2_1 _09069_ (.Y(_03851_),
    .A(_01713_),
    .B(_01751_));
 sg13g2_nand2_1 _09070_ (.Y(_03852_),
    .A(net3144),
    .B(net1749));
 sg13g2_o21ai_1 _09071_ (.B1(_03852_),
    .Y(_00550_),
    .A1(net2564),
    .A2(net1749));
 sg13g2_nand2_1 _09072_ (.Y(_03853_),
    .A(net1418),
    .B(net1752));
 sg13g2_o21ai_1 _09073_ (.B1(_03853_),
    .Y(_00551_),
    .A1(net2556),
    .A2(net1752));
 sg13g2_nand2_1 _09074_ (.Y(_03854_),
    .A(net1619),
    .B(net1758));
 sg13g2_o21ai_1 _09075_ (.B1(_03854_),
    .Y(_00552_),
    .A1(net2550),
    .A2(net1758));
 sg13g2_nand2_1 _09076_ (.Y(_03855_),
    .A(net3087),
    .B(net1756));
 sg13g2_o21ai_1 _09077_ (.B1(_03855_),
    .Y(_00553_),
    .A1(net2544),
    .A2(net1756));
 sg13g2_nand2_1 _09078_ (.Y(_03856_),
    .A(net1600),
    .B(net1756));
 sg13g2_o21ai_1 _09079_ (.B1(_03856_),
    .Y(_00554_),
    .A1(net2540),
    .A2(net1756));
 sg13g2_nand2_1 _09080_ (.Y(_03857_),
    .A(net2642),
    .B(net1756));
 sg13g2_o21ai_1 _09081_ (.B1(_03857_),
    .Y(_00555_),
    .A1(net2533),
    .A2(net1756));
 sg13g2_nand2_1 _09082_ (.Y(_03858_),
    .A(net1519),
    .B(net1758));
 sg13g2_o21ai_1 _09083_ (.B1(_03858_),
    .Y(_00556_),
    .A1(net2528),
    .A2(net1757));
 sg13g2_nand2_1 _09084_ (.Y(_03859_),
    .A(net2837),
    .B(net1757));
 sg13g2_o21ai_1 _09085_ (.B1(_03859_),
    .Y(_00557_),
    .A1(net2523),
    .A2(net1757));
 sg13g2_nand2_1 _09086_ (.Y(_03860_),
    .A(net3043),
    .B(net1757));
 sg13g2_o21ai_1 _09087_ (.B1(_03860_),
    .Y(_00558_),
    .A1(net2518),
    .A2(net1757));
 sg13g2_nand2_1 _09088_ (.Y(_03861_),
    .A(net1490),
    .B(net1755));
 sg13g2_o21ai_1 _09089_ (.B1(_03861_),
    .Y(_00559_),
    .A1(net2512),
    .A2(net1755));
 sg13g2_nand2_1 _09090_ (.Y(_03862_),
    .A(net1441),
    .B(net1754));
 sg13g2_o21ai_1 _09091_ (.B1(_03862_),
    .Y(_00560_),
    .A1(net2507),
    .A2(net1754));
 sg13g2_nand2_1 _09092_ (.Y(_03863_),
    .A(net3056),
    .B(net1755));
 sg13g2_o21ai_1 _09093_ (.B1(_03863_),
    .Y(_00561_),
    .A1(net2504),
    .A2(net1755));
 sg13g2_nand2_1 _09094_ (.Y(_03864_),
    .A(net1559),
    .B(net1755));
 sg13g2_o21ai_1 _09095_ (.B1(_03864_),
    .Y(_00562_),
    .A1(net2498),
    .A2(net1755));
 sg13g2_nand2_1 _09096_ (.Y(_03865_),
    .A(net3085),
    .B(net1757));
 sg13g2_o21ai_1 _09097_ (.B1(_03865_),
    .Y(_00563_),
    .A1(net2494),
    .A2(net1757));
 sg13g2_nand2_1 _09098_ (.Y(_03866_),
    .A(net2904),
    .B(net1750));
 sg13g2_o21ai_1 _09099_ (.B1(_03866_),
    .Y(_00564_),
    .A1(net2487),
    .A2(net1750));
 sg13g2_nand2_1 _09100_ (.Y(_03867_),
    .A(net2722),
    .B(net1754));
 sg13g2_o21ai_1 _09101_ (.B1(_03867_),
    .Y(_00565_),
    .A1(net2484),
    .A2(net1754));
 sg13g2_nand2_1 _09102_ (.Y(_03868_),
    .A(net3140),
    .B(net1756));
 sg13g2_o21ai_1 _09103_ (.B1(_03868_),
    .Y(_00566_),
    .A1(net2479),
    .A2(net1756));
 sg13g2_nand2_1 _09104_ (.Y(_03869_),
    .A(net1497),
    .B(net1754));
 sg13g2_o21ai_1 _09105_ (.B1(_03869_),
    .Y(_00567_),
    .A1(net2472),
    .A2(net1754));
 sg13g2_nand2_1 _09106_ (.Y(_03870_),
    .A(net2856),
    .B(net1754));
 sg13g2_o21ai_1 _09107_ (.B1(_03870_),
    .Y(_00568_),
    .A1(net2466),
    .A2(net1754));
 sg13g2_nand2_1 _09108_ (.Y(_03871_),
    .A(net2638),
    .B(net1750));
 sg13g2_o21ai_1 _09109_ (.B1(_03871_),
    .Y(_00569_),
    .A1(net2462),
    .A2(net1750));
 sg13g2_nand2_1 _09110_ (.Y(_03872_),
    .A(net2976),
    .B(net1750));
 sg13g2_o21ai_1 _09111_ (.B1(_03872_),
    .Y(_00570_),
    .A1(net2457),
    .A2(net1750));
 sg13g2_nand2_1 _09112_ (.Y(_03873_),
    .A(net1535),
    .B(net1752));
 sg13g2_o21ai_1 _09113_ (.B1(_03873_),
    .Y(_00571_),
    .A1(net2450),
    .A2(net1752));
 sg13g2_nand2_1 _09114_ (.Y(_03874_),
    .A(net2674),
    .B(net1758));
 sg13g2_o21ai_1 _09115_ (.B1(_03874_),
    .Y(_00572_),
    .A1(net2446),
    .A2(net1758));
 sg13g2_nand2_1 _09116_ (.Y(_03875_),
    .A(net3035),
    .B(net1752));
 sg13g2_o21ai_1 _09117_ (.B1(_03875_),
    .Y(_00573_),
    .A1(net2440),
    .A2(net1752));
 sg13g2_nand2_1 _09118_ (.Y(_03876_),
    .A(net2759),
    .B(net1758));
 sg13g2_o21ai_1 _09119_ (.B1(_03876_),
    .Y(_00574_),
    .A1(net2434),
    .A2(net1758));
 sg13g2_nand2_1 _09120_ (.Y(_03877_),
    .A(net1536),
    .B(net1751));
 sg13g2_o21ai_1 _09121_ (.B1(_03877_),
    .Y(_00575_),
    .A1(net2428),
    .A2(net1751));
 sg13g2_nand2_1 _09122_ (.Y(_03878_),
    .A(net2849),
    .B(net1751));
 sg13g2_o21ai_1 _09123_ (.B1(_03878_),
    .Y(_00576_),
    .A1(net2423),
    .A2(net1751));
 sg13g2_nand2_1 _09124_ (.Y(_03879_),
    .A(net1579),
    .B(net1751));
 sg13g2_o21ai_1 _09125_ (.B1(_03879_),
    .Y(_00577_),
    .A1(net2418),
    .A2(net1751));
 sg13g2_nand2_1 _09126_ (.Y(_03880_),
    .A(net1538),
    .B(net1751));
 sg13g2_o21ai_1 _09127_ (.B1(_03880_),
    .Y(_00578_),
    .A1(net2413),
    .A2(net1751));
 sg13g2_nand2_1 _09128_ (.Y(_03881_),
    .A(net3065),
    .B(net1749));
 sg13g2_o21ai_1 _09129_ (.B1(_03881_),
    .Y(_00579_),
    .A1(net2409),
    .A2(net1749));
 sg13g2_nand2_1 _09130_ (.Y(_03882_),
    .A(net1622),
    .B(net1749));
 sg13g2_o21ai_1 _09131_ (.B1(_03882_),
    .Y(_00580_),
    .A1(net2403),
    .A2(net1749));
 sg13g2_nand2_1 _09132_ (.Y(_03883_),
    .A(net1676),
    .B(net1749));
 sg13g2_o21ai_1 _09133_ (.B1(_03883_),
    .Y(_00581_),
    .A1(net2398),
    .A2(net1749));
 sg13g2_nor2_1 _09134_ (.A(_01334_),
    .B(_01485_),
    .Y(_03884_));
 sg13g2_a22oi_1 _09135_ (.Y(_03885_),
    .B1(net2336),
    .B2(net3472),
    .A2(net2342),
    .A1(\cpu.cpu.ctrl.pc [0]));
 sg13g2_inv_1 _09136_ (.Y(_00582_),
    .A(net3473));
 sg13g2_a22oi_1 _09137_ (.Y(_03886_),
    .B1(net2337),
    .B2(net3544),
    .A2(net2343),
    .A1(net3472));
 sg13g2_inv_1 _09138_ (.Y(_00583_),
    .A(_03886_));
 sg13g2_a22oi_1 _09139_ (.Y(_03887_),
    .B1(net2337),
    .B2(net3534),
    .A2(net2342),
    .A1(\cpu.arbiter.i_wb_cpu_ibus_adr[2] ));
 sg13g2_inv_1 _09140_ (.Y(_00584_),
    .A(net3535));
 sg13g2_a22oi_1 _09141_ (.Y(_03888_),
    .B1(net2336),
    .B2(net3630),
    .A2(net2342),
    .A1(net3534));
 sg13g2_inv_1 _09142_ (.Y(_00585_),
    .A(_03888_));
 sg13g2_a22oi_1 _09143_ (.Y(_03889_),
    .B1(net2336),
    .B2(net3634),
    .A2(net2342),
    .A1(net3630));
 sg13g2_inv_1 _09144_ (.Y(_00586_),
    .A(_03889_));
 sg13g2_a22oi_1 _09145_ (.Y(_03890_),
    .B1(net2336),
    .B2(net3596),
    .A2(net2342),
    .A1(\cpu.arbiter.i_wb_cpu_ibus_adr[5] ));
 sg13g2_inv_1 _09146_ (.Y(_00587_),
    .A(net3597));
 sg13g2_a22oi_1 _09147_ (.Y(_03891_),
    .B1(net2336),
    .B2(net3500),
    .A2(net2343),
    .A1(\cpu.arbiter.i_wb_cpu_ibus_adr[6] ));
 sg13g2_inv_1 _09148_ (.Y(_00588_),
    .A(net3501));
 sg13g2_a22oi_1 _09149_ (.Y(_03892_),
    .B1(net2337),
    .B2(net3527),
    .A2(net2343),
    .A1(net3500));
 sg13g2_inv_1 _09150_ (.Y(_00589_),
    .A(_03892_));
 sg13g2_a22oi_1 _09151_ (.Y(_03893_),
    .B1(net2336),
    .B2(net3666),
    .A2(net2342),
    .A1(net3527));
 sg13g2_inv_1 _09152_ (.Y(_00590_),
    .A(_03893_));
 sg13g2_a22oi_1 _09153_ (.Y(_03894_),
    .B1(net2336),
    .B2(net3569),
    .A2(net2342),
    .A1(\cpu.arbiter.i_wb_cpu_ibus_adr[9] ));
 sg13g2_inv_1 _09154_ (.Y(_00591_),
    .A(net3570));
 sg13g2_a22oi_1 _09155_ (.Y(_03895_),
    .B1(net2335),
    .B2(net3567),
    .A2(net2341),
    .A1(\cpu.arbiter.i_wb_cpu_ibus_adr[10] ));
 sg13g2_inv_1 _09156_ (.Y(_00592_),
    .A(net3568));
 sg13g2_a22oi_1 _09157_ (.Y(_03896_),
    .B1(net2335),
    .B2(net3542),
    .A2(net2341),
    .A1(\cpu.arbiter.i_wb_cpu_ibus_adr[11] ));
 sg13g2_inv_1 _09158_ (.Y(_00593_),
    .A(net3543));
 sg13g2_a22oi_1 _09159_ (.Y(_03897_),
    .B1(net2335),
    .B2(net3490),
    .A2(net2341),
    .A1(\cpu.arbiter.i_wb_cpu_ibus_adr[12] ));
 sg13g2_inv_1 _09160_ (.Y(_00594_),
    .A(net3491));
 sg13g2_a22oi_1 _09161_ (.Y(_03898_),
    .B1(net2334),
    .B2(net3479),
    .A2(net2341),
    .A1(\cpu.arbiter.i_wb_cpu_ibus_adr[13] ));
 sg13g2_inv_1 _09162_ (.Y(_00595_),
    .A(net3480));
 sg13g2_a22oi_1 _09163_ (.Y(_03899_),
    .B1(net2334),
    .B2(net3608),
    .A2(net2341),
    .A1(net3479));
 sg13g2_inv_1 _09164_ (.Y(_00596_),
    .A(_03899_));
 sg13g2_a22oi_1 _09165_ (.Y(_03900_),
    .B1(net2333),
    .B2(net3455),
    .A2(net2340),
    .A1(\cpu.arbiter.i_wb_cpu_ibus_adr[15] ));
 sg13g2_inv_1 _09166_ (.Y(_00597_),
    .A(net3456));
 sg13g2_a22oi_1 _09167_ (.Y(_03901_),
    .B1(net2333),
    .B2(net3325),
    .A2(net2339),
    .A1(\cpu.arbiter.i_wb_cpu_ibus_adr[16] ));
 sg13g2_inv_1 _09168_ (.Y(_00598_),
    .A(net3326));
 sg13g2_a22oi_1 _09169_ (.Y(_03902_),
    .B1(net2333),
    .B2(net3429),
    .A2(net2339),
    .A1(net3325));
 sg13g2_inv_1 _09170_ (.Y(_00599_),
    .A(_03902_));
 sg13g2_a22oi_1 _09171_ (.Y(_03903_),
    .B1(net2332),
    .B2(net3380),
    .A2(net2339),
    .A1(\cpu.arbiter.i_wb_cpu_ibus_adr[18] ));
 sg13g2_inv_1 _09172_ (.Y(_00600_),
    .A(net3381));
 sg13g2_a22oi_1 _09173_ (.Y(_03904_),
    .B1(net2334),
    .B2(net3518),
    .A2(net2339),
    .A1(net3380));
 sg13g2_inv_1 _09174_ (.Y(_00601_),
    .A(_03904_));
 sg13g2_a22oi_1 _09175_ (.Y(_03905_),
    .B1(net2332),
    .B2(net3474),
    .A2(net2338),
    .A1(\cpu.arbiter.i_wb_cpu_ibus_adr[20] ));
 sg13g2_inv_1 _09176_ (.Y(_00602_),
    .A(net3475));
 sg13g2_a22oi_1 _09177_ (.Y(_03906_),
    .B1(net2332),
    .B2(net3481),
    .A2(net2338),
    .A1(net3474));
 sg13g2_inv_1 _09178_ (.Y(_00603_),
    .A(_03906_));
 sg13g2_a22oi_1 _09179_ (.Y(_03907_),
    .B1(net2332),
    .B2(net3314),
    .A2(net2338),
    .A1(\cpu.arbiter.i_wb_cpu_ibus_adr[22] ));
 sg13g2_inv_1 _09180_ (.Y(_00604_),
    .A(net3315));
 sg13g2_a22oi_1 _09181_ (.Y(_03908_),
    .B1(net2333),
    .B2(net3400),
    .A2(net2340),
    .A1(net3314));
 sg13g2_inv_1 _09182_ (.Y(_00605_),
    .A(_03908_));
 sg13g2_a22oi_1 _09183_ (.Y(_03909_),
    .B1(net2333),
    .B2(net3484),
    .A2(net2340),
    .A1(net3400));
 sg13g2_inv_1 _09184_ (.Y(_00606_),
    .A(_03909_));
 sg13g2_a22oi_1 _09185_ (.Y(_03910_),
    .B1(net2333),
    .B2(net3367),
    .A2(net2340),
    .A1(\cpu.arbiter.i_wb_cpu_ibus_adr[25] ));
 sg13g2_inv_1 _09186_ (.Y(_00607_),
    .A(net3368));
 sg13g2_a22oi_1 _09187_ (.Y(_03911_),
    .B1(net2333),
    .B2(net3454),
    .A2(net2340),
    .A1(net3367));
 sg13g2_inv_1 _09188_ (.Y(_00608_),
    .A(_03911_));
 sg13g2_a22oi_1 _09189_ (.Y(_03912_),
    .B1(net2332),
    .B2(net3437),
    .A2(net2338),
    .A1(\cpu.arbiter.i_wb_cpu_ibus_adr[27] ));
 sg13g2_inv_1 _09190_ (.Y(_00609_),
    .A(net3438));
 sg13g2_a22oi_1 _09191_ (.Y(_03913_),
    .B1(net2332),
    .B2(net3382),
    .A2(net2338),
    .A1(\cpu.arbiter.i_wb_cpu_ibus_adr[28] ));
 sg13g2_inv_1 _09192_ (.Y(_00610_),
    .A(net3383));
 sg13g2_a22oi_1 _09193_ (.Y(_03914_),
    .B1(net2332),
    .B2(net3386),
    .A2(net2338),
    .A1(net3382));
 sg13g2_inv_1 _09194_ (.Y(_00611_),
    .A(_03914_));
 sg13g2_a22oi_1 _09195_ (.Y(_03915_),
    .B1(net2332),
    .B2(net3426),
    .A2(net2338),
    .A1(net3386));
 sg13g2_inv_1 _09196_ (.Y(_00612_),
    .A(_03915_));
 sg13g2_o21ai_1 _09197_ (.B1(net2336),
    .Y(_03916_),
    .A1(net3489),
    .A2(_01521_));
 sg13g2_a21oi_2 _09198_ (.B1(_03916_),
    .Y(_03917_),
    .A2(_01504_),
    .A1(net3489));
 sg13g2_a21o_1 _09199_ (.A2(net2338),
    .A1(net3426),
    .B1(_03917_),
    .X(_00613_));
 sg13g2_and3_2 _09200_ (.X(_03918_),
    .A(_01418_),
    .B(net2365),
    .C(_03650_));
 sg13g2_a21oi_2 _09201_ (.B1(net2348),
    .Y(_03919_),
    .A2(_03650_),
    .A1(_01418_));
 sg13g2_nand2_1 _09202_ (.Y(_03920_),
    .A(net3477),
    .B(_03919_));
 sg13g2_a22oi_1 _09203_ (.Y(_03921_),
    .B1(_03918_),
    .B2(\cpu.cpu.immdec.gen_immdec_w_eq_1.imm11_7[1] ),
    .A2(net2348),
    .A1(\cpu.arbiter.i_wb_mem_rdt[7] ));
 sg13g2_nand2_1 _09204_ (.Y(_00614_),
    .A(_03920_),
    .B(_03921_));
 sg13g2_nand2b_1 _09205_ (.Y(_03922_),
    .B(_03918_),
    .A_N(\cpu.cpu.immdec.gen_immdec_w_eq_1.imm11_7[2] ));
 sg13g2_o21ai_1 _09206_ (.B1(_03922_),
    .Y(_03923_),
    .A1(\cpu.arbiter.i_wb_mem_rdt[8] ),
    .A2(net2364));
 sg13g2_a21oi_1 _09207_ (.A1(_01365_),
    .A2(_03919_),
    .Y(_00615_),
    .B1(_03923_));
 sg13g2_a22oi_1 _09208_ (.Y(_03924_),
    .B1(_03919_),
    .B2(net3709),
    .A2(_03918_),
    .A1(\cpu.cpu.immdec.gen_immdec_w_eq_1.imm11_7[3] ));
 sg13g2_o21ai_1 _09209_ (.B1(net3710),
    .Y(_00616_),
    .A1(_01356_),
    .A2(net2364));
 sg13g2_a22oi_1 _09210_ (.Y(_03925_),
    .B1(_03919_),
    .B2(net3714),
    .A2(_03918_),
    .A1(\cpu.cpu.immdec.gen_immdec_w_eq_1.imm11_7[4] ));
 sg13g2_o21ai_1 _09211_ (.B1(net3715),
    .Y(_00617_),
    .A1(_01357_),
    .A2(net2364));
 sg13g2_a22oi_1 _09212_ (.Y(_03926_),
    .B1(_03919_),
    .B2(net3722),
    .A2(_03918_),
    .A1(net3696));
 sg13g2_o21ai_1 _09213_ (.B1(_03926_),
    .Y(_00618_),
    .A1(_01358_),
    .A2(net2364));
 sg13g2_dfrbpq_1 _09214_ (.RESET_B(net82),
    .D(net3033),
    .Q(\rf_ram.RAM[3][0] ),
    .CLK(clknet_leaf_14_clk_regs));
 sg13g2_dfrbpq_1 _09215_ (.RESET_B(net675),
    .D(_00621_),
    .Q(\rf_ram.RAM[3][1] ),
    .CLK(clknet_leaf_72_clk_regs));
 sg13g2_dfrbpq_1 _09216_ (.RESET_B(net674),
    .D(_00622_),
    .Q(\rf_ram.RAM[3][2] ),
    .CLK(clknet_leaf_76_clk_regs));
 sg13g2_dfrbpq_1 _09217_ (.RESET_B(net673),
    .D(_00623_),
    .Q(\rf_ram.RAM[3][3] ),
    .CLK(clknet_leaf_78_clk_regs));
 sg13g2_dfrbpq_1 _09218_ (.RESET_B(net672),
    .D(_00624_),
    .Q(\rf_ram.RAM[3][4] ),
    .CLK(clknet_leaf_82_clk_regs));
 sg13g2_dfrbpq_1 _09219_ (.RESET_B(net671),
    .D(_00625_),
    .Q(\rf_ram.RAM[3][5] ),
    .CLK(clknet_leaf_81_clk_regs));
 sg13g2_dfrbpq_1 _09220_ (.RESET_B(net670),
    .D(_00626_),
    .Q(\rf_ram.RAM[3][6] ),
    .CLK(clknet_leaf_101_clk_regs));
 sg13g2_dfrbpq_1 _09221_ (.RESET_B(net669),
    .D(_00627_),
    .Q(\rf_ram.RAM[3][7] ),
    .CLK(clknet_leaf_100_clk_regs));
 sg13g2_dfrbpq_1 _09222_ (.RESET_B(net668),
    .D(_00628_),
    .Q(\rf_ram.RAM[3][8] ),
    .CLK(clknet_leaf_111_clk_regs));
 sg13g2_dfrbpq_1 _09223_ (.RESET_B(net667),
    .D(_00629_),
    .Q(\rf_ram.RAM[3][9] ),
    .CLK(clknet_leaf_128_clk_regs));
 sg13g2_dfrbpq_1 _09224_ (.RESET_B(net666),
    .D(_00630_),
    .Q(\rf_ram.RAM[3][10] ),
    .CLK(clknet_leaf_120_clk_regs));
 sg13g2_dfrbpq_1 _09225_ (.RESET_B(net665),
    .D(_00631_),
    .Q(\rf_ram.RAM[3][11] ),
    .CLK(clknet_leaf_129_clk_regs));
 sg13g2_dfrbpq_1 _09226_ (.RESET_B(net664),
    .D(_00632_),
    .Q(\rf_ram.RAM[3][12] ),
    .CLK(clknet_leaf_128_clk_regs));
 sg13g2_dfrbpq_1 _09227_ (.RESET_B(net663),
    .D(_00633_),
    .Q(\rf_ram.RAM[3][13] ),
    .CLK(clknet_leaf_110_clk_regs));
 sg13g2_dfrbpq_1 _09228_ (.RESET_B(net662),
    .D(_00634_),
    .Q(\rf_ram.RAM[3][14] ),
    .CLK(clknet_leaf_161_clk_regs));
 sg13g2_dfrbpq_1 _09229_ (.RESET_B(net661),
    .D(_00635_),
    .Q(\rf_ram.RAM[3][15] ),
    .CLK(clknet_leaf_148_clk_regs));
 sg13g2_dfrbpq_1 _09230_ (.RESET_B(net660),
    .D(_00636_),
    .Q(\rf_ram.RAM[3][16] ),
    .CLK(clknet_leaf_102_clk_regs));
 sg13g2_dfrbpq_1 _09231_ (.RESET_B(net659),
    .D(_00637_),
    .Q(\rf_ram.RAM[3][17] ),
    .CLK(clknet_leaf_139_clk_regs));
 sg13g2_dfrbpq_1 _09232_ (.RESET_B(net658),
    .D(_00638_),
    .Q(\rf_ram.RAM[3][18] ),
    .CLK(clknet_leaf_137_clk_regs));
 sg13g2_dfrbpq_1 _09233_ (.RESET_B(net657),
    .D(_00639_),
    .Q(\rf_ram.RAM[3][19] ),
    .CLK(clknet_leaf_152_clk_regs));
 sg13g2_dfrbpq_1 _09234_ (.RESET_B(net656),
    .D(_00640_),
    .Q(\rf_ram.RAM[3][20] ),
    .CLK(clknet_leaf_153_clk_regs));
 sg13g2_dfrbpq_1 _09235_ (.RESET_B(net655),
    .D(_00641_),
    .Q(\rf_ram.RAM[3][21] ),
    .CLK(clknet_leaf_22_clk_regs));
 sg13g2_dfrbpq_1 _09236_ (.RESET_B(net654),
    .D(_00642_),
    .Q(\rf_ram.RAM[3][22] ),
    .CLK(clknet_leaf_64_clk_regs));
 sg13g2_dfrbpq_1 _09237_ (.RESET_B(net653),
    .D(_00643_),
    .Q(\rf_ram.RAM[3][23] ),
    .CLK(clknet_leaf_20_clk_regs));
 sg13g2_dfrbpq_1 _09238_ (.RESET_B(net652),
    .D(_00644_),
    .Q(\rf_ram.RAM[3][24] ),
    .CLK(clknet_leaf_74_clk_regs));
 sg13g2_dfrbpq_1 _09239_ (.RESET_B(net651),
    .D(_00645_),
    .Q(\rf_ram.RAM[3][25] ),
    .CLK(clknet_leaf_46_clk_regs));
 sg13g2_dfrbpq_1 _09240_ (.RESET_B(net650),
    .D(_00646_),
    .Q(\rf_ram.RAM[3][26] ),
    .CLK(clknet_leaf_50_clk_regs));
 sg13g2_dfrbpq_1 _09241_ (.RESET_B(net649),
    .D(_00647_),
    .Q(\rf_ram.RAM[3][27] ),
    .CLK(clknet_leaf_45_clk_regs));
 sg13g2_dfrbpq_1 _09242_ (.RESET_B(net648),
    .D(_00648_),
    .Q(\rf_ram.RAM[3][28] ),
    .CLK(clknet_leaf_27_clk_regs));
 sg13g2_dfrbpq_1 _09243_ (.RESET_B(net647),
    .D(_00649_),
    .Q(\rf_ram.RAM[3][29] ),
    .CLK(clknet_leaf_167_clk_regs));
 sg13g2_dfrbpq_1 _09244_ (.RESET_B(net646),
    .D(_00650_),
    .Q(\rf_ram.RAM[3][30] ),
    .CLK(clknet_leaf_165_clk_regs));
 sg13g2_dfrbpq_1 _09245_ (.RESET_B(net645),
    .D(_00651_),
    .Q(\rf_ram.RAM[3][31] ),
    .CLK(clknet_leaf_167_clk_regs));
 sg13g2_dfrbpq_1 _09246_ (.RESET_B(net644),
    .D(net1447),
    .Q(\rf_ram.RAM[4][0] ),
    .CLK(clknet_leaf_153_clk_regs));
 sg13g2_dfrbpq_1 _09247_ (.RESET_B(net643),
    .D(_00653_),
    .Q(\rf_ram.RAM[4][1] ),
    .CLK(clknet_leaf_55_clk_regs));
 sg13g2_dfrbpq_1 _09248_ (.RESET_B(net642),
    .D(_00654_),
    .Q(\rf_ram.RAM[4][2] ),
    .CLK(clknet_leaf_70_clk_regs));
 sg13g2_dfrbpq_1 _09249_ (.RESET_B(net641),
    .D(_00655_),
    .Q(\rf_ram.RAM[4][3] ),
    .CLK(clknet_leaf_89_clk_regs));
 sg13g2_dfrbpq_1 _09250_ (.RESET_B(net640),
    .D(_00656_),
    .Q(\rf_ram.RAM[4][4] ),
    .CLK(clknet_leaf_88_clk_regs));
 sg13g2_dfrbpq_1 _09251_ (.RESET_B(net639),
    .D(_00657_),
    .Q(\rf_ram.RAM[4][5] ),
    .CLK(clknet_leaf_88_clk_regs));
 sg13g2_dfrbpq_1 _09252_ (.RESET_B(net638),
    .D(_00658_),
    .Q(\rf_ram.RAM[4][6] ),
    .CLK(clknet_leaf_95_clk_regs));
 sg13g2_dfrbpq_1 _09253_ (.RESET_B(net637),
    .D(_00659_),
    .Q(\rf_ram.RAM[4][7] ),
    .CLK(clknet_leaf_99_clk_regs));
 sg13g2_dfrbpq_1 _09254_ (.RESET_B(net636),
    .D(_00660_),
    .Q(\rf_ram.RAM[4][8] ),
    .CLK(clknet_leaf_117_clk_regs));
 sg13g2_dfrbpq_1 _09255_ (.RESET_B(net635),
    .D(_00661_),
    .Q(\rf_ram.RAM[4][9] ),
    .CLK(clknet_leaf_126_clk_regs));
 sg13g2_dfrbpq_1 _09256_ (.RESET_B(net634),
    .D(_00662_),
    .Q(\rf_ram.RAM[4][10] ),
    .CLK(clknet_leaf_125_clk_regs));
 sg13g2_dfrbpq_1 _09257_ (.RESET_B(net633),
    .D(_00663_),
    .Q(\rf_ram.RAM[4][11] ),
    .CLK(clknet_leaf_133_clk_regs));
 sg13g2_dfrbpq_1 _09258_ (.RESET_B(net632),
    .D(_00664_),
    .Q(\rf_ram.RAM[4][12] ),
    .CLK(clknet_leaf_127_clk_regs));
 sg13g2_dfrbpq_1 _09259_ (.RESET_B(net631),
    .D(_00665_),
    .Q(\rf_ram.RAM[4][13] ),
    .CLK(clknet_leaf_143_clk_regs));
 sg13g2_dfrbpq_1 _09260_ (.RESET_B(net630),
    .D(_00666_),
    .Q(\rf_ram.RAM[4][14] ),
    .CLK(clknet_leaf_156_clk_regs));
 sg13g2_dfrbpq_1 _09261_ (.RESET_B(net629),
    .D(_00667_),
    .Q(\rf_ram.RAM[4][15] ),
    .CLK(clknet_leaf_145_clk_regs));
 sg13g2_dfrbpq_1 _09262_ (.RESET_B(net628),
    .D(_00668_),
    .Q(\rf_ram.RAM[4][16] ),
    .CLK(clknet_leaf_64_clk_regs));
 sg13g2_dfrbpq_1 _09263_ (.RESET_B(net627),
    .D(_00669_),
    .Q(\rf_ram.RAM[4][17] ),
    .CLK(clknet_leaf_138_clk_regs));
 sg13g2_dfrbpq_1 _09264_ (.RESET_B(net626),
    .D(_00670_),
    .Q(\rf_ram.RAM[4][18] ),
    .CLK(clknet_leaf_133_clk_regs));
 sg13g2_dfrbpq_1 _09265_ (.RESET_B(net625),
    .D(_00671_),
    .Q(\rf_ram.RAM[4][19] ),
    .CLK(clknet_leaf_162_clk_regs));
 sg13g2_dfrbpq_1 _09266_ (.RESET_B(net624),
    .D(_00672_),
    .Q(\rf_ram.RAM[4][20] ),
    .CLK(clknet_leaf_151_clk_regs));
 sg13g2_dfrbpq_1 _09267_ (.RESET_B(net623),
    .D(_00673_),
    .Q(\rf_ram.RAM[4][21] ),
    .CLK(clknet_leaf_63_clk_regs));
 sg13g2_dfrbpq_1 _09268_ (.RESET_B(net622),
    .D(_00674_),
    .Q(\rf_ram.RAM[4][22] ),
    .CLK(clknet_leaf_66_clk_regs));
 sg13g2_dfrbpq_1 _09269_ (.RESET_B(net621),
    .D(_00675_),
    .Q(\rf_ram.RAM[4][23] ),
    .CLK(clknet_leaf_21_clk_regs));
 sg13g2_dfrbpq_1 _09270_ (.RESET_B(net620),
    .D(_00676_),
    .Q(\rf_ram.RAM[4][24] ),
    .CLK(clknet_leaf_72_clk_regs));
 sg13g2_dfrbpq_1 _09271_ (.RESET_B(net619),
    .D(_00677_),
    .Q(\rf_ram.RAM[4][25] ),
    .CLK(clknet_leaf_57_clk_regs));
 sg13g2_dfrbpq_1 _09272_ (.RESET_B(net618),
    .D(_00678_),
    .Q(\rf_ram.RAM[4][26] ),
    .CLK(clknet_leaf_56_clk_regs));
 sg13g2_dfrbpq_1 _09273_ (.RESET_B(net617),
    .D(_00679_),
    .Q(\rf_ram.RAM[4][27] ),
    .CLK(clknet_leaf_46_clk_regs));
 sg13g2_dfrbpq_1 _09274_ (.RESET_B(net616),
    .D(_00680_),
    .Q(\rf_ram.RAM[4][28] ),
    .CLK(clknet_leaf_24_clk_regs));
 sg13g2_dfrbpq_1 _09275_ (.RESET_B(net615),
    .D(_00681_),
    .Q(\rf_ram.RAM[4][29] ),
    .CLK(clknet_leaf_167_clk_regs));
 sg13g2_dfrbpq_1 _09276_ (.RESET_B(net614),
    .D(_00682_),
    .Q(\rf_ram.RAM[4][30] ),
    .CLK(clknet_leaf_162_clk_regs));
 sg13g2_dfrbpq_1 _09277_ (.RESET_B(net83),
    .D(_00683_),
    .Q(\rf_ram.RAM[4][31] ),
    .CLK(clknet_leaf_169_clk_regs));
 sg13g2_dfrbpq_2 _09278_ (.RESET_B(net2599),
    .D(_00065_),
    .Q(\ram_spi_if.cycle_counter[0] ),
    .CLK(clknet_leaf_37_clk_regs));
 sg13g2_dfrbpq_2 _09279_ (.RESET_B(net2599),
    .D(_00066_),
    .Q(\ram_spi_if.cycle_counter[1] ),
    .CLK(clknet_leaf_38_clk_regs));
 sg13g2_dfrbpq_1 _09280_ (.RESET_B(net2599),
    .D(net3343),
    .Q(\ram_spi_if.cycle_counter[2] ),
    .CLK(clknet_leaf_37_clk_regs));
 sg13g2_dfrbpq_2 _09281_ (.RESET_B(net2599),
    .D(net3497),
    .Q(\ram_spi_if.cycle_counter[3] ),
    .CLK(clknet_leaf_37_clk_regs));
 sg13g2_dfrbpq_1 _09282_ (.RESET_B(net2599),
    .D(net3463),
    .Q(\ram_spi_if.cycle_counter[4] ),
    .CLK(clknet_leaf_37_clk_regs));
 sg13g2_dfrbpq_2 _09283_ (.RESET_B(net2599),
    .D(_00070_),
    .Q(\ram_spi_if.cycle_counter[5] ),
    .CLK(clknet_leaf_36_clk_regs));
 sg13g2_dfrbpq_1 _09284_ (.RESET_B(net2600),
    .D(_00684_),
    .Q(\ram_spi_if.state_reg[0] ),
    .CLK(clknet_leaf_36_clk_regs));
 sg13g2_dfrbpq_2 _09285_ (.RESET_B(net2600),
    .D(_00685_),
    .Q(\ram_spi_if.state_reg[1] ),
    .CLK(clknet_leaf_36_clk_regs));
 sg13g2_dfrbpq_2 _09286_ (.RESET_B(net2600),
    .D(net3706),
    .Q(\ram_spi_if.state_reg[2] ),
    .CLK(clknet_leaf_36_clk_regs));
 sg13g2_dfrbpq_1 _09287_ (.RESET_B(net2600),
    .D(net3727),
    .Q(\ram_spi_if.state_reg[3] ),
    .CLK(clknet_leaf_36_clk_regs));
 sg13g2_dfrbpq_1 _09288_ (.RESET_B(net613),
    .D(net3157),
    .Q(\rf_ram.RAM[15][0] ),
    .CLK(clknet_leaf_17_clk_regs));
 sg13g2_dfrbpq_1 _09289_ (.RESET_B(net612),
    .D(_00689_),
    .Q(\rf_ram.RAM[15][1] ),
    .CLK(clknet_leaf_53_clk_regs));
 sg13g2_dfrbpq_1 _09290_ (.RESET_B(net611),
    .D(_00690_),
    .Q(\rf_ram.RAM[15][2] ),
    .CLK(clknet_leaf_77_clk_regs));
 sg13g2_dfrbpq_1 _09291_ (.RESET_B(net610),
    .D(_00691_),
    .Q(\rf_ram.RAM[15][3] ),
    .CLK(clknet_leaf_84_clk_regs));
 sg13g2_dfrbpq_1 _09292_ (.RESET_B(net609),
    .D(_00692_),
    .Q(\rf_ram.RAM[15][4] ),
    .CLK(clknet_leaf_77_clk_regs));
 sg13g2_dfrbpq_1 _09293_ (.RESET_B(net608),
    .D(_00693_),
    .Q(\rf_ram.RAM[15][5] ),
    .CLK(clknet_leaf_84_clk_regs));
 sg13g2_dfrbpq_1 _09294_ (.RESET_B(net607),
    .D(_00694_),
    .Q(\rf_ram.RAM[15][6] ),
    .CLK(clknet_leaf_94_clk_regs));
 sg13g2_dfrbpq_1 _09295_ (.RESET_B(net606),
    .D(_00695_),
    .Q(\rf_ram.RAM[15][7] ),
    .CLK(clknet_leaf_94_clk_regs));
 sg13g2_dfrbpq_1 _09296_ (.RESET_B(net605),
    .D(_00696_),
    .Q(\rf_ram.RAM[15][8] ),
    .CLK(clknet_leaf_115_clk_regs));
 sg13g2_dfrbpq_1 _09297_ (.RESET_B(net604),
    .D(_00697_),
    .Q(\rf_ram.RAM[15][9] ),
    .CLK(clknet_leaf_124_clk_regs));
 sg13g2_dfrbpq_1 _09298_ (.RESET_B(net603),
    .D(_00698_),
    .Q(\rf_ram.RAM[15][10] ),
    .CLK(clknet_leaf_120_clk_regs));
 sg13g2_dfrbpq_1 _09299_ (.RESET_B(net602),
    .D(_00699_),
    .Q(\rf_ram.RAM[15][11] ),
    .CLK(clknet_leaf_132_clk_regs));
 sg13g2_dfrbpq_1 _09300_ (.RESET_B(net601),
    .D(_00700_),
    .Q(\rf_ram.RAM[15][12] ),
    .CLK(clknet_leaf_118_clk_regs));
 sg13g2_dfrbpq_1 _09301_ (.RESET_B(net600),
    .D(_00701_),
    .Q(\rf_ram.RAM[15][13] ),
    .CLK(clknet_leaf_103_clk_regs));
 sg13g2_dfrbpq_1 _09302_ (.RESET_B(net599),
    .D(_00702_),
    .Q(\rf_ram.RAM[15][14] ),
    .CLK(clknet_leaf_157_clk_regs));
 sg13g2_dfrbpq_1 _09303_ (.RESET_B(net598),
    .D(_00703_),
    .Q(\rf_ram.RAM[15][15] ),
    .CLK(clknet_leaf_147_clk_regs));
 sg13g2_dfrbpq_1 _09304_ (.RESET_B(net597),
    .D(_00704_),
    .Q(\rf_ram.RAM[15][16] ),
    .CLK(clknet_leaf_108_clk_regs));
 sg13g2_dfrbpq_1 _09305_ (.RESET_B(net596),
    .D(_00705_),
    .Q(\rf_ram.RAM[15][17] ),
    .CLK(clknet_leaf_141_clk_regs));
 sg13g2_dfrbpq_1 _09306_ (.RESET_B(net595),
    .D(_00706_),
    .Q(\rf_ram.RAM[15][18] ),
    .CLK(clknet_leaf_132_clk_regs));
 sg13g2_dfrbpq_1 _09307_ (.RESET_B(net594),
    .D(_00707_),
    .Q(\rf_ram.RAM[15][19] ),
    .CLK(clknet_leaf_155_clk_regs));
 sg13g2_dfrbpq_1 _09308_ (.RESET_B(net593),
    .D(_00708_),
    .Q(\rf_ram.RAM[15][20] ),
    .CLK(clknet_leaf_151_clk_regs));
 sg13g2_dfrbpq_1 _09309_ (.RESET_B(net592),
    .D(_00709_),
    .Q(\rf_ram.RAM[15][21] ),
    .CLK(clknet_leaf_60_clk_regs));
 sg13g2_dfrbpq_1 _09310_ (.RESET_B(net591),
    .D(_00710_),
    .Q(\rf_ram.RAM[15][22] ),
    .CLK(clknet_leaf_102_clk_regs));
 sg13g2_dfrbpq_1 _09311_ (.RESET_B(net590),
    .D(_00711_),
    .Q(\rf_ram.RAM[15][23] ),
    .CLK(clknet_leaf_25_clk_regs));
 sg13g2_dfrbpq_1 _09312_ (.RESET_B(net589),
    .D(_00712_),
    .Q(\rf_ram.RAM[15][24] ),
    .CLK(clknet_leaf_75_clk_regs));
 sg13g2_dfrbpq_1 _09313_ (.RESET_B(net588),
    .D(_00713_),
    .Q(\rf_ram.RAM[15][25] ),
    .CLK(clknet_leaf_53_clk_regs));
 sg13g2_dfrbpq_1 _09314_ (.RESET_B(net587),
    .D(_00714_),
    .Q(\rf_ram.RAM[15][26] ),
    .CLK(clknet_leaf_47_clk_regs));
 sg13g2_dfrbpq_1 _09315_ (.RESET_B(net586),
    .D(_00715_),
    .Q(\rf_ram.RAM[15][27] ),
    .CLK(clknet_leaf_44_clk_regs));
 sg13g2_dfrbpq_1 _09316_ (.RESET_B(net585),
    .D(_00716_),
    .Q(\rf_ram.RAM[15][28] ),
    .CLK(clknet_leaf_25_clk_regs));
 sg13g2_dfrbpq_1 _09317_ (.RESET_B(net584),
    .D(_00717_),
    .Q(\rf_ram.RAM[15][29] ),
    .CLK(clknet_leaf_5_clk_regs));
 sg13g2_dfrbpq_1 _09318_ (.RESET_B(net583),
    .D(_00718_),
    .Q(\rf_ram.RAM[15][30] ),
    .CLK(clknet_leaf_165_clk_regs));
 sg13g2_dfrbpq_1 _09319_ (.RESET_B(net582),
    .D(_00719_),
    .Q(\rf_ram.RAM[15][31] ),
    .CLK(clknet_leaf_166_clk_regs));
 sg13g2_dfrbpq_1 _09320_ (.RESET_B(net581),
    .D(net2919),
    .Q(\rf_ram.RAM[9][0] ),
    .CLK(clknet_leaf_16_clk_regs));
 sg13g2_dfrbpq_1 _09321_ (.RESET_B(net580),
    .D(_00721_),
    .Q(\rf_ram.RAM[9][1] ),
    .CLK(clknet_leaf_54_clk_regs));
 sg13g2_dfrbpq_1 _09322_ (.RESET_B(net579),
    .D(_00722_),
    .Q(\rf_ram.RAM[9][2] ),
    .CLK(clknet_leaf_75_clk_regs));
 sg13g2_dfrbpq_1 _09323_ (.RESET_B(net578),
    .D(_00723_),
    .Q(\rf_ram.RAM[9][3] ),
    .CLK(clknet_leaf_79_clk_regs));
 sg13g2_dfrbpq_1 _09324_ (.RESET_B(net577),
    .D(_00724_),
    .Q(\rf_ram.RAM[9][4] ),
    .CLK(clknet_leaf_82_clk_regs));
 sg13g2_dfrbpq_1 _09325_ (.RESET_B(net576),
    .D(_00725_),
    .Q(\rf_ram.RAM[9][5] ),
    .CLK(clknet_leaf_80_clk_regs));
 sg13g2_dfrbpq_1 _09326_ (.RESET_B(net575),
    .D(_00726_),
    .Q(\rf_ram.RAM[9][6] ),
    .CLK(clknet_leaf_100_clk_regs));
 sg13g2_dfrbpq_1 _09327_ (.RESET_B(net574),
    .D(_00727_),
    .Q(\rf_ram.RAM[9][7] ),
    .CLK(clknet_leaf_98_clk_regs));
 sg13g2_dfrbpq_1 _09328_ (.RESET_B(net573),
    .D(_00728_),
    .Q(\rf_ram.RAM[9][8] ),
    .CLK(clknet_leaf_113_clk_regs));
 sg13g2_dfrbpq_1 _09329_ (.RESET_B(net572),
    .D(_00729_),
    .Q(\rf_ram.RAM[9][9] ),
    .CLK(clknet_leaf_131_clk_regs));
 sg13g2_dfrbpq_1 _09330_ (.RESET_B(net571),
    .D(_00730_),
    .Q(\rf_ram.RAM[9][10] ),
    .CLK(clknet_leaf_111_clk_regs));
 sg13g2_dfrbpq_1 _09331_ (.RESET_B(net570),
    .D(_00731_),
    .Q(\rf_ram.RAM[9][11] ),
    .CLK(clknet_leaf_129_clk_regs));
 sg13g2_dfrbpq_1 _09332_ (.RESET_B(net569),
    .D(_00732_),
    .Q(\rf_ram.RAM[9][12] ),
    .CLK(clknet_leaf_130_clk_regs));
 sg13g2_dfrbpq_1 _09333_ (.RESET_B(net568),
    .D(_00733_),
    .Q(\rf_ram.RAM[9][13] ),
    .CLK(clknet_leaf_98_clk_regs));
 sg13g2_dfrbpq_1 _09334_ (.RESET_B(net567),
    .D(_00734_),
    .Q(\rf_ram.RAM[9][14] ),
    .CLK(clknet_leaf_161_clk_regs));
 sg13g2_dfrbpq_1 _09335_ (.RESET_B(net566),
    .D(_00735_),
    .Q(\rf_ram.RAM[9][15] ),
    .CLK(clknet_leaf_109_clk_regs));
 sg13g2_dfrbpq_1 _09336_ (.RESET_B(net565),
    .D(_00736_),
    .Q(\rf_ram.RAM[9][16] ),
    .CLK(clknet_leaf_68_clk_regs));
 sg13g2_dfrbpq_1 _09337_ (.RESET_B(net564),
    .D(_00737_),
    .Q(\rf_ram.RAM[9][17] ),
    .CLK(clknet_leaf_138_clk_regs));
 sg13g2_dfrbpq_1 _09338_ (.RESET_B(net563),
    .D(_00738_),
    .Q(\rf_ram.RAM[9][18] ),
    .CLK(clknet_leaf_136_clk_regs));
 sg13g2_dfrbpq_1 _09339_ (.RESET_B(net562),
    .D(_00739_),
    .Q(\rf_ram.RAM[9][19] ),
    .CLK(clknet_leaf_161_clk_regs));
 sg13g2_dfrbpq_1 _09340_ (.RESET_B(net561),
    .D(_00740_),
    .Q(\rf_ram.RAM[9][20] ),
    .CLK(clknet_leaf_152_clk_regs));
 sg13g2_dfrbpq_1 _09341_ (.RESET_B(net560),
    .D(_00741_),
    .Q(\rf_ram.RAM[9][21] ),
    .CLK(clknet_leaf_61_clk_regs));
 sg13g2_dfrbpq_1 _09342_ (.RESET_B(net559),
    .D(_00742_),
    .Q(\rf_ram.RAM[9][22] ),
    .CLK(clknet_leaf_105_clk_regs));
 sg13g2_dfrbpq_1 _09343_ (.RESET_B(net558),
    .D(_00743_),
    .Q(\rf_ram.RAM[9][23] ),
    .CLK(clknet_leaf_20_clk_regs));
 sg13g2_dfrbpq_1 _09344_ (.RESET_B(net557),
    .D(_00744_),
    .Q(\rf_ram.RAM[9][24] ),
    .CLK(clknet_leaf_72_clk_regs));
 sg13g2_dfrbpq_1 _09345_ (.RESET_B(net556),
    .D(_00745_),
    .Q(\rf_ram.RAM[9][25] ),
    .CLK(clknet_leaf_57_clk_regs));
 sg13g2_dfrbpq_1 _09346_ (.RESET_B(net555),
    .D(_00746_),
    .Q(\rf_ram.RAM[9][26] ),
    .CLK(clknet_leaf_58_clk_regs));
 sg13g2_dfrbpq_1 _09347_ (.RESET_B(net554),
    .D(_00747_),
    .Q(\rf_ram.RAM[9][27] ),
    .CLK(clknet_leaf_35_clk_regs));
 sg13g2_dfrbpq_1 _09348_ (.RESET_B(net553),
    .D(_00748_),
    .Q(\rf_ram.RAM[9][28] ),
    .CLK(clknet_leaf_28_clk_regs));
 sg13g2_dfrbpq_1 _09349_ (.RESET_B(net552),
    .D(_00749_),
    .Q(\rf_ram.RAM[9][29] ),
    .CLK(clknet_leaf_5_clk_regs));
 sg13g2_dfrbpq_1 _09350_ (.RESET_B(net551),
    .D(_00750_),
    .Q(\rf_ram.RAM[9][30] ),
    .CLK(clknet_leaf_164_clk_regs));
 sg13g2_dfrbpq_1 _09351_ (.RESET_B(net550),
    .D(_00751_),
    .Q(\rf_ram.RAM[9][31] ),
    .CLK(clknet_leaf_167_clk_regs));
 sg13g2_dfrbpq_1 _09352_ (.RESET_B(net549),
    .D(net2899),
    .Q(\rf_ram.RAM[14][0] ),
    .CLK(clknet_leaf_20_clk_regs));
 sg13g2_dfrbpq_1 _09353_ (.RESET_B(net548),
    .D(_00753_),
    .Q(\rf_ram.RAM[14][1] ),
    .CLK(clknet_leaf_53_clk_regs));
 sg13g2_dfrbpq_1 _09354_ (.RESET_B(net547),
    .D(_00754_),
    .Q(\rf_ram.RAM[14][2] ),
    .CLK(clknet_leaf_77_clk_regs));
 sg13g2_dfrbpq_1 _09355_ (.RESET_B(net546),
    .D(_00755_),
    .Q(\rf_ram.RAM[14][3] ),
    .CLK(clknet_leaf_83_clk_regs));
 sg13g2_dfrbpq_1 _09356_ (.RESET_B(net545),
    .D(_00756_),
    .Q(\rf_ram.RAM[14][4] ),
    .CLK(clknet_leaf_82_clk_regs));
 sg13g2_dfrbpq_1 _09357_ (.RESET_B(net544),
    .D(_00757_),
    .Q(\rf_ram.RAM[14][5] ),
    .CLK(clknet_leaf_85_clk_regs));
 sg13g2_dfrbpq_1 _09358_ (.RESET_B(net543),
    .D(_00758_),
    .Q(\rf_ram.RAM[14][6] ),
    .CLK(clknet_leaf_91_clk_regs));
 sg13g2_dfrbpq_1 _09359_ (.RESET_B(net542),
    .D(_00759_),
    .Q(\rf_ram.RAM[14][7] ),
    .CLK(clknet_leaf_92_clk_regs));
 sg13g2_dfrbpq_1 _09360_ (.RESET_B(net541),
    .D(_00760_),
    .Q(\rf_ram.RAM[14][8] ),
    .CLK(clknet_leaf_114_clk_regs));
 sg13g2_dfrbpq_1 _09361_ (.RESET_B(net540),
    .D(_00761_),
    .Q(\rf_ram.RAM[14][9] ),
    .CLK(clknet_leaf_124_clk_regs));
 sg13g2_dfrbpq_1 _09362_ (.RESET_B(net539),
    .D(_00762_),
    .Q(\rf_ram.RAM[14][10] ),
    .CLK(clknet_leaf_120_clk_regs));
 sg13g2_dfrbpq_1 _09363_ (.RESET_B(net538),
    .D(_00763_),
    .Q(\rf_ram.RAM[14][11] ),
    .CLK(clknet_leaf_131_clk_regs));
 sg13g2_dfrbpq_1 _09364_ (.RESET_B(net537),
    .D(_00764_),
    .Q(\rf_ram.RAM[14][12] ),
    .CLK(clknet_leaf_118_clk_regs));
 sg13g2_dfrbpq_1 _09365_ (.RESET_B(net536),
    .D(_00765_),
    .Q(\rf_ram.RAM[14][13] ),
    .CLK(clknet_leaf_103_clk_regs));
 sg13g2_dfrbpq_1 _09366_ (.RESET_B(net535),
    .D(_00766_),
    .Q(\rf_ram.RAM[14][14] ),
    .CLK(clknet_leaf_157_clk_regs));
 sg13g2_dfrbpq_1 _09367_ (.RESET_B(net534),
    .D(_00767_),
    .Q(\rf_ram.RAM[14][15] ),
    .CLK(clknet_leaf_148_clk_regs));
 sg13g2_dfrbpq_1 _09368_ (.RESET_B(net533),
    .D(_00768_),
    .Q(\rf_ram.RAM[14][16] ),
    .CLK(clknet_leaf_108_clk_regs));
 sg13g2_dfrbpq_1 _09369_ (.RESET_B(net532),
    .D(_00769_),
    .Q(\rf_ram.RAM[14][17] ),
    .CLK(clknet_leaf_140_clk_regs));
 sg13g2_dfrbpq_1 _09370_ (.RESET_B(net531),
    .D(_00770_),
    .Q(\rf_ram.RAM[14][18] ),
    .CLK(clknet_leaf_132_clk_regs));
 sg13g2_dfrbpq_1 _09371_ (.RESET_B(net530),
    .D(_00771_),
    .Q(\rf_ram.RAM[14][19] ),
    .CLK(clknet_leaf_155_clk_regs));
 sg13g2_dfrbpq_1 _09372_ (.RESET_B(net529),
    .D(_00772_),
    .Q(\rf_ram.RAM[14][20] ),
    .CLK(clknet_leaf_150_clk_regs));
 sg13g2_dfrbpq_1 _09373_ (.RESET_B(net528),
    .D(_00773_),
    .Q(\rf_ram.RAM[14][21] ),
    .CLK(clknet_leaf_60_clk_regs));
 sg13g2_dfrbpq_1 _09374_ (.RESET_B(net527),
    .D(_00774_),
    .Q(\rf_ram.RAM[14][22] ),
    .CLK(clknet_leaf_67_clk_regs));
 sg13g2_dfrbpq_1 _09375_ (.RESET_B(net526),
    .D(_00775_),
    .Q(\rf_ram.RAM[14][23] ),
    .CLK(clknet_leaf_19_clk_regs));
 sg13g2_dfrbpq_1 _09376_ (.RESET_B(net525),
    .D(_00776_),
    .Q(\rf_ram.RAM[14][24] ),
    .CLK(clknet_leaf_74_clk_regs));
 sg13g2_dfrbpq_1 _09377_ (.RESET_B(net524),
    .D(_00777_),
    .Q(\rf_ram.RAM[14][25] ),
    .CLK(clknet_leaf_53_clk_regs));
 sg13g2_dfrbpq_1 _09378_ (.RESET_B(net523),
    .D(_00778_),
    .Q(\rf_ram.RAM[14][26] ),
    .CLK(clknet_leaf_50_clk_regs));
 sg13g2_dfrbpq_1 _09379_ (.RESET_B(net522),
    .D(_00779_),
    .Q(\rf_ram.RAM[14][27] ),
    .CLK(clknet_leaf_48_clk_regs));
 sg13g2_dfrbpq_1 _09380_ (.RESET_B(net521),
    .D(_00780_),
    .Q(\rf_ram.RAM[14][28] ),
    .CLK(clknet_leaf_26_clk_regs));
 sg13g2_dfrbpq_1 _09381_ (.RESET_B(net520),
    .D(_00781_),
    .Q(\rf_ram.RAM[14][29] ),
    .CLK(clknet_leaf_5_clk_regs));
 sg13g2_dfrbpq_1 _09382_ (.RESET_B(net519),
    .D(_00782_),
    .Q(\rf_ram.RAM[14][30] ),
    .CLK(clknet_leaf_164_clk_regs));
 sg13g2_dfrbpq_1 _09383_ (.RESET_B(net518),
    .D(_00783_),
    .Q(\rf_ram.RAM[14][31] ),
    .CLK(clknet_leaf_166_clk_regs));
 sg13g2_dfrbpq_1 _09384_ (.RESET_B(net517),
    .D(_00784_),
    .Q(uo_out[4]),
    .CLK(clknet_leaf_40_clk_regs));
 sg13g2_dfrbpq_1 _09385_ (.RESET_B(net515),
    .D(_00785_),
    .Q(uo_out[5]),
    .CLK(clknet_leaf_41_clk_regs));
 sg13g2_dfrbpq_1 _09386_ (.RESET_B(net513),
    .D(_00786_),
    .Q(uo_out[6]),
    .CLK(clknet_leaf_42_clk_regs));
 sg13g2_dfrbpq_1 _09387_ (.RESET_B(net511),
    .D(_00787_),
    .Q(uo_out[7]),
    .CLK(clknet_leaf_42_clk_regs));
 sg13g2_dfrbpq_1 _09388_ (.RESET_B(net509),
    .D(net2914),
    .Q(\rf_ram.RAM[7][0] ),
    .CLK(clknet_leaf_153_clk_regs));
 sg13g2_dfrbpq_1 _09389_ (.RESET_B(net508),
    .D(_00789_),
    .Q(\rf_ram.RAM[7][1] ),
    .CLK(clknet_leaf_54_clk_regs));
 sg13g2_dfrbpq_1 _09390_ (.RESET_B(net507),
    .D(_00790_),
    .Q(\rf_ram.RAM[7][2] ),
    .CLK(clknet_leaf_69_clk_regs));
 sg13g2_dfrbpq_1 _09391_ (.RESET_B(net506),
    .D(_00791_),
    .Q(\rf_ram.RAM[7][3] ),
    .CLK(clknet_leaf_89_clk_regs));
 sg13g2_dfrbpq_1 _09392_ (.RESET_B(net505),
    .D(_00792_),
    .Q(\rf_ram.RAM[7][4] ),
    .CLK(clknet_leaf_88_clk_regs));
 sg13g2_dfrbpq_1 _09393_ (.RESET_B(net504),
    .D(_00793_),
    .Q(\rf_ram.RAM[7][5] ),
    .CLK(clknet_leaf_88_clk_regs));
 sg13g2_dfrbpq_1 _09394_ (.RESET_B(net503),
    .D(_00794_),
    .Q(\rf_ram.RAM[7][6] ),
    .CLK(clknet_leaf_96_clk_regs));
 sg13g2_dfrbpq_1 _09395_ (.RESET_B(net502),
    .D(_00795_),
    .Q(\rf_ram.RAM[7][7] ),
    .CLK(clknet_leaf_91_clk_regs));
 sg13g2_dfrbpq_1 _09396_ (.RESET_B(net501),
    .D(_00796_),
    .Q(\rf_ram.RAM[7][8] ),
    .CLK(clknet_leaf_117_clk_regs));
 sg13g2_dfrbpq_1 _09397_ (.RESET_B(net500),
    .D(_00797_),
    .Q(\rf_ram.RAM[7][9] ),
    .CLK(clknet_leaf_126_clk_regs));
 sg13g2_dfrbpq_1 _09398_ (.RESET_B(net499),
    .D(_00798_),
    .Q(\rf_ram.RAM[7][10] ),
    .CLK(clknet_leaf_125_clk_regs));
 sg13g2_dfrbpq_1 _09399_ (.RESET_B(net498),
    .D(_00799_),
    .Q(\rf_ram.RAM[7][11] ),
    .CLK(clknet_leaf_133_clk_regs));
 sg13g2_dfrbpq_1 _09400_ (.RESET_B(net497),
    .D(_00800_),
    .Q(\rf_ram.RAM[7][12] ),
    .CLK(clknet_leaf_127_clk_regs));
 sg13g2_dfrbpq_1 _09401_ (.RESET_B(net496),
    .D(_00801_),
    .Q(\rf_ram.RAM[7][13] ),
    .CLK(clknet_leaf_143_clk_regs));
 sg13g2_dfrbpq_1 _09402_ (.RESET_B(net495),
    .D(_00802_),
    .Q(\rf_ram.RAM[7][14] ),
    .CLK(clknet_leaf_157_clk_regs));
 sg13g2_dfrbpq_1 _09403_ (.RESET_B(net494),
    .D(_00803_),
    .Q(\rf_ram.RAM[7][15] ),
    .CLK(clknet_leaf_145_clk_regs));
 sg13g2_dfrbpq_1 _09404_ (.RESET_B(net493),
    .D(_00804_),
    .Q(\rf_ram.RAM[7][16] ),
    .CLK(clknet_leaf_105_clk_regs));
 sg13g2_dfrbpq_1 _09405_ (.RESET_B(net492),
    .D(_00805_),
    .Q(\rf_ram.RAM[7][17] ),
    .CLK(clknet_leaf_159_clk_regs));
 sg13g2_dfrbpq_1 _09406_ (.RESET_B(net491),
    .D(_00806_),
    .Q(\rf_ram.RAM[7][18] ),
    .CLK(clknet_leaf_133_clk_regs));
 sg13g2_dfrbpq_1 _09407_ (.RESET_B(net490),
    .D(_00807_),
    .Q(\rf_ram.RAM[7][19] ),
    .CLK(clknet_leaf_162_clk_regs));
 sg13g2_dfrbpq_1 _09408_ (.RESET_B(net489),
    .D(_00808_),
    .Q(\rf_ram.RAM[7][20] ),
    .CLK(clknet_leaf_151_clk_regs));
 sg13g2_dfrbpq_1 _09409_ (.RESET_B(net488),
    .D(_00809_),
    .Q(\rf_ram.RAM[7][21] ),
    .CLK(clknet_leaf_62_clk_regs));
 sg13g2_dfrbpq_1 _09410_ (.RESET_B(net487),
    .D(_00810_),
    .Q(\rf_ram.RAM[7][22] ),
    .CLK(clknet_leaf_66_clk_regs));
 sg13g2_dfrbpq_1 _09411_ (.RESET_B(net486),
    .D(_00811_),
    .Q(\rf_ram.RAM[7][23] ),
    .CLK(clknet_leaf_21_clk_regs));
 sg13g2_dfrbpq_1 _09412_ (.RESET_B(net485),
    .D(_00812_),
    .Q(\rf_ram.RAM[7][24] ),
    .CLK(clknet_leaf_69_clk_regs));
 sg13g2_dfrbpq_1 _09413_ (.RESET_B(net484),
    .D(_00813_),
    .Q(\rf_ram.RAM[7][25] ),
    .CLK(clknet_leaf_58_clk_regs));
 sg13g2_dfrbpq_1 _09414_ (.RESET_B(net483),
    .D(_00814_),
    .Q(\rf_ram.RAM[7][26] ),
    .CLK(clknet_leaf_57_clk_regs));
 sg13g2_dfrbpq_1 _09415_ (.RESET_B(net482),
    .D(_00815_),
    .Q(\rf_ram.RAM[7][27] ),
    .CLK(clknet_leaf_46_clk_regs));
 sg13g2_dfrbpq_1 _09416_ (.RESET_B(net481),
    .D(_00816_),
    .Q(\rf_ram.RAM[7][28] ),
    .CLK(clknet_leaf_24_clk_regs));
 sg13g2_dfrbpq_1 _09417_ (.RESET_B(net480),
    .D(_00817_),
    .Q(\rf_ram.RAM[7][29] ),
    .CLK(clknet_leaf_167_clk_regs));
 sg13g2_dfrbpq_1 _09418_ (.RESET_B(net479),
    .D(_00818_),
    .Q(\rf_ram.RAM[7][30] ),
    .CLK(clknet_leaf_162_clk_regs));
 sg13g2_dfrbpq_1 _09419_ (.RESET_B(net478),
    .D(_00819_),
    .Q(\rf_ram.RAM[7][31] ),
    .CLK(clknet_leaf_169_clk_regs));
 sg13g2_dfrbpq_1 _09420_ (.RESET_B(net477),
    .D(_00820_),
    .Q(\rf_ram.RAM[26][0] ),
    .CLK(clknet_leaf_17_clk_regs));
 sg13g2_dfrbpq_1 _09421_ (.RESET_B(net476),
    .D(_00821_),
    .Q(\rf_ram.RAM[26][1] ),
    .CLK(clknet_leaf_52_clk_regs));
 sg13g2_dfrbpq_1 _09422_ (.RESET_B(net475),
    .D(_00822_),
    .Q(\rf_ram.RAM[26][2] ),
    .CLK(clknet_leaf_75_clk_regs));
 sg13g2_dfrbpq_1 _09423_ (.RESET_B(net474),
    .D(_00823_),
    .Q(\rf_ram.RAM[26][3] ),
    .CLK(clknet_leaf_79_clk_regs));
 sg13g2_dfrbpq_1 _09424_ (.RESET_B(net473),
    .D(_00824_),
    .Q(\rf_ram.RAM[26][4] ),
    .CLK(clknet_leaf_83_clk_regs));
 sg13g2_dfrbpq_1 _09425_ (.RESET_B(net472),
    .D(_00825_),
    .Q(\rf_ram.RAM[26][5] ),
    .CLK(clknet_leaf_81_clk_regs));
 sg13g2_dfrbpq_1 _09426_ (.RESET_B(net471),
    .D(_00826_),
    .Q(\rf_ram.RAM[26][6] ),
    .CLK(clknet_leaf_90_clk_regs));
 sg13g2_dfrbpq_1 _09427_ (.RESET_B(net470),
    .D(_00827_),
    .Q(\rf_ram.RAM[26][7] ),
    .CLK(clknet_leaf_96_clk_regs));
 sg13g2_dfrbpq_1 _09428_ (.RESET_B(net469),
    .D(_00828_),
    .Q(\rf_ram.RAM[26][8] ),
    .CLK(clknet_leaf_114_clk_regs));
 sg13g2_dfrbpq_1 _09429_ (.RESET_B(net468),
    .D(_00829_),
    .Q(\rf_ram.RAM[26][9] ),
    .CLK(clknet_leaf_130_clk_regs));
 sg13g2_dfrbpq_1 _09430_ (.RESET_B(net467),
    .D(_00830_),
    .Q(\rf_ram.RAM[26][10] ),
    .CLK(clknet_leaf_119_clk_regs));
 sg13g2_dfrbpq_1 _09431_ (.RESET_B(net466),
    .D(_00831_),
    .Q(\rf_ram.RAM[26][11] ),
    .CLK(clknet_leaf_131_clk_regs));
 sg13g2_dfrbpq_1 _09432_ (.RESET_B(net465),
    .D(_00832_),
    .Q(\rf_ram.RAM[26][12] ),
    .CLK(clknet_leaf_122_clk_regs));
 sg13g2_dfrbpq_1 _09433_ (.RESET_B(net464),
    .D(_00833_),
    .Q(\rf_ram.RAM[26][13] ),
    .CLK(clknet_leaf_98_clk_regs));
 sg13g2_dfrbpq_1 _09434_ (.RESET_B(net463),
    .D(_00834_),
    .Q(\rf_ram.RAM[26][14] ),
    .CLK(clknet_leaf_158_clk_regs));
 sg13g2_dfrbpq_1 _09435_ (.RESET_B(net462),
    .D(_00835_),
    .Q(\rf_ram.RAM[26][15] ),
    .CLK(clknet_leaf_148_clk_regs));
 sg13g2_dfrbpq_1 _09436_ (.RESET_B(net461),
    .D(_00836_),
    .Q(\rf_ram.RAM[26][16] ),
    .CLK(clknet_leaf_107_clk_regs));
 sg13g2_dfrbpq_1 _09437_ (.RESET_B(net460),
    .D(_00837_),
    .Q(\rf_ram.RAM[26][17] ),
    .CLK(clknet_leaf_159_clk_regs));
 sg13g2_dfrbpq_1 _09438_ (.RESET_B(net459),
    .D(_00838_),
    .Q(\rf_ram.RAM[26][18] ),
    .CLK(clknet_leaf_142_clk_regs));
 sg13g2_dfrbpq_1 _09439_ (.RESET_B(net458),
    .D(_00839_),
    .Q(\rf_ram.RAM[26][19] ),
    .CLK(clknet_leaf_20_clk_regs));
 sg13g2_dfrbpq_1 _09440_ (.RESET_B(net457),
    .D(_00840_),
    .Q(\rf_ram.RAM[26][20] ),
    .CLK(clknet_leaf_149_clk_regs));
 sg13g2_dfrbpq_1 _09441_ (.RESET_B(net456),
    .D(_00841_),
    .Q(\rf_ram.RAM[26][21] ),
    .CLK(clknet_leaf_60_clk_regs));
 sg13g2_dfrbpq_1 _09442_ (.RESET_B(net455),
    .D(_00842_),
    .Q(\rf_ram.RAM[26][22] ),
    .CLK(clknet_leaf_70_clk_regs));
 sg13g2_dfrbpq_1 _09443_ (.RESET_B(net454),
    .D(_00843_),
    .Q(\rf_ram.RAM[26][23] ),
    .CLK(clknet_leaf_24_clk_regs));
 sg13g2_dfrbpq_1 _09444_ (.RESET_B(net453),
    .D(_00844_),
    .Q(\rf_ram.RAM[26][24] ),
    .CLK(clknet_leaf_74_clk_regs));
 sg13g2_dfrbpq_1 _09445_ (.RESET_B(net452),
    .D(_00845_),
    .Q(\rf_ram.RAM[26][25] ),
    .CLK(clknet_leaf_47_clk_regs));
 sg13g2_dfrbpq_1 _09446_ (.RESET_B(net451),
    .D(_00846_),
    .Q(\rf_ram.RAM[26][26] ),
    .CLK(clknet_leaf_54_clk_regs));
 sg13g2_dfrbpq_1 _09447_ (.RESET_B(net450),
    .D(_00847_),
    .Q(\rf_ram.RAM[26][27] ),
    .CLK(clknet_leaf_44_clk_regs));
 sg13g2_dfrbpq_1 _09448_ (.RESET_B(net449),
    .D(_00848_),
    .Q(\rf_ram.RAM[26][28] ),
    .CLK(clknet_leaf_27_clk_regs));
 sg13g2_dfrbpq_1 _09449_ (.RESET_B(net448),
    .D(_00849_),
    .Q(\rf_ram.RAM[26][29] ),
    .CLK(clknet_leaf_16_clk_regs));
 sg13g2_dfrbpq_1 _09450_ (.RESET_B(net447),
    .D(_00850_),
    .Q(\rf_ram.RAM[26][30] ),
    .CLK(clknet_leaf_164_clk_regs));
 sg13g2_dfrbpq_1 _09451_ (.RESET_B(net446),
    .D(_00851_),
    .Q(\rf_ram.RAM[26][31] ),
    .CLK(clknet_leaf_166_clk_regs));
 sg13g2_dfrbpq_1 _09452_ (.RESET_B(net445),
    .D(net2825),
    .Q(\rf_ram.RAM[6][0] ),
    .CLK(clknet_leaf_19_clk_regs));
 sg13g2_dfrbpq_1 _09453_ (.RESET_B(net444),
    .D(_00853_),
    .Q(\rf_ram.RAM[6][1] ),
    .CLK(clknet_leaf_55_clk_regs));
 sg13g2_dfrbpq_1 _09454_ (.RESET_B(net443),
    .D(_00854_),
    .Q(\rf_ram.RAM[6][2] ),
    .CLK(clknet_leaf_70_clk_regs));
 sg13g2_dfrbpq_1 _09455_ (.RESET_B(net442),
    .D(_00855_),
    .Q(\rf_ram.RAM[6][3] ),
    .CLK(clknet_leaf_89_clk_regs));
 sg13g2_dfrbpq_1 _09456_ (.RESET_B(net441),
    .D(_00856_),
    .Q(\rf_ram.RAM[6][4] ),
    .CLK(clknet_leaf_88_clk_regs));
 sg13g2_dfrbpq_1 _09457_ (.RESET_B(net440),
    .D(_00857_),
    .Q(\rf_ram.RAM[6][5] ),
    .CLK(clknet_leaf_91_clk_regs));
 sg13g2_dfrbpq_1 _09458_ (.RESET_B(net439),
    .D(_00858_),
    .Q(\rf_ram.RAM[6][6] ),
    .CLK(clknet_leaf_96_clk_regs));
 sg13g2_dfrbpq_1 _09459_ (.RESET_B(net438),
    .D(_00859_),
    .Q(\rf_ram.RAM[6][7] ),
    .CLK(clknet_leaf_99_clk_regs));
 sg13g2_dfrbpq_1 _09460_ (.RESET_B(net437),
    .D(_00860_),
    .Q(\rf_ram.RAM[6][8] ),
    .CLK(clknet_leaf_116_clk_regs));
 sg13g2_dfrbpq_1 _09461_ (.RESET_B(net436),
    .D(_00861_),
    .Q(\rf_ram.RAM[6][9] ),
    .CLK(clknet_leaf_127_clk_regs));
 sg13g2_dfrbpq_1 _09462_ (.RESET_B(net435),
    .D(_00862_),
    .Q(\rf_ram.RAM[6][10] ),
    .CLK(clknet_leaf_122_clk_regs));
 sg13g2_dfrbpq_1 _09463_ (.RESET_B(net434),
    .D(_00863_),
    .Q(\rf_ram.RAM[6][11] ),
    .CLK(clknet_leaf_134_clk_regs));
 sg13g2_dfrbpq_1 _09464_ (.RESET_B(net433),
    .D(_00864_),
    .Q(\rf_ram.RAM[6][12] ),
    .CLK(clknet_leaf_127_clk_regs));
 sg13g2_dfrbpq_1 _09465_ (.RESET_B(net432),
    .D(_00865_),
    .Q(\rf_ram.RAM[6][13] ),
    .CLK(clknet_leaf_143_clk_regs));
 sg13g2_dfrbpq_1 _09466_ (.RESET_B(net431),
    .D(_00866_),
    .Q(\rf_ram.RAM[6][14] ),
    .CLK(clknet_leaf_157_clk_regs));
 sg13g2_dfrbpq_1 _09467_ (.RESET_B(net430),
    .D(_00867_),
    .Q(\rf_ram.RAM[6][15] ),
    .CLK(clknet_leaf_144_clk_regs));
 sg13g2_dfrbpq_1 _09468_ (.RESET_B(net429),
    .D(_00868_),
    .Q(\rf_ram.RAM[6][16] ),
    .CLK(clknet_leaf_105_clk_regs));
 sg13g2_dfrbpq_1 _09469_ (.RESET_B(net428),
    .D(_00869_),
    .Q(\rf_ram.RAM[6][17] ),
    .CLK(clknet_leaf_159_clk_regs));
 sg13g2_dfrbpq_1 _09470_ (.RESET_B(net427),
    .D(_00870_),
    .Q(\rf_ram.RAM[6][18] ),
    .CLK(clknet_leaf_133_clk_regs));
 sg13g2_dfrbpq_1 _09471_ (.RESET_B(net426),
    .D(_00871_),
    .Q(\rf_ram.RAM[6][19] ),
    .CLK(clknet_leaf_161_clk_regs));
 sg13g2_dfrbpq_1 _09472_ (.RESET_B(net425),
    .D(_00872_),
    .Q(\rf_ram.RAM[6][20] ),
    .CLK(clknet_leaf_149_clk_regs));
 sg13g2_dfrbpq_1 _09473_ (.RESET_B(net424),
    .D(_00873_),
    .Q(\rf_ram.RAM[6][21] ),
    .CLK(clknet_leaf_60_clk_regs));
 sg13g2_dfrbpq_1 _09474_ (.RESET_B(net423),
    .D(_00874_),
    .Q(\rf_ram.RAM[6][22] ),
    .CLK(clknet_leaf_66_clk_regs));
 sg13g2_dfrbpq_1 _09475_ (.RESET_B(net422),
    .D(_00875_),
    .Q(\rf_ram.RAM[6][23] ),
    .CLK(clknet_leaf_20_clk_regs));
 sg13g2_dfrbpq_1 _09476_ (.RESET_B(net421),
    .D(_00876_),
    .Q(\rf_ram.RAM[6][24] ),
    .CLK(clknet_leaf_70_clk_regs));
 sg13g2_dfrbpq_1 _09477_ (.RESET_B(net420),
    .D(_00877_),
    .Q(\rf_ram.RAM[6][25] ),
    .CLK(clknet_leaf_58_clk_regs));
 sg13g2_dfrbpq_1 _09478_ (.RESET_B(net419),
    .D(_00878_),
    .Q(\rf_ram.RAM[6][26] ),
    .CLK(clknet_leaf_55_clk_regs));
 sg13g2_dfrbpq_1 _09479_ (.RESET_B(net418),
    .D(_00879_),
    .Q(\rf_ram.RAM[6][27] ),
    .CLK(clknet_leaf_46_clk_regs));
 sg13g2_dfrbpq_1 _09480_ (.RESET_B(net417),
    .D(_00880_),
    .Q(\rf_ram.RAM[6][28] ),
    .CLK(clknet_leaf_24_clk_regs));
 sg13g2_dfrbpq_1 _09481_ (.RESET_B(net416),
    .D(_00881_),
    .Q(\rf_ram.RAM[6][29] ),
    .CLK(clknet_leaf_170_clk_regs));
 sg13g2_dfrbpq_1 _09482_ (.RESET_B(net415),
    .D(_00882_),
    .Q(\rf_ram.RAM[6][30] ),
    .CLK(clknet_leaf_162_clk_regs));
 sg13g2_dfrbpq_1 _09483_ (.RESET_B(net414),
    .D(_00883_),
    .Q(\rf_ram.RAM[6][31] ),
    .CLK(clknet_leaf_169_clk_regs));
 sg13g2_dfrbpq_1 _09484_ (.RESET_B(net413),
    .D(_00884_),
    .Q(\rf_ram.RAM[25][0] ),
    .CLK(clknet_leaf_18_clk_regs));
 sg13g2_dfrbpq_1 _09485_ (.RESET_B(net412),
    .D(_00885_),
    .Q(\rf_ram.RAM[25][1] ),
    .CLK(clknet_leaf_52_clk_regs));
 sg13g2_dfrbpq_1 _09486_ (.RESET_B(net411),
    .D(_00886_),
    .Q(\rf_ram.RAM[25][2] ),
    .CLK(clknet_leaf_78_clk_regs));
 sg13g2_dfrbpq_1 _09487_ (.RESET_B(net410),
    .D(_00887_),
    .Q(\rf_ram.RAM[25][3] ),
    .CLK(clknet_leaf_78_clk_regs));
 sg13g2_dfrbpq_1 _09488_ (.RESET_B(net409),
    .D(_00888_),
    .Q(\rf_ram.RAM[25][4] ),
    .CLK(clknet_leaf_83_clk_regs));
 sg13g2_dfrbpq_1 _09489_ (.RESET_B(net408),
    .D(_00889_),
    .Q(\rf_ram.RAM[25][5] ),
    .CLK(clknet_leaf_81_clk_regs));
 sg13g2_dfrbpq_1 _09490_ (.RESET_B(net407),
    .D(_00890_),
    .Q(\rf_ram.RAM[25][6] ),
    .CLK(clknet_leaf_90_clk_regs));
 sg13g2_dfrbpq_1 _09491_ (.RESET_B(net406),
    .D(_00891_),
    .Q(\rf_ram.RAM[25][7] ),
    .CLK(clknet_leaf_96_clk_regs));
 sg13g2_dfrbpq_1 _09492_ (.RESET_B(net405),
    .D(_00892_),
    .Q(\rf_ram.RAM[25][8] ),
    .CLK(clknet_leaf_113_clk_regs));
 sg13g2_dfrbpq_1 _09493_ (.RESET_B(net404),
    .D(_00893_),
    .Q(\rf_ram.RAM[25][9] ),
    .CLK(clknet_leaf_130_clk_regs));
 sg13g2_dfrbpq_1 _09494_ (.RESET_B(net403),
    .D(_00894_),
    .Q(\rf_ram.RAM[25][10] ),
    .CLK(clknet_leaf_119_clk_regs));
 sg13g2_dfrbpq_1 _09495_ (.RESET_B(net402),
    .D(_00895_),
    .Q(\rf_ram.RAM[25][11] ),
    .CLK(clknet_leaf_131_clk_regs));
 sg13g2_dfrbpq_1 _09496_ (.RESET_B(net401),
    .D(_00896_),
    .Q(\rf_ram.RAM[25][12] ),
    .CLK(clknet_leaf_125_clk_regs));
 sg13g2_dfrbpq_1 _09497_ (.RESET_B(net400),
    .D(_00897_),
    .Q(\rf_ram.RAM[25][13] ),
    .CLK(clknet_leaf_98_clk_regs));
 sg13g2_dfrbpq_1 _09498_ (.RESET_B(net399),
    .D(_00898_),
    .Q(\rf_ram.RAM[25][14] ),
    .CLK(clknet_leaf_158_clk_regs));
 sg13g2_dfrbpq_1 _09499_ (.RESET_B(net398),
    .D(_00899_),
    .Q(\rf_ram.RAM[25][15] ),
    .CLK(clknet_leaf_107_clk_regs));
 sg13g2_dfrbpq_1 _09500_ (.RESET_B(net397),
    .D(_00900_),
    .Q(\rf_ram.RAM[25][16] ),
    .CLK(clknet_leaf_107_clk_regs));
 sg13g2_dfrbpq_1 _09501_ (.RESET_B(net396),
    .D(_00901_),
    .Q(\rf_ram.RAM[25][17] ),
    .CLK(clknet_leaf_159_clk_regs));
 sg13g2_dfrbpq_1 _09502_ (.RESET_B(net395),
    .D(_00902_),
    .Q(\rf_ram.RAM[25][18] ),
    .CLK(clknet_leaf_142_clk_regs));
 sg13g2_dfrbpq_1 _09503_ (.RESET_B(net394),
    .D(_00903_),
    .Q(\rf_ram.RAM[25][19] ),
    .CLK(clknet_leaf_21_clk_regs));
 sg13g2_dfrbpq_1 _09504_ (.RESET_B(net393),
    .D(_00904_),
    .Q(\rf_ram.RAM[25][20] ),
    .CLK(clknet_leaf_150_clk_regs));
 sg13g2_dfrbpq_1 _09505_ (.RESET_B(net392),
    .D(_00905_),
    .Q(\rf_ram.RAM[25][21] ),
    .CLK(clknet_leaf_60_clk_regs));
 sg13g2_dfrbpq_1 _09506_ (.RESET_B(net391),
    .D(_00906_),
    .Q(\rf_ram.RAM[25][22] ),
    .CLK(clknet_leaf_70_clk_regs));
 sg13g2_dfrbpq_1 _09507_ (.RESET_B(net390),
    .D(_00907_),
    .Q(\rf_ram.RAM[25][23] ),
    .CLK(clknet_leaf_18_clk_regs));
 sg13g2_dfrbpq_1 _09508_ (.RESET_B(net389),
    .D(_00908_),
    .Q(\rf_ram.RAM[25][24] ),
    .CLK(clknet_leaf_74_clk_regs));
 sg13g2_dfrbpq_1 _09509_ (.RESET_B(net388),
    .D(_00909_),
    .Q(\rf_ram.RAM[25][25] ),
    .CLK(clknet_leaf_47_clk_regs));
 sg13g2_dfrbpq_1 _09510_ (.RESET_B(net387),
    .D(_00910_),
    .Q(\rf_ram.RAM[25][26] ),
    .CLK(clknet_leaf_54_clk_regs));
 sg13g2_dfrbpq_1 _09511_ (.RESET_B(net386),
    .D(_00911_),
    .Q(\rf_ram.RAM[25][27] ),
    .CLK(clknet_leaf_44_clk_regs));
 sg13g2_dfrbpq_1 _09512_ (.RESET_B(net385),
    .D(_00912_),
    .Q(\rf_ram.RAM[25][28] ),
    .CLK(clknet_leaf_27_clk_regs));
 sg13g2_dfrbpq_1 _09513_ (.RESET_B(net384),
    .D(_00913_),
    .Q(\rf_ram.RAM[25][29] ),
    .CLK(clknet_leaf_16_clk_regs));
 sg13g2_dfrbpq_1 _09514_ (.RESET_B(net383),
    .D(_00914_),
    .Q(\rf_ram.RAM[25][30] ),
    .CLK(clknet_leaf_164_clk_regs));
 sg13g2_dfrbpq_1 _09515_ (.RESET_B(net382),
    .D(_00915_),
    .Q(\rf_ram.RAM[25][31] ),
    .CLK(clknet_leaf_167_clk_regs));
 sg13g2_dfrbpq_1 _09516_ (.RESET_B(net381),
    .D(net3143),
    .Q(\rf_ram.RAM[5][0] ),
    .CLK(clknet_leaf_19_clk_regs));
 sg13g2_dfrbpq_1 _09517_ (.RESET_B(net380),
    .D(_00917_),
    .Q(\rf_ram.RAM[5][1] ),
    .CLK(clknet_leaf_55_clk_regs));
 sg13g2_dfrbpq_1 _09518_ (.RESET_B(net379),
    .D(_00918_),
    .Q(\rf_ram.RAM[5][2] ),
    .CLK(clknet_leaf_69_clk_regs));
 sg13g2_dfrbpq_1 _09519_ (.RESET_B(net378),
    .D(_00919_),
    .Q(\rf_ram.RAM[5][3] ),
    .CLK(clknet_leaf_89_clk_regs));
 sg13g2_dfrbpq_1 _09520_ (.RESET_B(net377),
    .D(_00920_),
    .Q(\rf_ram.RAM[5][4] ),
    .CLK(clknet_leaf_89_clk_regs));
 sg13g2_dfrbpq_1 _09521_ (.RESET_B(net376),
    .D(_00921_),
    .Q(\rf_ram.RAM[5][5] ),
    .CLK(clknet_leaf_89_clk_regs));
 sg13g2_dfrbpq_1 _09522_ (.RESET_B(net375),
    .D(_00922_),
    .Q(\rf_ram.RAM[5][6] ),
    .CLK(clknet_leaf_96_clk_regs));
 sg13g2_dfrbpq_1 _09523_ (.RESET_B(net374),
    .D(_00923_),
    .Q(\rf_ram.RAM[5][7] ),
    .CLK(clknet_leaf_99_clk_regs));
 sg13g2_dfrbpq_1 _09524_ (.RESET_B(net373),
    .D(_00924_),
    .Q(\rf_ram.RAM[5][8] ),
    .CLK(clknet_leaf_117_clk_regs));
 sg13g2_dfrbpq_1 _09525_ (.RESET_B(net372),
    .D(_00925_),
    .Q(\rf_ram.RAM[5][9] ),
    .CLK(clknet_leaf_127_clk_regs));
 sg13g2_dfrbpq_1 _09526_ (.RESET_B(net371),
    .D(_00926_),
    .Q(\rf_ram.RAM[5][10] ),
    .CLK(clknet_leaf_123_clk_regs));
 sg13g2_dfrbpq_1 _09527_ (.RESET_B(net370),
    .D(_00927_),
    .Q(\rf_ram.RAM[5][11] ),
    .CLK(clknet_leaf_134_clk_regs));
 sg13g2_dfrbpq_1 _09528_ (.RESET_B(net369),
    .D(_00928_),
    .Q(\rf_ram.RAM[5][12] ),
    .CLK(clknet_leaf_127_clk_regs));
 sg13g2_dfrbpq_1 _09529_ (.RESET_B(net368),
    .D(_00929_),
    .Q(\rf_ram.RAM[5][13] ),
    .CLK(clknet_leaf_143_clk_regs));
 sg13g2_dfrbpq_1 _09530_ (.RESET_B(net367),
    .D(_00930_),
    .Q(\rf_ram.RAM[5][14] ),
    .CLK(clknet_leaf_157_clk_regs));
 sg13g2_dfrbpq_1 _09531_ (.RESET_B(net366),
    .D(_00931_),
    .Q(\rf_ram.RAM[5][15] ),
    .CLK(clknet_leaf_144_clk_regs));
 sg13g2_dfrbpq_1 _09532_ (.RESET_B(net365),
    .D(_00932_),
    .Q(\rf_ram.RAM[5][16] ),
    .CLK(clknet_leaf_105_clk_regs));
 sg13g2_dfrbpq_1 _09533_ (.RESET_B(net364),
    .D(_00933_),
    .Q(\rf_ram.RAM[5][17] ),
    .CLK(clknet_leaf_159_clk_regs));
 sg13g2_dfrbpq_1 _09534_ (.RESET_B(net363),
    .D(_00934_),
    .Q(\rf_ram.RAM[5][18] ),
    .CLK(clknet_leaf_134_clk_regs));
 sg13g2_dfrbpq_1 _09535_ (.RESET_B(net362),
    .D(_00935_),
    .Q(\rf_ram.RAM[5][19] ),
    .CLK(clknet_leaf_160_clk_regs));
 sg13g2_dfrbpq_1 _09536_ (.RESET_B(net361),
    .D(_00936_),
    .Q(\rf_ram.RAM[5][20] ),
    .CLK(clknet_leaf_150_clk_regs));
 sg13g2_dfrbpq_1 _09537_ (.RESET_B(net360),
    .D(_00937_),
    .Q(\rf_ram.RAM[5][21] ),
    .CLK(clknet_leaf_61_clk_regs));
 sg13g2_dfrbpq_1 _09538_ (.RESET_B(net359),
    .D(_00938_),
    .Q(\rf_ram.RAM[5][22] ),
    .CLK(clknet_leaf_64_clk_regs));
 sg13g2_dfrbpq_1 _09539_ (.RESET_B(net358),
    .D(_00939_),
    .Q(\rf_ram.RAM[5][23] ),
    .CLK(clknet_leaf_20_clk_regs));
 sg13g2_dfrbpq_1 _09540_ (.RESET_B(net357),
    .D(_00940_),
    .Q(\rf_ram.RAM[5][24] ),
    .CLK(clknet_leaf_69_clk_regs));
 sg13g2_dfrbpq_1 _09541_ (.RESET_B(net356),
    .D(net1675),
    .Q(\rf_ram.RAM[5][25] ),
    .CLK(clknet_leaf_58_clk_regs));
 sg13g2_dfrbpq_1 _09542_ (.RESET_B(net355),
    .D(_00942_),
    .Q(\rf_ram.RAM[5][26] ),
    .CLK(clknet_leaf_55_clk_regs));
 sg13g2_dfrbpq_1 _09543_ (.RESET_B(net354),
    .D(_00943_),
    .Q(\rf_ram.RAM[5][27] ),
    .CLK(clknet_leaf_46_clk_regs));
 sg13g2_dfrbpq_1 _09544_ (.RESET_B(net353),
    .D(_00944_),
    .Q(\rf_ram.RAM[5][28] ),
    .CLK(clknet_leaf_24_clk_regs));
 sg13g2_dfrbpq_1 _09545_ (.RESET_B(net352),
    .D(_00945_),
    .Q(\rf_ram.RAM[5][29] ),
    .CLK(clknet_leaf_169_clk_regs));
 sg13g2_dfrbpq_1 _09546_ (.RESET_B(net351),
    .D(_00946_),
    .Q(\rf_ram.RAM[5][30] ),
    .CLK(clknet_leaf_162_clk_regs));
 sg13g2_dfrbpq_1 _09547_ (.RESET_B(net350),
    .D(_00947_),
    .Q(\rf_ram.RAM[5][31] ),
    .CLK(clknet_leaf_169_clk_regs));
 sg13g2_dfrbpq_1 _09548_ (.RESET_B(net349),
    .D(_00948_),
    .Q(\rf_ram.RAM[24][0] ),
    .CLK(clknet_leaf_17_clk_regs));
 sg13g2_dfrbpq_1 _09549_ (.RESET_B(net348),
    .D(_00949_),
    .Q(\rf_ram.RAM[24][1] ),
    .CLK(clknet_leaf_52_clk_regs));
 sg13g2_dfrbpq_1 _09550_ (.RESET_B(net347),
    .D(_00950_),
    .Q(\rf_ram.RAM[24][2] ),
    .CLK(clknet_leaf_78_clk_regs));
 sg13g2_dfrbpq_1 _09551_ (.RESET_B(net346),
    .D(_00951_),
    .Q(\rf_ram.RAM[24][3] ),
    .CLK(clknet_leaf_79_clk_regs));
 sg13g2_dfrbpq_1 _09552_ (.RESET_B(net345),
    .D(_00952_),
    .Q(\rf_ram.RAM[24][4] ),
    .CLK(clknet_leaf_86_clk_regs));
 sg13g2_dfrbpq_1 _09553_ (.RESET_B(net344),
    .D(_00953_),
    .Q(\rf_ram.RAM[24][5] ),
    .CLK(clknet_leaf_86_clk_regs));
 sg13g2_dfrbpq_1 _09554_ (.RESET_B(net343),
    .D(_00954_),
    .Q(\rf_ram.RAM[24][6] ),
    .CLK(clknet_leaf_91_clk_regs));
 sg13g2_dfrbpq_1 _09555_ (.RESET_B(net342),
    .D(_00955_),
    .Q(\rf_ram.RAM[24][7] ),
    .CLK(clknet_leaf_94_clk_regs));
 sg13g2_dfrbpq_1 _09556_ (.RESET_B(net341),
    .D(_00956_),
    .Q(\rf_ram.RAM[24][8] ),
    .CLK(clknet_leaf_113_clk_regs));
 sg13g2_dfrbpq_1 _09557_ (.RESET_B(net340),
    .D(_00957_),
    .Q(\rf_ram.RAM[24][9] ),
    .CLK(clknet_leaf_122_clk_regs));
 sg13g2_dfrbpq_1 _09558_ (.RESET_B(net339),
    .D(_00958_),
    .Q(\rf_ram.RAM[24][10] ),
    .CLK(clknet_leaf_122_clk_regs));
 sg13g2_dfrbpq_1 _09559_ (.RESET_B(net338),
    .D(_00959_),
    .Q(\rf_ram.RAM[24][11] ),
    .CLK(clknet_leaf_131_clk_regs));
 sg13g2_dfrbpq_1 _09560_ (.RESET_B(net337),
    .D(_00960_),
    .Q(\rf_ram.RAM[24][12] ),
    .CLK(clknet_leaf_125_clk_regs));
 sg13g2_dfrbpq_1 _09561_ (.RESET_B(net336),
    .D(_00961_),
    .Q(\rf_ram.RAM[24][13] ),
    .CLK(clknet_leaf_113_clk_regs));
 sg13g2_dfrbpq_1 _09562_ (.RESET_B(net335),
    .D(_00962_),
    .Q(\rf_ram.RAM[24][14] ),
    .CLK(clknet_leaf_158_clk_regs));
 sg13g2_dfrbpq_1 _09563_ (.RESET_B(net334),
    .D(_00963_),
    .Q(\rf_ram.RAM[24][15] ),
    .CLK(clknet_leaf_148_clk_regs));
 sg13g2_dfrbpq_1 _09564_ (.RESET_B(net333),
    .D(_00964_),
    .Q(\rf_ram.RAM[24][16] ),
    .CLK(clknet_leaf_108_clk_regs));
 sg13g2_dfrbpq_1 _09565_ (.RESET_B(net332),
    .D(_00965_),
    .Q(\rf_ram.RAM[24][17] ),
    .CLK(clknet_leaf_159_clk_regs));
 sg13g2_dfrbpq_1 _09566_ (.RESET_B(net331),
    .D(_00966_),
    .Q(\rf_ram.RAM[24][18] ),
    .CLK(clknet_leaf_142_clk_regs));
 sg13g2_dfrbpq_1 _09567_ (.RESET_B(net330),
    .D(_00967_),
    .Q(\rf_ram.RAM[24][19] ),
    .CLK(clknet_leaf_21_clk_regs));
 sg13g2_dfrbpq_1 _09568_ (.RESET_B(net329),
    .D(_00968_),
    .Q(\rf_ram.RAM[24][20] ),
    .CLK(clknet_leaf_149_clk_regs));
 sg13g2_dfrbpq_1 _09569_ (.RESET_B(net328),
    .D(_00969_),
    .Q(\rf_ram.RAM[24][21] ),
    .CLK(clknet_leaf_70_clk_regs));
 sg13g2_dfrbpq_1 _09570_ (.RESET_B(net327),
    .D(_00970_),
    .Q(\rf_ram.RAM[24][22] ),
    .CLK(clknet_leaf_70_clk_regs));
 sg13g2_dfrbpq_1 _09571_ (.RESET_B(net326),
    .D(_00971_),
    .Q(\rf_ram.RAM[24][23] ),
    .CLK(clknet_leaf_24_clk_regs));
 sg13g2_dfrbpq_1 _09572_ (.RESET_B(net325),
    .D(_00972_),
    .Q(\rf_ram.RAM[24][24] ),
    .CLK(clknet_leaf_72_clk_regs));
 sg13g2_dfrbpq_1 _09573_ (.RESET_B(net324),
    .D(_00973_),
    .Q(\rf_ram.RAM[24][25] ),
    .CLK(clknet_leaf_49_clk_regs));
 sg13g2_dfrbpq_1 _09574_ (.RESET_B(net323),
    .D(_00974_),
    .Q(\rf_ram.RAM[24][26] ),
    .CLK(clknet_leaf_71_clk_regs));
 sg13g2_dfrbpq_1 _09575_ (.RESET_B(net322),
    .D(_00975_),
    .Q(\rf_ram.RAM[24][27] ),
    .CLK(clknet_leaf_43_clk_regs));
 sg13g2_dfrbpq_1 _09576_ (.RESET_B(net321),
    .D(_00976_),
    .Q(\rf_ram.RAM[24][28] ),
    .CLK(clknet_leaf_35_clk_regs));
 sg13g2_dfrbpq_1 _09577_ (.RESET_B(net320),
    .D(_00977_),
    .Q(\rf_ram.RAM[24][29] ),
    .CLK(clknet_leaf_15_clk_regs));
 sg13g2_dfrbpq_1 _09578_ (.RESET_B(net319),
    .D(_00978_),
    .Q(\rf_ram.RAM[24][30] ),
    .CLK(clknet_leaf_164_clk_regs));
 sg13g2_dfrbpq_1 _09579_ (.RESET_B(net318),
    .D(_00979_),
    .Q(\rf_ram.RAM[24][31] ),
    .CLK(clknet_leaf_168_clk_regs));
 sg13g2_dfrbpq_1 _09580_ (.RESET_B(net317),
    .D(net3198),
    .Q(\rf_ram.RAM[30][0] ),
    .CLK(clknet_leaf_155_clk_regs));
 sg13g2_dfrbpq_1 _09581_ (.RESET_B(net316),
    .D(_00981_),
    .Q(\rf_ram.RAM[30][1] ),
    .CLK(clknet_leaf_52_clk_regs));
 sg13g2_dfrbpq_1 _09582_ (.RESET_B(net315),
    .D(_00982_),
    .Q(\rf_ram.RAM[30][2] ),
    .CLK(clknet_leaf_68_clk_regs));
 sg13g2_dfrbpq_1 _09583_ (.RESET_B(net314),
    .D(_00983_),
    .Q(\rf_ram.RAM[30][3] ),
    .CLK(clknet_leaf_86_clk_regs));
 sg13g2_dfrbpq_1 _09584_ (.RESET_B(net313),
    .D(_00984_),
    .Q(\rf_ram.RAM[30][4] ),
    .CLK(clknet_leaf_87_clk_regs));
 sg13g2_dfrbpq_1 _09585_ (.RESET_B(net312),
    .D(_00985_),
    .Q(\rf_ram.RAM[30][5] ),
    .CLK(clknet_leaf_92_clk_regs));
 sg13g2_dfrbpq_1 _09586_ (.RESET_B(net311),
    .D(_00986_),
    .Q(\rf_ram.RAM[30][6] ),
    .CLK(clknet_leaf_93_clk_regs));
 sg13g2_dfrbpq_1 _09587_ (.RESET_B(net310),
    .D(_00987_),
    .Q(\rf_ram.RAM[30][7] ),
    .CLK(clknet_leaf_95_clk_regs));
 sg13g2_dfrbpq_1 _09588_ (.RESET_B(net309),
    .D(_00988_),
    .Q(\rf_ram.RAM[30][8] ),
    .CLK(clknet_leaf_116_clk_regs));
 sg13g2_dfrbpq_1 _09589_ (.RESET_B(net308),
    .D(_00989_),
    .Q(\rf_ram.RAM[30][9] ),
    .CLK(clknet_leaf_124_clk_regs));
 sg13g2_dfrbpq_1 _09590_ (.RESET_B(net307),
    .D(_00990_),
    .Q(\rf_ram.RAM[30][10] ),
    .CLK(clknet_leaf_118_clk_regs));
 sg13g2_dfrbpq_1 _09591_ (.RESET_B(net306),
    .D(_00991_),
    .Q(\rf_ram.RAM[30][11] ),
    .CLK(clknet_leaf_135_clk_regs));
 sg13g2_dfrbpq_1 _09592_ (.RESET_B(net305),
    .D(_00992_),
    .Q(\rf_ram.RAM[30][12] ),
    .CLK(clknet_leaf_123_clk_regs));
 sg13g2_dfrbpq_1 _09593_ (.RESET_B(net304),
    .D(_00993_),
    .Q(\rf_ram.RAM[30][13] ),
    .CLK(clknet_leaf_90_clk_regs));
 sg13g2_dfrbpq_1 _09594_ (.RESET_B(net303),
    .D(_00994_),
    .Q(\rf_ram.RAM[30][14] ),
    .CLK(clknet_leaf_140_clk_regs));
 sg13g2_dfrbpq_1 _09595_ (.RESET_B(net302),
    .D(_00995_),
    .Q(\rf_ram.RAM[30][15] ),
    .CLK(clknet_leaf_109_clk_regs));
 sg13g2_dfrbpq_1 _09596_ (.RESET_B(net301),
    .D(_00996_),
    .Q(\rf_ram.RAM[30][16] ),
    .CLK(clknet_leaf_107_clk_regs));
 sg13g2_dfrbpq_1 _09597_ (.RESET_B(net300),
    .D(_00997_),
    .Q(\rf_ram.RAM[30][17] ),
    .CLK(clknet_leaf_139_clk_regs));
 sg13g2_dfrbpq_1 _09598_ (.RESET_B(net299),
    .D(_00998_),
    .Q(\rf_ram.RAM[30][18] ),
    .CLK(clknet_leaf_135_clk_regs));
 sg13g2_dfrbpq_1 _09599_ (.RESET_B(net298),
    .D(_00999_),
    .Q(\rf_ram.RAM[30][19] ),
    .CLK(clknet_leaf_155_clk_regs));
 sg13g2_dfrbpq_1 _09600_ (.RESET_B(net297),
    .D(_01000_),
    .Q(\rf_ram.RAM[30][20] ),
    .CLK(clknet_leaf_151_clk_regs));
 sg13g2_dfrbpq_1 _09601_ (.RESET_B(net296),
    .D(_01001_),
    .Q(\rf_ram.RAM[30][21] ),
    .CLK(clknet_leaf_65_clk_regs));
 sg13g2_dfrbpq_1 _09602_ (.RESET_B(net295),
    .D(_01002_),
    .Q(\rf_ram.RAM[30][22] ),
    .CLK(clknet_leaf_102_clk_regs));
 sg13g2_dfrbpq_1 _09603_ (.RESET_B(net294),
    .D(_01003_),
    .Q(\rf_ram.RAM[30][23] ),
    .CLK(clknet_leaf_59_clk_regs));
 sg13g2_dfrbpq_1 _09604_ (.RESET_B(net293),
    .D(_01004_),
    .Q(\rf_ram.RAM[30][24] ),
    .CLK(clknet_leaf_73_clk_regs));
 sg13g2_dfrbpq_1 _09605_ (.RESET_B(net292),
    .D(_01005_),
    .Q(\rf_ram.RAM[30][25] ),
    .CLK(clknet_leaf_50_clk_regs));
 sg13g2_dfrbpq_1 _09606_ (.RESET_B(net291),
    .D(_01006_),
    .Q(\rf_ram.RAM[30][26] ),
    .CLK(clknet_leaf_51_clk_regs));
 sg13g2_dfrbpq_1 _09607_ (.RESET_B(net290),
    .D(_01007_),
    .Q(\rf_ram.RAM[30][27] ),
    .CLK(clknet_leaf_43_clk_regs));
 sg13g2_dfrbpq_1 _09608_ (.RESET_B(net289),
    .D(_01008_),
    .Q(\rf_ram.RAM[30][28] ),
    .CLK(clknet_leaf_25_clk_regs));
 sg13g2_dfrbpq_1 _09609_ (.RESET_B(net288),
    .D(_01009_),
    .Q(\rf_ram.RAM[30][29] ),
    .CLK(clknet_leaf_154_clk_regs));
 sg13g2_dfrbpq_1 _09610_ (.RESET_B(net287),
    .D(_01010_),
    .Q(\rf_ram.RAM[30][30] ),
    .CLK(clknet_leaf_163_clk_regs));
 sg13g2_dfrbpq_1 _09611_ (.RESET_B(net286),
    .D(_01011_),
    .Q(\rf_ram.RAM[30][31] ),
    .CLK(clknet_leaf_168_clk_regs));
 sg13g2_dfrbpq_1 _09612_ (.RESET_B(net285),
    .D(net3595),
    .Q(\cpu.arbiter.i_wb_mem_rdt[0] ),
    .CLK(clknet_leaf_41_clk_regs));
 sg13g2_dfrbpq_1 _09613_ (.RESET_B(net284),
    .D(_01013_),
    .Q(\cpu.arbiter.i_wb_mem_rdt[1] ),
    .CLK(clknet_leaf_41_clk_regs));
 sg13g2_dfrbpq_2 _09614_ (.RESET_B(net283),
    .D(net3638),
    .Q(\cpu.arbiter.i_wb_mem_rdt[2] ),
    .CLK(clknet_leaf_41_clk_regs));
 sg13g2_dfrbpq_2 _09615_ (.RESET_B(net282),
    .D(_01015_),
    .Q(\cpu.arbiter.i_wb_mem_rdt[3] ),
    .CLK(clknet_leaf_41_clk_regs));
 sg13g2_dfrbpq_2 _09616_ (.RESET_B(net281),
    .D(_01016_),
    .Q(\cpu.arbiter.i_wb_mem_rdt[4] ),
    .CLK(clknet_leaf_39_clk_regs));
 sg13g2_dfrbpq_2 _09617_ (.RESET_B(net280),
    .D(net3679),
    .Q(\cpu.arbiter.i_wb_mem_rdt[5] ),
    .CLK(clknet_leaf_39_clk_regs));
 sg13g2_dfrbpq_2 _09618_ (.RESET_B(net279),
    .D(_01018_),
    .Q(\cpu.arbiter.i_wb_mem_rdt[6] ),
    .CLK(clknet_leaf_38_clk_regs));
 sg13g2_dfrbpq_2 _09619_ (.RESET_B(net278),
    .D(net3750),
    .Q(\cpu.arbiter.i_wb_mem_rdt[7] ),
    .CLK(clknet_leaf_38_clk_regs));
 sg13g2_dfrbpq_2 _09620_ (.RESET_B(net277),
    .D(net3693),
    .Q(\cpu.arbiter.i_wb_mem_rdt[8] ),
    .CLK(clknet_leaf_30_clk_regs));
 sg13g2_dfrbpq_1 _09621_ (.RESET_B(net276),
    .D(_01021_),
    .Q(\cpu.arbiter.i_wb_mem_rdt[9] ),
    .CLK(clknet_leaf_30_clk_regs));
 sg13g2_dfrbpq_1 _09622_ (.RESET_B(net275),
    .D(net3627),
    .Q(\cpu.arbiter.i_wb_mem_rdt[10] ),
    .CLK(clknet_leaf_11_clk_regs));
 sg13g2_dfrbpq_1 _09623_ (.RESET_B(net274),
    .D(_01023_),
    .Q(\cpu.arbiter.i_wb_mem_rdt[11] ),
    .CLK(clknet_leaf_10_clk_regs));
 sg13g2_dfrbpq_2 _09624_ (.RESET_B(net273),
    .D(_01024_),
    .Q(\cpu.arbiter.i_wb_mem_rdt[12] ),
    .CLK(clknet_leaf_9_clk_regs));
 sg13g2_dfrbpq_2 _09625_ (.RESET_B(net272),
    .D(net3695),
    .Q(\cpu.arbiter.i_wb_mem_rdt[13] ),
    .CLK(clknet_leaf_8_clk_regs));
 sg13g2_dfrbpq_2 _09626_ (.RESET_B(net271),
    .D(net3629),
    .Q(\cpu.arbiter.i_wb_mem_rdt[14] ),
    .CLK(clknet_leaf_9_clk_regs));
 sg13g2_dfrbpq_2 _09627_ (.RESET_B(net270),
    .D(_01027_),
    .Q(\cpu.arbiter.i_wb_mem_rdt[15] ),
    .CLK(clknet_leaf_11_clk_regs));
 sg13g2_dfrbpq_1 _09628_ (.RESET_B(net269),
    .D(net1573),
    .Q(\rf_ram.RAM[2][0] ),
    .CLK(clknet_leaf_14_clk_regs));
 sg13g2_dfrbpq_1 _09629_ (.RESET_B(net268),
    .D(_01029_),
    .Q(\rf_ram.RAM[2][1] ),
    .CLK(clknet_leaf_53_clk_regs));
 sg13g2_dfrbpq_1 _09630_ (.RESET_B(net267),
    .D(_01030_),
    .Q(\rf_ram.RAM[2][2] ),
    .CLK(clknet_leaf_76_clk_regs));
 sg13g2_dfrbpq_1 _09631_ (.RESET_B(net266),
    .D(_01031_),
    .Q(\rf_ram.RAM[2][3] ),
    .CLK(clknet_leaf_79_clk_regs));
 sg13g2_dfrbpq_1 _09632_ (.RESET_B(net265),
    .D(_01032_),
    .Q(\rf_ram.RAM[2][4] ),
    .CLK(clknet_leaf_82_clk_regs));
 sg13g2_dfrbpq_1 _09633_ (.RESET_B(net264),
    .D(_01033_),
    .Q(\rf_ram.RAM[2][5] ),
    .CLK(clknet_leaf_83_clk_regs));
 sg13g2_dfrbpq_1 _09634_ (.RESET_B(net263),
    .D(_01034_),
    .Q(\rf_ram.RAM[2][6] ),
    .CLK(clknet_leaf_101_clk_regs));
 sg13g2_dfrbpq_1 _09635_ (.RESET_B(net262),
    .D(_01035_),
    .Q(\rf_ram.RAM[2][7] ),
    .CLK(clknet_leaf_100_clk_regs));
 sg13g2_dfrbpq_1 _09636_ (.RESET_B(net261),
    .D(_01036_),
    .Q(\rf_ram.RAM[2][8] ),
    .CLK(clknet_leaf_114_clk_regs));
 sg13g2_dfrbpq_1 _09637_ (.RESET_B(net260),
    .D(_01037_),
    .Q(\rf_ram.RAM[2][9] ),
    .CLK(clknet_leaf_128_clk_regs));
 sg13g2_dfrbpq_1 _09638_ (.RESET_B(net259),
    .D(_01038_),
    .Q(\rf_ram.RAM[2][10] ),
    .CLK(clknet_leaf_121_clk_regs));
 sg13g2_dfrbpq_1 _09639_ (.RESET_B(net258),
    .D(_01039_),
    .Q(\rf_ram.RAM[2][11] ),
    .CLK(clknet_leaf_129_clk_regs));
 sg13g2_dfrbpq_1 _09640_ (.RESET_B(net257),
    .D(_01040_),
    .Q(\rf_ram.RAM[2][12] ),
    .CLK(clknet_leaf_128_clk_regs));
 sg13g2_dfrbpq_1 _09641_ (.RESET_B(net256),
    .D(_01041_),
    .Q(\rf_ram.RAM[2][13] ),
    .CLK(clknet_leaf_110_clk_regs));
 sg13g2_dfrbpq_1 _09642_ (.RESET_B(net255),
    .D(_01042_),
    .Q(\rf_ram.RAM[2][14] ),
    .CLK(clknet_leaf_158_clk_regs));
 sg13g2_dfrbpq_1 _09643_ (.RESET_B(net254),
    .D(_01043_),
    .Q(\rf_ram.RAM[2][15] ),
    .CLK(clknet_leaf_148_clk_regs));
 sg13g2_dfrbpq_1 _09644_ (.RESET_B(net253),
    .D(_01044_),
    .Q(\rf_ram.RAM[2][16] ),
    .CLK(clknet_leaf_102_clk_regs));
 sg13g2_dfrbpq_1 _09645_ (.RESET_B(net252),
    .D(_01045_),
    .Q(\rf_ram.RAM[2][17] ),
    .CLK(clknet_leaf_137_clk_regs));
 sg13g2_dfrbpq_1 _09646_ (.RESET_B(net251),
    .D(_01046_),
    .Q(\rf_ram.RAM[2][18] ),
    .CLK(clknet_leaf_136_clk_regs));
 sg13g2_dfrbpq_1 _09647_ (.RESET_B(net250),
    .D(_01047_),
    .Q(\rf_ram.RAM[2][19] ),
    .CLK(clknet_leaf_156_clk_regs));
 sg13g2_dfrbpq_1 _09648_ (.RESET_B(net249),
    .D(_01048_),
    .Q(\rf_ram.RAM[2][20] ),
    .CLK(clknet_leaf_20_clk_regs));
 sg13g2_dfrbpq_1 _09649_ (.RESET_B(net248),
    .D(_01049_),
    .Q(\rf_ram.RAM[2][21] ),
    .CLK(clknet_leaf_61_clk_regs));
 sg13g2_dfrbpq_1 _09650_ (.RESET_B(net247),
    .D(_01050_),
    .Q(\rf_ram.RAM[2][22] ),
    .CLK(clknet_leaf_64_clk_regs));
 sg13g2_dfrbpq_1 _09651_ (.RESET_B(net246),
    .D(_01051_),
    .Q(\rf_ram.RAM[2][23] ),
    .CLK(clknet_leaf_17_clk_regs));
 sg13g2_dfrbpq_1 _09652_ (.RESET_B(net245),
    .D(_01052_),
    .Q(\rf_ram.RAM[2][24] ),
    .CLK(clknet_leaf_74_clk_regs));
 sg13g2_dfrbpq_1 _09653_ (.RESET_B(net244),
    .D(_01053_),
    .Q(\rf_ram.RAM[2][25] ),
    .CLK(clknet_leaf_47_clk_regs));
 sg13g2_dfrbpq_1 _09654_ (.RESET_B(net243),
    .D(_01054_),
    .Q(\rf_ram.RAM[2][26] ),
    .CLK(clknet_leaf_56_clk_regs));
 sg13g2_dfrbpq_1 _09655_ (.RESET_B(net242),
    .D(_01055_),
    .Q(\rf_ram.RAM[2][27] ),
    .CLK(clknet_leaf_45_clk_regs));
 sg13g2_dfrbpq_1 _09656_ (.RESET_B(net241),
    .D(_01056_),
    .Q(\rf_ram.RAM[2][28] ),
    .CLK(clknet_leaf_27_clk_regs));
 sg13g2_dfrbpq_1 _09657_ (.RESET_B(net240),
    .D(_01057_),
    .Q(\rf_ram.RAM[2][29] ),
    .CLK(clknet_leaf_170_clk_regs));
 sg13g2_dfrbpq_1 _09658_ (.RESET_B(net239),
    .D(_01058_),
    .Q(\rf_ram.RAM[2][30] ),
    .CLK(clknet_leaf_168_clk_regs));
 sg13g2_dfrbpq_1 _09659_ (.RESET_B(net238),
    .D(_01059_),
    .Q(\rf_ram.RAM[2][31] ),
    .CLK(clknet_leaf_3_clk_regs));
 sg13g2_dfrbpq_1 _09660_ (.RESET_B(net237),
    .D(net2720),
    .Q(\rf_ram.RAM[28][0] ),
    .CLK(clknet_leaf_154_clk_regs));
 sg13g2_dfrbpq_1 _09661_ (.RESET_B(net236),
    .D(_01061_),
    .Q(\rf_ram.RAM[28][1] ),
    .CLK(clknet_leaf_52_clk_regs));
 sg13g2_dfrbpq_1 _09662_ (.RESET_B(net235),
    .D(_01062_),
    .Q(\rf_ram.RAM[28][2] ),
    .CLK(clknet_leaf_78_clk_regs));
 sg13g2_dfrbpq_1 _09663_ (.RESET_B(net234),
    .D(_01063_),
    .Q(\rf_ram.RAM[28][3] ),
    .CLK(clknet_leaf_86_clk_regs));
 sg13g2_dfrbpq_1 _09664_ (.RESET_B(net233),
    .D(_01064_),
    .Q(\rf_ram.RAM[28][4] ),
    .CLK(clknet_leaf_86_clk_regs));
 sg13g2_dfrbpq_1 _09665_ (.RESET_B(net232),
    .D(_01065_),
    .Q(\rf_ram.RAM[28][5] ),
    .CLK(clknet_leaf_92_clk_regs));
 sg13g2_dfrbpq_1 _09666_ (.RESET_B(net231),
    .D(_01066_),
    .Q(\rf_ram.RAM[28][6] ),
    .CLK(clknet_leaf_93_clk_regs));
 sg13g2_dfrbpq_1 _09667_ (.RESET_B(net230),
    .D(_01067_),
    .Q(\rf_ram.RAM[28][7] ),
    .CLK(clknet_leaf_93_clk_regs));
 sg13g2_dfrbpq_1 _09668_ (.RESET_B(net229),
    .D(_01068_),
    .Q(\rf_ram.RAM[28][8] ),
    .CLK(clknet_leaf_116_clk_regs));
 sg13g2_dfrbpq_1 _09669_ (.RESET_B(net228),
    .D(_01069_),
    .Q(\rf_ram.RAM[28][9] ),
    .CLK(clknet_leaf_124_clk_regs));
 sg13g2_dfrbpq_1 _09670_ (.RESET_B(net227),
    .D(_01070_),
    .Q(\rf_ram.RAM[28][10] ),
    .CLK(clknet_leaf_117_clk_regs));
 sg13g2_dfrbpq_1 _09671_ (.RESET_B(net226),
    .D(_01071_),
    .Q(\rf_ram.RAM[28][11] ),
    .CLK(clknet_leaf_134_clk_regs));
 sg13g2_dfrbpq_1 _09672_ (.RESET_B(net225),
    .D(_01072_),
    .Q(\rf_ram.RAM[28][12] ),
    .CLK(clknet_leaf_123_clk_regs));
 sg13g2_dfrbpq_1 _09673_ (.RESET_B(net224),
    .D(_01073_),
    .Q(\rf_ram.RAM[28][13] ),
    .CLK(clknet_leaf_101_clk_regs));
 sg13g2_dfrbpq_1 _09674_ (.RESET_B(net223),
    .D(_01074_),
    .Q(\rf_ram.RAM[28][14] ),
    .CLK(clknet_leaf_141_clk_regs));
 sg13g2_dfrbpq_1 _09675_ (.RESET_B(net222),
    .D(_01075_),
    .Q(\rf_ram.RAM[28][15] ),
    .CLK(clknet_leaf_109_clk_regs));
 sg13g2_dfrbpq_1 _09676_ (.RESET_B(net221),
    .D(_01076_),
    .Q(\rf_ram.RAM[28][16] ),
    .CLK(clknet_leaf_109_clk_regs));
 sg13g2_dfrbpq_1 _09677_ (.RESET_B(net220),
    .D(_01077_),
    .Q(\rf_ram.RAM[28][17] ),
    .CLK(clknet_leaf_138_clk_regs));
 sg13g2_dfrbpq_1 _09678_ (.RESET_B(net219),
    .D(_01078_),
    .Q(\rf_ram.RAM[28][18] ),
    .CLK(clknet_leaf_135_clk_regs));
 sg13g2_dfrbpq_1 _09679_ (.RESET_B(net218),
    .D(_01079_),
    .Q(\rf_ram.RAM[28][19] ),
    .CLK(clknet_leaf_155_clk_regs));
 sg13g2_dfrbpq_1 _09680_ (.RESET_B(net217),
    .D(_01080_),
    .Q(\rf_ram.RAM[28][20] ),
    .CLK(clknet_leaf_152_clk_regs));
 sg13g2_dfrbpq_1 _09681_ (.RESET_B(net216),
    .D(_01081_),
    .Q(\rf_ram.RAM[28][21] ),
    .CLK(clknet_leaf_63_clk_regs));
 sg13g2_dfrbpq_1 _09682_ (.RESET_B(net215),
    .D(_01082_),
    .Q(\rf_ram.RAM[28][22] ),
    .CLK(clknet_leaf_67_clk_regs));
 sg13g2_dfrbpq_1 _09683_ (.RESET_B(net214),
    .D(_01083_),
    .Q(\rf_ram.RAM[28][23] ),
    .CLK(clknet_leaf_59_clk_regs));
 sg13g2_dfrbpq_1 _09684_ (.RESET_B(net213),
    .D(_01084_),
    .Q(\rf_ram.RAM[28][24] ),
    .CLK(clknet_leaf_73_clk_regs));
 sg13g2_dfrbpq_1 _09685_ (.RESET_B(net212),
    .D(_01085_),
    .Q(\rf_ram.RAM[28][25] ),
    .CLK(clknet_leaf_49_clk_regs));
 sg13g2_dfrbpq_1 _09686_ (.RESET_B(net211),
    .D(_01086_),
    .Q(\rf_ram.RAM[28][26] ),
    .CLK(clknet_leaf_51_clk_regs));
 sg13g2_dfrbpq_1 _09687_ (.RESET_B(net210),
    .D(_01087_),
    .Q(\rf_ram.RAM[28][27] ),
    .CLK(clknet_leaf_48_clk_regs));
 sg13g2_dfrbpq_1 _09688_ (.RESET_B(net209),
    .D(_01088_),
    .Q(\rf_ram.RAM[28][28] ),
    .CLK(clknet_leaf_26_clk_regs));
 sg13g2_dfrbpq_1 _09689_ (.RESET_B(net208),
    .D(_01089_),
    .Q(\rf_ram.RAM[28][29] ),
    .CLK(clknet_leaf_154_clk_regs));
 sg13g2_dfrbpq_1 _09690_ (.RESET_B(net207),
    .D(_01090_),
    .Q(\rf_ram.RAM[28][30] ),
    .CLK(clknet_leaf_163_clk_regs));
 sg13g2_dfrbpq_1 _09691_ (.RESET_B(net206),
    .D(_01091_),
    .Q(\rf_ram.RAM[28][31] ),
    .CLK(clknet_leaf_168_clk_regs));
 sg13g2_dfrbpq_1 _09692_ (.RESET_B(net205),
    .D(net2712),
    .Q(\rf_ram.RAM[13][0] ),
    .CLK(clknet_leaf_17_clk_regs));
 sg13g2_dfrbpq_1 _09693_ (.RESET_B(net204),
    .D(_01093_),
    .Q(\rf_ram.RAM[13][1] ),
    .CLK(clknet_leaf_52_clk_regs));
 sg13g2_dfrbpq_1 _09694_ (.RESET_B(net203),
    .D(_01094_),
    .Q(\rf_ram.RAM[13][2] ),
    .CLK(clknet_leaf_77_clk_regs));
 sg13g2_dfrbpq_1 _09695_ (.RESET_B(net202),
    .D(_01095_),
    .Q(\rf_ram.RAM[13][3] ),
    .CLK(clknet_leaf_84_clk_regs));
 sg13g2_dfrbpq_1 _09696_ (.RESET_B(net201),
    .D(_01096_),
    .Q(\rf_ram.RAM[13][4] ),
    .CLK(clknet_leaf_82_clk_regs));
 sg13g2_dfrbpq_1 _09697_ (.RESET_B(net200),
    .D(_01097_),
    .Q(\rf_ram.RAM[13][5] ),
    .CLK(clknet_leaf_85_clk_regs));
 sg13g2_dfrbpq_1 _09698_ (.RESET_B(net199),
    .D(_01098_),
    .Q(\rf_ram.RAM[13][6] ),
    .CLK(clknet_leaf_94_clk_regs));
 sg13g2_dfrbpq_1 _09699_ (.RESET_B(net198),
    .D(_01099_),
    .Q(\rf_ram.RAM[13][7] ),
    .CLK(clknet_leaf_96_clk_regs));
 sg13g2_dfrbpq_1 _09700_ (.RESET_B(net197),
    .D(_01100_),
    .Q(\rf_ram.RAM[13][8] ),
    .CLK(clknet_leaf_114_clk_regs));
 sg13g2_dfrbpq_1 _09701_ (.RESET_B(net196),
    .D(_01101_),
    .Q(\rf_ram.RAM[13][9] ),
    .CLK(clknet_leaf_124_clk_regs));
 sg13g2_dfrbpq_1 _09702_ (.RESET_B(net195),
    .D(_01102_),
    .Q(\rf_ram.RAM[13][10] ),
    .CLK(clknet_leaf_120_clk_regs));
 sg13g2_dfrbpq_1 _09703_ (.RESET_B(net194),
    .D(_01103_),
    .Q(\rf_ram.RAM[13][11] ),
    .CLK(clknet_leaf_131_clk_regs));
 sg13g2_dfrbpq_1 _09704_ (.RESET_B(net193),
    .D(_01104_),
    .Q(\rf_ram.RAM[13][12] ),
    .CLK(clknet_leaf_123_clk_regs));
 sg13g2_dfrbpq_1 _09705_ (.RESET_B(net192),
    .D(_01105_),
    .Q(\rf_ram.RAM[13][13] ),
    .CLK(clknet_leaf_103_clk_regs));
 sg13g2_dfrbpq_1 _09706_ (.RESET_B(net191),
    .D(_01106_),
    .Q(\rf_ram.RAM[13][14] ),
    .CLK(clknet_leaf_157_clk_regs));
 sg13g2_dfrbpq_1 _09707_ (.RESET_B(net190),
    .D(_01107_),
    .Q(\rf_ram.RAM[13][15] ),
    .CLK(clknet_leaf_148_clk_regs));
 sg13g2_dfrbpq_1 _09708_ (.RESET_B(net189),
    .D(_01108_),
    .Q(\rf_ram.RAM[13][16] ),
    .CLK(clknet_leaf_108_clk_regs));
 sg13g2_dfrbpq_1 _09709_ (.RESET_B(net188),
    .D(_01109_),
    .Q(\rf_ram.RAM[13][17] ),
    .CLK(clknet_leaf_140_clk_regs));
 sg13g2_dfrbpq_1 _09710_ (.RESET_B(net187),
    .D(_01110_),
    .Q(\rf_ram.RAM[13][18] ),
    .CLK(clknet_leaf_133_clk_regs));
 sg13g2_dfrbpq_1 _09711_ (.RESET_B(net186),
    .D(_01111_),
    .Q(\rf_ram.RAM[13][19] ),
    .CLK(clknet_leaf_155_clk_regs));
 sg13g2_dfrbpq_1 _09712_ (.RESET_B(net185),
    .D(_01112_),
    .Q(\rf_ram.RAM[13][20] ),
    .CLK(clknet_leaf_150_clk_regs));
 sg13g2_dfrbpq_1 _09713_ (.RESET_B(net184),
    .D(_01113_),
    .Q(\rf_ram.RAM[13][21] ),
    .CLK(clknet_leaf_55_clk_regs));
 sg13g2_dfrbpq_1 _09714_ (.RESET_B(net183),
    .D(_01114_),
    .Q(\rf_ram.RAM[13][22] ),
    .CLK(clknet_leaf_66_clk_regs));
 sg13g2_dfrbpq_1 _09715_ (.RESET_B(net182),
    .D(_01115_),
    .Q(\rf_ram.RAM[13][23] ),
    .CLK(clknet_leaf_23_clk_regs));
 sg13g2_dfrbpq_1 _09716_ (.RESET_B(net181),
    .D(_01116_),
    .Q(\rf_ram.RAM[13][24] ),
    .CLK(clknet_leaf_75_clk_regs));
 sg13g2_dfrbpq_1 _09717_ (.RESET_B(net180),
    .D(_01117_),
    .Q(\rf_ram.RAM[13][25] ),
    .CLK(clknet_leaf_54_clk_regs));
 sg13g2_dfrbpq_1 _09718_ (.RESET_B(net179),
    .D(_01118_),
    .Q(\rf_ram.RAM[13][26] ),
    .CLK(clknet_leaf_47_clk_regs));
 sg13g2_dfrbpq_1 _09719_ (.RESET_B(net178),
    .D(_01119_),
    .Q(\rf_ram.RAM[13][27] ),
    .CLK(clknet_leaf_44_clk_regs));
 sg13g2_dfrbpq_1 _09720_ (.RESET_B(net177),
    .D(_01120_),
    .Q(\rf_ram.RAM[13][28] ),
    .CLK(clknet_leaf_26_clk_regs));
 sg13g2_dfrbpq_1 _09721_ (.RESET_B(net176),
    .D(_01121_),
    .Q(\rf_ram.RAM[13][29] ),
    .CLK(clknet_leaf_5_clk_regs));
 sg13g2_dfrbpq_1 _09722_ (.RESET_B(net175),
    .D(_01122_),
    .Q(\rf_ram.RAM[13][30] ),
    .CLK(clknet_leaf_165_clk_regs));
 sg13g2_dfrbpq_1 _09723_ (.RESET_B(net174),
    .D(_01123_),
    .Q(\rf_ram.RAM[13][31] ),
    .CLK(clknet_leaf_166_clk_regs));
 sg13g2_dfrbpq_1 _09724_ (.RESET_B(net173),
    .D(net1631),
    .Q(\rf_ram.RAM[12][0] ),
    .CLK(clknet_leaf_17_clk_regs));
 sg13g2_dfrbpq_1 _09725_ (.RESET_B(net172),
    .D(_01125_),
    .Q(\rf_ram.RAM[12][1] ),
    .CLK(clknet_leaf_53_clk_regs));
 sg13g2_dfrbpq_1 _09726_ (.RESET_B(net171),
    .D(_01126_),
    .Q(\rf_ram.RAM[12][2] ),
    .CLK(clknet_leaf_77_clk_regs));
 sg13g2_dfrbpq_1 _09727_ (.RESET_B(net170),
    .D(_01127_),
    .Q(\rf_ram.RAM[12][3] ),
    .CLK(clknet_leaf_84_clk_regs));
 sg13g2_dfrbpq_1 _09728_ (.RESET_B(net169),
    .D(_01128_),
    .Q(\rf_ram.RAM[12][4] ),
    .CLK(clknet_leaf_77_clk_regs));
 sg13g2_dfrbpq_1 _09729_ (.RESET_B(net168),
    .D(_01129_),
    .Q(\rf_ram.RAM[12][5] ),
    .CLK(clknet_leaf_85_clk_regs));
 sg13g2_dfrbpq_1 _09730_ (.RESET_B(net167),
    .D(_01130_),
    .Q(\rf_ram.RAM[12][6] ),
    .CLK(clknet_leaf_94_clk_regs));
 sg13g2_dfrbpq_1 _09731_ (.RESET_B(net166),
    .D(_01131_),
    .Q(\rf_ram.RAM[12][7] ),
    .CLK(clknet_leaf_94_clk_regs));
 sg13g2_dfrbpq_1 _09732_ (.RESET_B(net165),
    .D(_01132_),
    .Q(\rf_ram.RAM[12][8] ),
    .CLK(clknet_leaf_115_clk_regs));
 sg13g2_dfrbpq_1 _09733_ (.RESET_B(net164),
    .D(_01133_),
    .Q(\rf_ram.RAM[12][9] ),
    .CLK(clknet_leaf_125_clk_regs));
 sg13g2_dfrbpq_1 _09734_ (.RESET_B(net163),
    .D(_01134_),
    .Q(\rf_ram.RAM[12][10] ),
    .CLK(clknet_leaf_120_clk_regs));
 sg13g2_dfrbpq_1 _09735_ (.RESET_B(net162),
    .D(_01135_),
    .Q(\rf_ram.RAM[12][11] ),
    .CLK(clknet_leaf_132_clk_regs));
 sg13g2_dfrbpq_1 _09736_ (.RESET_B(net161),
    .D(_01136_),
    .Q(\rf_ram.RAM[12][12] ),
    .CLK(clknet_leaf_118_clk_regs));
 sg13g2_dfrbpq_1 _09737_ (.RESET_B(net160),
    .D(_01137_),
    .Q(\rf_ram.RAM[12][13] ),
    .CLK(clknet_leaf_103_clk_regs));
 sg13g2_dfrbpq_1 _09738_ (.RESET_B(net159),
    .D(_01138_),
    .Q(\rf_ram.RAM[12][14] ),
    .CLK(clknet_leaf_157_clk_regs));
 sg13g2_dfrbpq_1 _09739_ (.RESET_B(net158),
    .D(_01139_),
    .Q(\rf_ram.RAM[12][15] ),
    .CLK(clknet_leaf_147_clk_regs));
 sg13g2_dfrbpq_1 _09740_ (.RESET_B(net157),
    .D(_01140_),
    .Q(\rf_ram.RAM[12][16] ),
    .CLK(clknet_leaf_108_clk_regs));
 sg13g2_dfrbpq_1 _09741_ (.RESET_B(net156),
    .D(_01141_),
    .Q(\rf_ram.RAM[12][17] ),
    .CLK(clknet_leaf_141_clk_regs));
 sg13g2_dfrbpq_1 _09742_ (.RESET_B(net155),
    .D(_01142_),
    .Q(\rf_ram.RAM[12][18] ),
    .CLK(clknet_leaf_132_clk_regs));
 sg13g2_dfrbpq_1 _09743_ (.RESET_B(net154),
    .D(_01143_),
    .Q(\rf_ram.RAM[12][19] ),
    .CLK(clknet_leaf_164_clk_regs));
 sg13g2_dfrbpq_1 _09744_ (.RESET_B(net153),
    .D(_01144_),
    .Q(\rf_ram.RAM[12][20] ),
    .CLK(clknet_leaf_150_clk_regs));
 sg13g2_dfrbpq_1 _09745_ (.RESET_B(net152),
    .D(_01145_),
    .Q(\rf_ram.RAM[12][21] ),
    .CLK(clknet_leaf_60_clk_regs));
 sg13g2_dfrbpq_1 _09746_ (.RESET_B(net151),
    .D(_01146_),
    .Q(\rf_ram.RAM[12][22] ),
    .CLK(clknet_leaf_104_clk_regs));
 sg13g2_dfrbpq_1 _09747_ (.RESET_B(net150),
    .D(_01147_),
    .Q(\rf_ram.RAM[12][23] ),
    .CLK(clknet_leaf_59_clk_regs));
 sg13g2_dfrbpq_1 _09748_ (.RESET_B(net149),
    .D(_01148_),
    .Q(\rf_ram.RAM[12][24] ),
    .CLK(clknet_leaf_75_clk_regs));
 sg13g2_dfrbpq_1 _09749_ (.RESET_B(net148),
    .D(_01149_),
    .Q(\rf_ram.RAM[12][25] ),
    .CLK(clknet_leaf_53_clk_regs));
 sg13g2_dfrbpq_1 _09750_ (.RESET_B(net147),
    .D(_01150_),
    .Q(\rf_ram.RAM[12][26] ),
    .CLK(clknet_leaf_47_clk_regs));
 sg13g2_dfrbpq_1 _09751_ (.RESET_B(net146),
    .D(_01151_),
    .Q(\rf_ram.RAM[12][27] ),
    .CLK(clknet_leaf_44_clk_regs));
 sg13g2_dfrbpq_1 _09752_ (.RESET_B(net145),
    .D(_01152_),
    .Q(\rf_ram.RAM[12][28] ),
    .CLK(clknet_leaf_58_clk_regs));
 sg13g2_dfrbpq_1 _09753_ (.RESET_B(net144),
    .D(_01153_),
    .Q(\rf_ram.RAM[12][29] ),
    .CLK(clknet_leaf_16_clk_regs));
 sg13g2_dfrbpq_1 _09754_ (.RESET_B(net143),
    .D(_01154_),
    .Q(\rf_ram.RAM[12][30] ),
    .CLK(clknet_leaf_165_clk_regs));
 sg13g2_dfrbpq_1 _09755_ (.RESET_B(net142),
    .D(_01155_),
    .Q(\rf_ram.RAM[12][31] ),
    .CLK(clknet_leaf_166_clk_regs));
 sg13g2_dfrbpq_1 _09756_ (.RESET_B(net141),
    .D(_01156_),
    .Q(\rf_ram.RAM[27][0] ),
    .CLK(clknet_leaf_17_clk_regs));
 sg13g2_dfrbpq_1 _09757_ (.RESET_B(net140),
    .D(_01157_),
    .Q(\rf_ram.RAM[27][1] ),
    .CLK(clknet_leaf_51_clk_regs));
 sg13g2_dfrbpq_1 _09758_ (.RESET_B(net139),
    .D(_01158_),
    .Q(\rf_ram.RAM[27][2] ),
    .CLK(clknet_leaf_78_clk_regs));
 sg13g2_dfrbpq_1 _09759_ (.RESET_B(net138),
    .D(_01159_),
    .Q(\rf_ram.RAM[27][3] ),
    .CLK(clknet_leaf_79_clk_regs));
 sg13g2_dfrbpq_1 _09760_ (.RESET_B(net137),
    .D(_01160_),
    .Q(\rf_ram.RAM[27][4] ),
    .CLK(clknet_leaf_86_clk_regs));
 sg13g2_dfrbpq_1 _09761_ (.RESET_B(net136),
    .D(_01161_),
    .Q(\rf_ram.RAM[27][5] ),
    .CLK(clknet_leaf_84_clk_regs));
 sg13g2_dfrbpq_1 _09762_ (.RESET_B(net135),
    .D(_01162_),
    .Q(\rf_ram.RAM[27][6] ),
    .CLK(clknet_leaf_91_clk_regs));
 sg13g2_dfrbpq_1 _09763_ (.RESET_B(net134),
    .D(_01163_),
    .Q(\rf_ram.RAM[27][7] ),
    .CLK(clknet_leaf_94_clk_regs));
 sg13g2_dfrbpq_1 _09764_ (.RESET_B(net133),
    .D(_01164_),
    .Q(\rf_ram.RAM[27][8] ),
    .CLK(clknet_leaf_113_clk_regs));
 sg13g2_dfrbpq_1 _09765_ (.RESET_B(net132),
    .D(_01165_),
    .Q(\rf_ram.RAM[27][9] ),
    .CLK(clknet_leaf_127_clk_regs));
 sg13g2_dfrbpq_1 _09766_ (.RESET_B(net131),
    .D(_01166_),
    .Q(\rf_ram.RAM[27][10] ),
    .CLK(clknet_leaf_125_clk_regs));
 sg13g2_dfrbpq_1 _09767_ (.RESET_B(net130),
    .D(_01167_),
    .Q(\rf_ram.RAM[27][11] ),
    .CLK(clknet_leaf_130_clk_regs));
 sg13g2_dfrbpq_1 _09768_ (.RESET_B(net129),
    .D(_01168_),
    .Q(\rf_ram.RAM[27][12] ),
    .CLK(clknet_leaf_125_clk_regs));
 sg13g2_dfrbpq_1 _09769_ (.RESET_B(net128),
    .D(_01169_),
    .Q(\rf_ram.RAM[27][13] ),
    .CLK(clknet_leaf_108_clk_regs));
 sg13g2_dfrbpq_1 _09770_ (.RESET_B(net127),
    .D(_01170_),
    .Q(\rf_ram.RAM[27][14] ),
    .CLK(clknet_leaf_158_clk_regs));
 sg13g2_dfrbpq_1 _09771_ (.RESET_B(net126),
    .D(_01171_),
    .Q(\rf_ram.RAM[27][15] ),
    .CLK(clknet_leaf_148_clk_regs));
 sg13g2_dfrbpq_1 _09772_ (.RESET_B(net125),
    .D(_01172_),
    .Q(\rf_ram.RAM[27][16] ),
    .CLK(clknet_leaf_108_clk_regs));
 sg13g2_dfrbpq_1 _09773_ (.RESET_B(net124),
    .D(_01173_),
    .Q(\rf_ram.RAM[27][17] ),
    .CLK(clknet_leaf_159_clk_regs));
 sg13g2_dfrbpq_1 _09774_ (.RESET_B(net123),
    .D(_01174_),
    .Q(\rf_ram.RAM[27][18] ),
    .CLK(clknet_leaf_142_clk_regs));
 sg13g2_dfrbpq_1 _09775_ (.RESET_B(net122),
    .D(_01175_),
    .Q(\rf_ram.RAM[27][19] ),
    .CLK(clknet_leaf_21_clk_regs));
 sg13g2_dfrbpq_1 _09776_ (.RESET_B(net121),
    .D(_01176_),
    .Q(\rf_ram.RAM[27][20] ),
    .CLK(clknet_leaf_150_clk_regs));
 sg13g2_dfrbpq_1 _09777_ (.RESET_B(net120),
    .D(_01177_),
    .Q(\rf_ram.RAM[27][21] ),
    .CLK(clknet_leaf_65_clk_regs));
 sg13g2_dfrbpq_1 _09778_ (.RESET_B(net119),
    .D(_01178_),
    .Q(\rf_ram.RAM[27][22] ),
    .CLK(clknet_leaf_70_clk_regs));
 sg13g2_dfrbpq_1 _09779_ (.RESET_B(net118),
    .D(_01179_),
    .Q(\rf_ram.RAM[27][23] ),
    .CLK(clknet_leaf_18_clk_regs));
 sg13g2_dfrbpq_1 _09780_ (.RESET_B(net117),
    .D(_01180_),
    .Q(\rf_ram.RAM[27][24] ),
    .CLK(clknet_leaf_72_clk_regs));
 sg13g2_dfrbpq_1 _09781_ (.RESET_B(net116),
    .D(_01181_),
    .Q(\rf_ram.RAM[27][25] ),
    .CLK(clknet_leaf_49_clk_regs));
 sg13g2_dfrbpq_1 _09782_ (.RESET_B(net115),
    .D(_01182_),
    .Q(\rf_ram.RAM[27][26] ),
    .CLK(clknet_leaf_71_clk_regs));
 sg13g2_dfrbpq_1 _09783_ (.RESET_B(net114),
    .D(_01183_),
    .Q(\rf_ram.RAM[27][27] ),
    .CLK(clknet_leaf_43_clk_regs));
 sg13g2_dfrbpq_1 _09784_ (.RESET_B(net113),
    .D(_01184_),
    .Q(\rf_ram.RAM[27][28] ),
    .CLK(clknet_leaf_34_clk_regs));
 sg13g2_dfrbpq_1 _09785_ (.RESET_B(net112),
    .D(_01185_),
    .Q(\rf_ram.RAM[27][29] ),
    .CLK(clknet_leaf_15_clk_regs));
 sg13g2_dfrbpq_1 _09786_ (.RESET_B(net111),
    .D(_01186_),
    .Q(\rf_ram.RAM[27][30] ),
    .CLK(clknet_leaf_164_clk_regs));
 sg13g2_dfrbpq_1 _09787_ (.RESET_B(net110),
    .D(_01187_),
    .Q(\rf_ram.RAM[27][31] ),
    .CLK(clknet_leaf_166_clk_regs));
 sg13g2_dfrbpq_1 _09788_ (.RESET_B(net109),
    .D(net3022),
    .Q(\rf_ram.RAM[11][0] ),
    .CLK(clknet_leaf_153_clk_regs));
 sg13g2_dfrbpq_1 _09789_ (.RESET_B(net108),
    .D(_01189_),
    .Q(\rf_ram.RAM[11][1] ),
    .CLK(clknet_leaf_55_clk_regs));
 sg13g2_dfrbpq_1 _09790_ (.RESET_B(net107),
    .D(_01190_),
    .Q(\rf_ram.RAM[11][2] ),
    .CLK(clknet_leaf_69_clk_regs));
 sg13g2_dfrbpq_1 _09791_ (.RESET_B(net106),
    .D(_01191_),
    .Q(\rf_ram.RAM[11][3] ),
    .CLK(clknet_leaf_79_clk_regs));
 sg13g2_dfrbpq_1 _09792_ (.RESET_B(net105),
    .D(_01192_),
    .Q(\rf_ram.RAM[11][4] ),
    .CLK(clknet_leaf_82_clk_regs));
 sg13g2_dfrbpq_1 _09793_ (.RESET_B(net104),
    .D(_01193_),
    .Q(\rf_ram.RAM[11][5] ),
    .CLK(clknet_leaf_80_clk_regs));
 sg13g2_dfrbpq_1 _09794_ (.RESET_B(net103),
    .D(_01194_),
    .Q(\rf_ram.RAM[11][6] ),
    .CLK(clknet_leaf_100_clk_regs));
 sg13g2_dfrbpq_1 _09795_ (.RESET_B(net102),
    .D(_01195_),
    .Q(\rf_ram.RAM[11][7] ),
    .CLK(clknet_leaf_99_clk_regs));
 sg13g2_dfrbpq_1 _09796_ (.RESET_B(net101),
    .D(_01196_),
    .Q(\rf_ram.RAM[11][8] ),
    .CLK(clknet_leaf_112_clk_regs));
 sg13g2_dfrbpq_1 _09797_ (.RESET_B(net100),
    .D(_01197_),
    .Q(\rf_ram.RAM[11][9] ),
    .CLK(clknet_leaf_131_clk_regs));
 sg13g2_dfrbpq_1 _09798_ (.RESET_B(net99),
    .D(_01198_),
    .Q(\rf_ram.RAM[11][10] ),
    .CLK(clknet_leaf_112_clk_regs));
 sg13g2_dfrbpq_1 _09799_ (.RESET_B(net98),
    .D(_01199_),
    .Q(\rf_ram.RAM[11][11] ),
    .CLK(clknet_leaf_129_clk_regs));
 sg13g2_dfrbpq_1 _09800_ (.RESET_B(net97),
    .D(_01200_),
    .Q(\rf_ram.RAM[11][12] ),
    .CLK(clknet_leaf_128_clk_regs));
 sg13g2_dfrbpq_1 _09801_ (.RESET_B(net96),
    .D(_01201_),
    .Q(\rf_ram.RAM[11][13] ),
    .CLK(clknet_leaf_103_clk_regs));
 sg13g2_dfrbpq_1 _09802_ (.RESET_B(net95),
    .D(_01202_),
    .Q(\rf_ram.RAM[11][14] ),
    .CLK(clknet_leaf_158_clk_regs));
 sg13g2_dfrbpq_1 _09803_ (.RESET_B(net94),
    .D(_01203_),
    .Q(\rf_ram.RAM[11][15] ),
    .CLK(clknet_leaf_107_clk_regs));
 sg13g2_dfrbpq_1 _09804_ (.RESET_B(net93),
    .D(_01204_),
    .Q(\rf_ram.RAM[11][16] ),
    .CLK(clknet_leaf_101_clk_regs));
 sg13g2_dfrbpq_1 _09805_ (.RESET_B(net92),
    .D(_01205_),
    .Q(\rf_ram.RAM[11][17] ),
    .CLK(clknet_leaf_139_clk_regs));
 sg13g2_dfrbpq_1 _09806_ (.RESET_B(net91),
    .D(_01206_),
    .Q(\rf_ram.RAM[11][18] ),
    .CLK(clknet_leaf_133_clk_regs));
 sg13g2_dfrbpq_1 _09807_ (.RESET_B(net90),
    .D(_01207_),
    .Q(\rf_ram.RAM[11][19] ),
    .CLK(clknet_leaf_158_clk_regs));
 sg13g2_dfrbpq_1 _09808_ (.RESET_B(net89),
    .D(_01208_),
    .Q(\rf_ram.RAM[11][20] ),
    .CLK(clknet_leaf_153_clk_regs));
 sg13g2_dfrbpq_1 _09809_ (.RESET_B(net88),
    .D(_01209_),
    .Q(\rf_ram.RAM[11][21] ),
    .CLK(clknet_leaf_62_clk_regs));
 sg13g2_dfrbpq_1 _09810_ (.RESET_B(net87),
    .D(_01210_),
    .Q(\rf_ram.RAM[11][22] ),
    .CLK(clknet_leaf_64_clk_regs));
 sg13g2_dfrbpq_1 _09811_ (.RESET_B(net86),
    .D(_01211_),
    .Q(\rf_ram.RAM[11][23] ),
    .CLK(clknet_leaf_18_clk_regs));
 sg13g2_dfrbpq_1 _09812_ (.RESET_B(net85),
    .D(_01212_),
    .Q(\rf_ram.RAM[11][24] ),
    .CLK(clknet_leaf_72_clk_regs));
 sg13g2_dfrbpq_1 _09813_ (.RESET_B(net84),
    .D(_01213_),
    .Q(\rf_ram.RAM[11][25] ),
    .CLK(clknet_leaf_57_clk_regs));
 sg13g2_dfrbpq_1 _09814_ (.RESET_B(net81),
    .D(_01214_),
    .Q(\rf_ram.RAM[11][26] ),
    .CLK(clknet_leaf_59_clk_regs));
 sg13g2_dfrbpq_1 _09815_ (.RESET_B(net80),
    .D(_01215_),
    .Q(\rf_ram.RAM[11][27] ),
    .CLK(clknet_leaf_46_clk_regs));
 sg13g2_dfrbpq_1 _09816_ (.RESET_B(net79),
    .D(_01216_),
    .Q(\rf_ram.RAM[11][28] ),
    .CLK(clknet_leaf_28_clk_regs));
 sg13g2_dfrbpq_1 _09817_ (.RESET_B(net78),
    .D(_01217_),
    .Q(\rf_ram.RAM[11][29] ),
    .CLK(clknet_leaf_166_clk_regs));
 sg13g2_dfrbpq_1 _09818_ (.RESET_B(net77),
    .D(_01218_),
    .Q(\rf_ram.RAM[11][30] ),
    .CLK(clknet_leaf_161_clk_regs));
 sg13g2_dfrbpq_1 _09819_ (.RESET_B(net76),
    .D(_01219_),
    .Q(\rf_ram.RAM[11][31] ),
    .CLK(clknet_leaf_168_clk_regs));
 sg13g2_dfrbpq_1 _09820_ (.RESET_B(net75),
    .D(net2840),
    .Q(\rf_ram.RAM[0][0] ),
    .CLK(clknet_leaf_14_clk_regs));
 sg13g2_dfrbpq_1 _09821_ (.RESET_B(net74),
    .D(_01221_),
    .Q(\rf_ram.RAM[0][1] ),
    .CLK(clknet_leaf_73_clk_regs));
 sg13g2_dfrbpq_1 _09822_ (.RESET_B(net73),
    .D(_01222_),
    .Q(\rf_ram.RAM[0][2] ),
    .CLK(clknet_leaf_78_clk_regs));
 sg13g2_dfrbpq_1 _09823_ (.RESET_B(net72),
    .D(_01223_),
    .Q(\rf_ram.RAM[0][3] ),
    .CLK(clknet_leaf_77_clk_regs));
 sg13g2_dfrbpq_1 _09824_ (.RESET_B(net71),
    .D(_01224_),
    .Q(\rf_ram.RAM[0][4] ),
    .CLK(clknet_leaf_82_clk_regs));
 sg13g2_dfrbpq_1 _09825_ (.RESET_B(net70),
    .D(_01225_),
    .Q(\rf_ram.RAM[0][5] ),
    .CLK(clknet_leaf_81_clk_regs));
 sg13g2_dfrbpq_1 _09826_ (.RESET_B(net69),
    .D(_01226_),
    .Q(\rf_ram.RAM[0][6] ),
    .CLK(clknet_leaf_101_clk_regs));
 sg13g2_dfrbpq_1 _09827_ (.RESET_B(net68),
    .D(_01227_),
    .Q(\rf_ram.RAM[0][7] ),
    .CLK(clknet_leaf_99_clk_regs));
 sg13g2_dfrbpq_1 _09828_ (.RESET_B(net67),
    .D(_01228_),
    .Q(\rf_ram.RAM[0][8] ),
    .CLK(clknet_leaf_112_clk_regs));
 sg13g2_dfrbpq_1 _09829_ (.RESET_B(net66),
    .D(_01229_),
    .Q(\rf_ram.RAM[0][9] ),
    .CLK(clknet_leaf_127_clk_regs));
 sg13g2_dfrbpq_1 _09830_ (.RESET_B(net65),
    .D(_01230_),
    .Q(\rf_ram.RAM[0][10] ),
    .CLK(clknet_leaf_120_clk_regs));
 sg13g2_dfrbpq_1 _09831_ (.RESET_B(net64),
    .D(_01231_),
    .Q(\rf_ram.RAM[0][11] ),
    .CLK(clknet_leaf_129_clk_regs));
 sg13g2_dfrbpq_1 _09832_ (.RESET_B(net63),
    .D(_01232_),
    .Q(\rf_ram.RAM[0][12] ),
    .CLK(clknet_leaf_128_clk_regs));
 sg13g2_dfrbpq_1 _09833_ (.RESET_B(net62),
    .D(_01233_),
    .Q(\rf_ram.RAM[0][13] ),
    .CLK(clknet_leaf_110_clk_regs));
 sg13g2_dfrbpq_1 _09834_ (.RESET_B(net61),
    .D(_01234_),
    .Q(\rf_ram.RAM[0][14] ),
    .CLK(clknet_leaf_161_clk_regs));
 sg13g2_dfrbpq_1 _09835_ (.RESET_B(net60),
    .D(_01235_),
    .Q(\rf_ram.RAM[0][15] ),
    .CLK(clknet_leaf_147_clk_regs));
 sg13g2_dfrbpq_1 _09836_ (.RESET_B(net59),
    .D(_01236_),
    .Q(\rf_ram.RAM[0][16] ),
    .CLK(clknet_leaf_101_clk_regs));
 sg13g2_dfrbpq_1 _09837_ (.RESET_B(net58),
    .D(_01237_),
    .Q(\rf_ram.RAM[0][17] ),
    .CLK(clknet_leaf_139_clk_regs));
 sg13g2_dfrbpq_1 _09838_ (.RESET_B(net57),
    .D(_01238_),
    .Q(\rf_ram.RAM[0][18] ),
    .CLK(clknet_leaf_137_clk_regs));
 sg13g2_dfrbpq_1 _09839_ (.RESET_B(net56),
    .D(_01239_),
    .Q(\rf_ram.RAM[0][19] ),
    .CLK(clknet_leaf_152_clk_regs));
 sg13g2_dfrbpq_1 _09840_ (.RESET_B(net55),
    .D(_01240_),
    .Q(\rf_ram.RAM[0][20] ),
    .CLK(clknet_leaf_153_clk_regs));
 sg13g2_dfrbpq_1 _09841_ (.RESET_B(net54),
    .D(_01241_),
    .Q(\rf_ram.RAM[0][21] ),
    .CLK(clknet_leaf_22_clk_regs));
 sg13g2_dfrbpq_1 _09842_ (.RESET_B(net53),
    .D(_01242_),
    .Q(\rf_ram.RAM[0][22] ),
    .CLK(clknet_leaf_64_clk_regs));
 sg13g2_dfrbpq_1 _09843_ (.RESET_B(net52),
    .D(_01243_),
    .Q(\rf_ram.RAM[0][23] ),
    .CLK(clknet_leaf_19_clk_regs));
 sg13g2_dfrbpq_1 _09844_ (.RESET_B(net51),
    .D(_01244_),
    .Q(\rf_ram.RAM[0][24] ),
    .CLK(clknet_leaf_74_clk_regs));
 sg13g2_dfrbpq_1 _09845_ (.RESET_B(net50),
    .D(_01245_),
    .Q(\rf_ram.RAM[0][25] ),
    .CLK(clknet_leaf_47_clk_regs));
 sg13g2_dfrbpq_1 _09846_ (.RESET_B(net49),
    .D(_01246_),
    .Q(\rf_ram.RAM[0][26] ),
    .CLK(clknet_leaf_50_clk_regs));
 sg13g2_dfrbpq_1 _09847_ (.RESET_B(net48),
    .D(_01247_),
    .Q(\rf_ram.RAM[0][27] ),
    .CLK(clknet_leaf_45_clk_regs));
 sg13g2_dfrbpq_1 _09848_ (.RESET_B(net47),
    .D(_01248_),
    .Q(\rf_ram.RAM[0][28] ),
    .CLK(clknet_leaf_27_clk_regs));
 sg13g2_dfrbpq_1 _09849_ (.RESET_B(net46),
    .D(_01249_),
    .Q(\rf_ram.RAM[0][29] ),
    .CLK(clknet_leaf_167_clk_regs));
 sg13g2_dfrbpq_1 _09850_ (.RESET_B(net45),
    .D(_01250_),
    .Q(\rf_ram.RAM[0][30] ),
    .CLK(clknet_leaf_165_clk_regs));
 sg13g2_dfrbpq_1 _09851_ (.RESET_B(net44),
    .D(_01251_),
    .Q(\rf_ram.RAM[0][31] ),
    .CLK(clknet_leaf_4_clk_regs));
 sg13g2_dfrbpq_1 _09852_ (.RESET_B(net43),
    .D(_01252_),
    .Q(\rf_ram.RAM[19][0] ),
    .CLK(clknet_leaf_19_clk_regs));
 sg13g2_dfrbpq_1 _09853_ (.RESET_B(net42),
    .D(_01253_),
    .Q(\rf_ram.RAM[19][1] ),
    .CLK(clknet_leaf_54_clk_regs));
 sg13g2_dfrbpq_1 _09854_ (.RESET_B(net41),
    .D(_01254_),
    .Q(\rf_ram.RAM[19][2] ),
    .CLK(clknet_leaf_69_clk_regs));
 sg13g2_dfrbpq_1 _09855_ (.RESET_B(net40),
    .D(_01255_),
    .Q(\rf_ram.RAM[19][3] ),
    .CLK(clknet_leaf_88_clk_regs));
 sg13g2_dfrbpq_1 _09856_ (.RESET_B(net39),
    .D(_01256_),
    .Q(\rf_ram.RAM[19][4] ),
    .CLK(clknet_leaf_87_clk_regs));
 sg13g2_dfrbpq_1 _09857_ (.RESET_B(net38),
    .D(_01257_),
    .Q(\rf_ram.RAM[19][5] ),
    .CLK(clknet_leaf_93_clk_regs));
 sg13g2_dfrbpq_1 _09858_ (.RESET_B(net37),
    .D(_01258_),
    .Q(\rf_ram.RAM[19][6] ),
    .CLK(clknet_leaf_92_clk_regs));
 sg13g2_dfrbpq_1 _09859_ (.RESET_B(net36),
    .D(_01259_),
    .Q(\rf_ram.RAM[19][7] ),
    .CLK(clknet_leaf_95_clk_regs));
 sg13g2_dfrbpq_1 _09860_ (.RESET_B(net35),
    .D(_01260_),
    .Q(\rf_ram.RAM[19][8] ),
    .CLK(clknet_leaf_116_clk_regs));
 sg13g2_dfrbpq_1 _09861_ (.RESET_B(net34),
    .D(_01261_),
    .Q(\rf_ram.RAM[19][9] ),
    .CLK(clknet_leaf_126_clk_regs));
 sg13g2_dfrbpq_1 _09862_ (.RESET_B(net33),
    .D(_01262_),
    .Q(\rf_ram.RAM[19][10] ),
    .CLK(clknet_leaf_117_clk_regs));
 sg13g2_dfrbpq_1 _09863_ (.RESET_B(net32),
    .D(_01263_),
    .Q(\rf_ram.RAM[19][11] ),
    .CLK(clknet_leaf_135_clk_regs));
 sg13g2_dfrbpq_1 _09864_ (.RESET_B(net31),
    .D(_01264_),
    .Q(\rf_ram.RAM[19][12] ),
    .CLK(clknet_leaf_126_clk_regs));
 sg13g2_dfrbpq_1 _09865_ (.RESET_B(net30),
    .D(_01265_),
    .Q(\rf_ram.RAM[19][13] ),
    .CLK(clknet_leaf_143_clk_regs));
 sg13g2_dfrbpq_1 _09866_ (.RESET_B(net29),
    .D(_01266_),
    .Q(\rf_ram.RAM[19][14] ),
    .CLK(clknet_leaf_160_clk_regs));
 sg13g2_dfrbpq_1 _09867_ (.RESET_B(net28),
    .D(_01267_),
    .Q(\rf_ram.RAM[19][15] ),
    .CLK(clknet_leaf_144_clk_regs));
 sg13g2_dfrbpq_1 _09868_ (.RESET_B(net27),
    .D(_01268_),
    .Q(\rf_ram.RAM[19][16] ),
    .CLK(clknet_leaf_103_clk_regs));
 sg13g2_dfrbpq_1 _09869_ (.RESET_B(net26),
    .D(_01269_),
    .Q(\rf_ram.RAM[19][17] ),
    .CLK(clknet_leaf_138_clk_regs));
 sg13g2_dfrbpq_1 _09870_ (.RESET_B(net25),
    .D(_01270_),
    .Q(\rf_ram.RAM[19][18] ),
    .CLK(clknet_leaf_136_clk_regs));
 sg13g2_dfrbpq_1 _09871_ (.RESET_B(net24),
    .D(_01271_),
    .Q(\rf_ram.RAM[19][19] ),
    .CLK(clknet_leaf_160_clk_regs));
 sg13g2_dfrbpq_1 _09872_ (.RESET_B(net23),
    .D(_01272_),
    .Q(\rf_ram.RAM[19][20] ),
    .CLK(clknet_leaf_147_clk_regs));
 sg13g2_dfrbpq_1 _09873_ (.RESET_B(net22),
    .D(_01273_),
    .Q(\rf_ram.RAM[19][21] ),
    .CLK(clknet_leaf_61_clk_regs));
 sg13g2_dfrbpq_1 _09874_ (.RESET_B(net21),
    .D(_01274_),
    .Q(\rf_ram.RAM[19][22] ),
    .CLK(clknet_leaf_102_clk_regs));
 sg13g2_dfrbpq_1 _09875_ (.RESET_B(net20),
    .D(_01275_),
    .Q(\rf_ram.RAM[19][23] ),
    .CLK(clknet_leaf_22_clk_regs));
 sg13g2_dfrbpq_1 _09876_ (.RESET_B(net19),
    .D(_01276_),
    .Q(\rf_ram.RAM[19][24] ),
    .CLK(clknet_leaf_73_clk_regs));
 sg13g2_dfrbpq_1 _09877_ (.RESET_B(net18),
    .D(_01277_),
    .Q(\rf_ram.RAM[19][25] ),
    .CLK(clknet_leaf_50_clk_regs));
 sg13g2_dfrbpq_1 _09878_ (.RESET_B(net1373),
    .D(_01278_),
    .Q(\rf_ram.RAM[19][26] ),
    .CLK(clknet_leaf_58_clk_regs));
 sg13g2_dfrbpq_1 _09879_ (.RESET_B(net1372),
    .D(_01279_),
    .Q(\rf_ram.RAM[19][27] ),
    .CLK(clknet_leaf_48_clk_regs));
 sg13g2_dfrbpq_1 _09880_ (.RESET_B(net1371),
    .D(_01280_),
    .Q(\rf_ram.RAM[19][28] ),
    .CLK(clknet_leaf_25_clk_regs));
 sg13g2_dfrbpq_1 _09881_ (.RESET_B(net1370),
    .D(_01281_),
    .Q(\rf_ram.RAM[19][29] ),
    .CLK(clknet_leaf_170_clk_regs));
 sg13g2_dfrbpq_1 _09882_ (.RESET_B(net1369),
    .D(_01282_),
    .Q(\rf_ram.RAM[19][30] ),
    .CLK(clknet_leaf_163_clk_regs));
 sg13g2_dfrbpq_1 _09883_ (.RESET_B(net1368),
    .D(_01283_),
    .Q(\rf_ram.RAM[19][31] ),
    .CLK(clknet_leaf_169_clk_regs));
 sg13g2_dfrbpq_1 _09884_ (.RESET_B(net1366),
    .D(net2830),
    .Q(\rf_ram.RAM[8][0] ),
    .CLK(clknet_leaf_153_clk_regs));
 sg13g2_dfrbpq_1 _09885_ (.RESET_B(net1365),
    .D(_01285_),
    .Q(\rf_ram.RAM[8][1] ),
    .CLK(clknet_leaf_55_clk_regs));
 sg13g2_dfrbpq_1 _09886_ (.RESET_B(net1364),
    .D(_01286_),
    .Q(\rf_ram.RAM[8][2] ),
    .CLK(clknet_leaf_69_clk_regs));
 sg13g2_dfrbpq_1 _09887_ (.RESET_B(net1363),
    .D(_01287_),
    .Q(\rf_ram.RAM[8][3] ),
    .CLK(clknet_leaf_79_clk_regs));
 sg13g2_dfrbpq_1 _09888_ (.RESET_B(net1362),
    .D(_01288_),
    .Q(\rf_ram.RAM[8][4] ),
    .CLK(clknet_leaf_80_clk_regs));
 sg13g2_dfrbpq_1 _09889_ (.RESET_B(net1361),
    .D(_01289_),
    .Q(\rf_ram.RAM[8][5] ),
    .CLK(clknet_leaf_80_clk_regs));
 sg13g2_dfrbpq_1 _09890_ (.RESET_B(net1360),
    .D(_01290_),
    .Q(\rf_ram.RAM[8][6] ),
    .CLK(clknet_leaf_101_clk_regs));
 sg13g2_dfrbpq_1 _09891_ (.RESET_B(net1359),
    .D(_01291_),
    .Q(\rf_ram.RAM[8][7] ),
    .CLK(clknet_leaf_99_clk_regs));
 sg13g2_dfrbpq_1 _09892_ (.RESET_B(net1358),
    .D(_01292_),
    .Q(\rf_ram.RAM[8][8] ),
    .CLK(clknet_leaf_112_clk_regs));
 sg13g2_dfrbpq_1 _09893_ (.RESET_B(net1357),
    .D(_01293_),
    .Q(\rf_ram.RAM[8][9] ),
    .CLK(clknet_leaf_130_clk_regs));
 sg13g2_dfrbpq_1 _09894_ (.RESET_B(net1356),
    .D(_01294_),
    .Q(\rf_ram.RAM[8][10] ),
    .CLK(clknet_leaf_113_clk_regs));
 sg13g2_dfrbpq_1 _09895_ (.RESET_B(net1355),
    .D(_01295_),
    .Q(\rf_ram.RAM[8][11] ),
    .CLK(clknet_leaf_129_clk_regs));
 sg13g2_dfrbpq_1 _09896_ (.RESET_B(net1354),
    .D(_01296_),
    .Q(\rf_ram.RAM[8][12] ),
    .CLK(clknet_leaf_128_clk_regs));
 sg13g2_dfrbpq_1 _09897_ (.RESET_B(net1353),
    .D(_01297_),
    .Q(\rf_ram.RAM[8][13] ),
    .CLK(clknet_leaf_103_clk_regs));
 sg13g2_dfrbpq_1 _09898_ (.RESET_B(net1352),
    .D(_01298_),
    .Q(\rf_ram.RAM[8][14] ),
    .CLK(clknet_leaf_156_clk_regs));
 sg13g2_dfrbpq_1 _09899_ (.RESET_B(net1351),
    .D(_01299_),
    .Q(\rf_ram.RAM[8][15] ),
    .CLK(clknet_leaf_107_clk_regs));
 sg13g2_dfrbpq_1 _09900_ (.RESET_B(net1350),
    .D(_01300_),
    .Q(\rf_ram.RAM[8][16] ),
    .CLK(clknet_leaf_68_clk_regs));
 sg13g2_dfrbpq_1 _09901_ (.RESET_B(net1349),
    .D(_01301_),
    .Q(\rf_ram.RAM[8][17] ),
    .CLK(clknet_leaf_139_clk_regs));
 sg13g2_dfrbpq_1 _09902_ (.RESET_B(net1348),
    .D(_01302_),
    .Q(\rf_ram.RAM[8][18] ),
    .CLK(clknet_leaf_133_clk_regs));
 sg13g2_dfrbpq_1 _09903_ (.RESET_B(net1347),
    .D(_01303_),
    .Q(\rf_ram.RAM[8][19] ),
    .CLK(clknet_leaf_155_clk_regs));
 sg13g2_dfrbpq_1 _09904_ (.RESET_B(net1346),
    .D(_01304_),
    .Q(\rf_ram.RAM[8][20] ),
    .CLK(clknet_leaf_152_clk_regs));
 sg13g2_dfrbpq_1 _09905_ (.RESET_B(net1345),
    .D(_01305_),
    .Q(\rf_ram.RAM[8][21] ),
    .CLK(clknet_leaf_61_clk_regs));
 sg13g2_dfrbpq_1 _09906_ (.RESET_B(net1344),
    .D(_01306_),
    .Q(\rf_ram.RAM[8][22] ),
    .CLK(clknet_leaf_63_clk_regs));
 sg13g2_dfrbpq_1 _09907_ (.RESET_B(net1343),
    .D(_01307_),
    .Q(\rf_ram.RAM[8][23] ),
    .CLK(clknet_leaf_18_clk_regs));
 sg13g2_dfrbpq_1 _09908_ (.RESET_B(net1342),
    .D(_01308_),
    .Q(\rf_ram.RAM[8][24] ),
    .CLK(clknet_leaf_71_clk_regs));
 sg13g2_dfrbpq_1 _09909_ (.RESET_B(net1341),
    .D(_01309_),
    .Q(\rf_ram.RAM[8][25] ),
    .CLK(clknet_leaf_57_clk_regs));
 sg13g2_dfrbpq_1 _09910_ (.RESET_B(net1340),
    .D(_01310_),
    .Q(\rf_ram.RAM[8][26] ),
    .CLK(clknet_leaf_59_clk_regs));
 sg13g2_dfrbpq_1 _09911_ (.RESET_B(net1339),
    .D(_01311_),
    .Q(\rf_ram.RAM[8][27] ),
    .CLK(clknet_leaf_35_clk_regs));
 sg13g2_dfrbpq_1 _09912_ (.RESET_B(net1338),
    .D(_01312_),
    .Q(\rf_ram.RAM[8][28] ),
    .CLK(clknet_leaf_28_clk_regs));
 sg13g2_dfrbpq_1 _09913_ (.RESET_B(net1337),
    .D(_01313_),
    .Q(\rf_ram.RAM[8][29] ),
    .CLK(clknet_leaf_166_clk_regs));
 sg13g2_dfrbpq_1 _09914_ (.RESET_B(net1336),
    .D(_01314_),
    .Q(\rf_ram.RAM[8][30] ),
    .CLK(clknet_leaf_162_clk_regs));
 sg13g2_dfrbpq_1 _09915_ (.RESET_B(net1335),
    .D(_01315_),
    .Q(\rf_ram.RAM[8][31] ),
    .CLK(clknet_leaf_168_clk_regs));
 sg13g2_dfrbpq_1 _09916_ (.RESET_B(net1332),
    .D(_01316_),
    .Q(\rf_ram.RAM[16][0] ),
    .CLK(clknet_leaf_23_clk_regs));
 sg13g2_dfrbpq_1 _09917_ (.RESET_B(net1331),
    .D(_01317_),
    .Q(\rf_ram.RAM[16][1] ),
    .CLK(clknet_leaf_53_clk_regs));
 sg13g2_dfrbpq_1 _09918_ (.RESET_B(net1330),
    .D(_01318_),
    .Q(\rf_ram.RAM[16][2] ),
    .CLK(clknet_leaf_69_clk_regs));
 sg13g2_dfrbpq_1 _09919_ (.RESET_B(net1329),
    .D(_01319_),
    .Q(\rf_ram.RAM[16][3] ),
    .CLK(clknet_leaf_89_clk_regs));
 sg13g2_dfrbpq_1 _09920_ (.RESET_B(net1328),
    .D(_01320_),
    .Q(\rf_ram.RAM[16][4] ),
    .CLK(clknet_leaf_87_clk_regs));
 sg13g2_dfrbpq_1 _09921_ (.RESET_B(net1327),
    .D(_01321_),
    .Q(\rf_ram.RAM[16][5] ),
    .CLK(clknet_leaf_93_clk_regs));
 sg13g2_dfrbpq_1 _09922_ (.RESET_B(net1326),
    .D(_01322_),
    .Q(\rf_ram.RAM[16][6] ),
    .CLK(clknet_leaf_92_clk_regs));
 sg13g2_dfrbpq_1 _09923_ (.RESET_B(net1325),
    .D(_01323_),
    .Q(\rf_ram.RAM[16][7] ),
    .CLK(clknet_leaf_95_clk_regs));
 sg13g2_dfrbpq_1 _09924_ (.RESET_B(net1324),
    .D(_01324_),
    .Q(\rf_ram.RAM[16][8] ),
    .CLK(clknet_leaf_116_clk_regs));
 sg13g2_dfrbpq_1 _09925_ (.RESET_B(net1323),
    .D(_01325_),
    .Q(\rf_ram.RAM[16][9] ),
    .CLK(clknet_leaf_124_clk_regs));
 sg13g2_dfrbpq_1 _09926_ (.RESET_B(net1322),
    .D(_01326_),
    .Q(\rf_ram.RAM[16][10] ),
    .CLK(clknet_leaf_117_clk_regs));
 sg13g2_dfrbpq_1 _09927_ (.RESET_B(net1321),
    .D(_01327_),
    .Q(\rf_ram.RAM[16][11] ),
    .CLK(clknet_leaf_135_clk_regs));
 sg13g2_dfrbpq_1 _09928_ (.RESET_B(net1320),
    .D(_01328_),
    .Q(\rf_ram.RAM[16][12] ),
    .CLK(clknet_leaf_126_clk_regs));
 sg13g2_dfrbpq_1 _09929_ (.RESET_B(net1319),
    .D(_01329_),
    .Q(\rf_ram.RAM[16][13] ),
    .CLK(clknet_leaf_143_clk_regs));
 sg13g2_dfrbpq_1 _09930_ (.RESET_B(net1318),
    .D(_01330_),
    .Q(\rf_ram.RAM[16][14] ),
    .CLK(clknet_leaf_160_clk_regs));
 sg13g2_dfrbpq_1 _09931_ (.RESET_B(net1317),
    .D(_01331_),
    .Q(\rf_ram.RAM[16][15] ),
    .CLK(clknet_leaf_144_clk_regs));
 sg13g2_dfrbpq_1 _09932_ (.RESET_B(net1316),
    .D(_01332_),
    .Q(\rf_ram.RAM[16][16] ),
    .CLK(clknet_leaf_102_clk_regs));
 sg13g2_dfrbpq_1 _09933_ (.RESET_B(net1315),
    .D(_00072_),
    .Q(\rf_ram.RAM[16][17] ),
    .CLK(clknet_leaf_138_clk_regs));
 sg13g2_dfrbpq_1 _09934_ (.RESET_B(net1314),
    .D(_00073_),
    .Q(\rf_ram.RAM[16][18] ),
    .CLK(clknet_leaf_136_clk_regs));
 sg13g2_dfrbpq_1 _09935_ (.RESET_B(net1313),
    .D(_00074_),
    .Q(\rf_ram.RAM[16][19] ),
    .CLK(clknet_leaf_160_clk_regs));
 sg13g2_dfrbpq_1 _09936_ (.RESET_B(net1312),
    .D(_00075_),
    .Q(\rf_ram.RAM[16][20] ),
    .CLK(clknet_leaf_151_clk_regs));
 sg13g2_dfrbpq_1 _09937_ (.RESET_B(net1311),
    .D(_00076_),
    .Q(\rf_ram.RAM[16][21] ),
    .CLK(clknet_leaf_62_clk_regs));
 sg13g2_dfrbpq_1 _09938_ (.RESET_B(net1310),
    .D(_00077_),
    .Q(\rf_ram.RAM[16][22] ),
    .CLK(clknet_leaf_104_clk_regs));
 sg13g2_dfrbpq_1 _09939_ (.RESET_B(net1309),
    .D(_00078_),
    .Q(\rf_ram.RAM[16][23] ),
    .CLK(clknet_leaf_22_clk_regs));
 sg13g2_dfrbpq_1 _09940_ (.RESET_B(net1308),
    .D(_00079_),
    .Q(\rf_ram.RAM[16][24] ),
    .CLK(clknet_leaf_72_clk_regs));
 sg13g2_dfrbpq_1 _09941_ (.RESET_B(net1307),
    .D(_00080_),
    .Q(\rf_ram.RAM[16][25] ),
    .CLK(clknet_leaf_49_clk_regs));
 sg13g2_dfrbpq_1 _09942_ (.RESET_B(net1306),
    .D(_00081_),
    .Q(\rf_ram.RAM[16][26] ),
    .CLK(clknet_leaf_57_clk_regs));
 sg13g2_dfrbpq_1 _09943_ (.RESET_B(net1305),
    .D(_00082_),
    .Q(\rf_ram.RAM[16][27] ),
    .CLK(clknet_leaf_48_clk_regs));
 sg13g2_dfrbpq_1 _09944_ (.RESET_B(net1304),
    .D(_00083_),
    .Q(\rf_ram.RAM[16][28] ),
    .CLK(clknet_leaf_25_clk_regs));
 sg13g2_dfrbpq_1 _09945_ (.RESET_B(net1303),
    .D(_00084_),
    .Q(\rf_ram.RAM[16][29] ),
    .CLK(clknet_leaf_170_clk_regs));
 sg13g2_dfrbpq_1 _09946_ (.RESET_B(net1302),
    .D(_00085_),
    .Q(\rf_ram.RAM[16][30] ),
    .CLK(clknet_leaf_163_clk_regs));
 sg13g2_dfrbpq_1 _09947_ (.RESET_B(net1301),
    .D(_00086_),
    .Q(\rf_ram.RAM[16][31] ),
    .CLK(clknet_leaf_169_clk_regs));
 sg13g2_dfrbpq_1 _09948_ (.RESET_B(net1300),
    .D(_00087_),
    .Q(\rf_ram.RAM[17][0] ),
    .CLK(clknet_leaf_19_clk_regs));
 sg13g2_dfrbpq_1 _09949_ (.RESET_B(net1299),
    .D(_00088_),
    .Q(\rf_ram.RAM[17][1] ),
    .CLK(clknet_leaf_56_clk_regs));
 sg13g2_dfrbpq_1 _09950_ (.RESET_B(net1298),
    .D(_00089_),
    .Q(\rf_ram.RAM[17][2] ),
    .CLK(clknet_leaf_68_clk_regs));
 sg13g2_dfrbpq_1 _09951_ (.RESET_B(net1297),
    .D(_00090_),
    .Q(\rf_ram.RAM[17][3] ),
    .CLK(clknet_leaf_87_clk_regs));
 sg13g2_dfrbpq_1 _09952_ (.RESET_B(net1296),
    .D(_00091_),
    .Q(\rf_ram.RAM[17][4] ),
    .CLK(clknet_leaf_87_clk_regs));
 sg13g2_dfrbpq_1 _09953_ (.RESET_B(net1295),
    .D(_00092_),
    .Q(\rf_ram.RAM[17][5] ),
    .CLK(clknet_leaf_88_clk_regs));
 sg13g2_dfrbpq_1 _09954_ (.RESET_B(net1294),
    .D(_00093_),
    .Q(\rf_ram.RAM[17][6] ),
    .CLK(clknet_leaf_93_clk_regs));
 sg13g2_dfrbpq_1 _09955_ (.RESET_B(net1293),
    .D(_00094_),
    .Q(\rf_ram.RAM[17][7] ),
    .CLK(clknet_leaf_95_clk_regs));
 sg13g2_dfrbpq_1 _09956_ (.RESET_B(net1292),
    .D(_00095_),
    .Q(\rf_ram.RAM[17][8] ),
    .CLK(clknet_leaf_115_clk_regs));
 sg13g2_dfrbpq_1 _09957_ (.RESET_B(net1291),
    .D(_00096_),
    .Q(\rf_ram.RAM[17][9] ),
    .CLK(clknet_leaf_126_clk_regs));
 sg13g2_dfrbpq_1 _09958_ (.RESET_B(net1289),
    .D(_00097_),
    .Q(\rf_ram.RAM[17][10] ),
    .CLK(clknet_leaf_118_clk_regs));
 sg13g2_dfrbpq_1 _09959_ (.RESET_B(net1288),
    .D(_00098_),
    .Q(\rf_ram.RAM[17][11] ),
    .CLK(clknet_leaf_135_clk_regs));
 sg13g2_dfrbpq_1 _09960_ (.RESET_B(net1287),
    .D(_00099_),
    .Q(\rf_ram.RAM[17][12] ),
    .CLK(clknet_leaf_125_clk_regs));
 sg13g2_dfrbpq_1 _09961_ (.RESET_B(net1286),
    .D(_00100_),
    .Q(\rf_ram.RAM[17][13] ),
    .CLK(clknet_leaf_144_clk_regs));
 sg13g2_dfrbpq_1 _09962_ (.RESET_B(net1285),
    .D(_00101_),
    .Q(\rf_ram.RAM[17][14] ),
    .CLK(clknet_leaf_160_clk_regs));
 sg13g2_dfrbpq_1 _09963_ (.RESET_B(net1284),
    .D(_00102_),
    .Q(\rf_ram.RAM[17][15] ),
    .CLK(clknet_leaf_144_clk_regs));
 sg13g2_dfrbpq_1 _09964_ (.RESET_B(net1283),
    .D(_00103_),
    .Q(\rf_ram.RAM[17][16] ),
    .CLK(clknet_leaf_104_clk_regs));
 sg13g2_dfrbpq_1 _09965_ (.RESET_B(net1282),
    .D(_00104_),
    .Q(\rf_ram.RAM[17][17] ),
    .CLK(clknet_leaf_138_clk_regs));
 sg13g2_dfrbpq_1 _09966_ (.RESET_B(net1281),
    .D(_00105_),
    .Q(\rf_ram.RAM[17][18] ),
    .CLK(clknet_leaf_137_clk_regs));
 sg13g2_dfrbpq_1 _09967_ (.RESET_B(net1280),
    .D(_00106_),
    .Q(\rf_ram.RAM[17][19] ),
    .CLK(clknet_leaf_160_clk_regs));
 sg13g2_dfrbpq_1 _09968_ (.RESET_B(net1279),
    .D(_00107_),
    .Q(\rf_ram.RAM[17][20] ),
    .CLK(clknet_leaf_149_clk_regs));
 sg13g2_dfrbpq_1 _09969_ (.RESET_B(net1278),
    .D(_00108_),
    .Q(\rf_ram.RAM[17][21] ),
    .CLK(clknet_leaf_62_clk_regs));
 sg13g2_dfrbpq_1 _09970_ (.RESET_B(net1277),
    .D(_00109_),
    .Q(\rf_ram.RAM[17][22] ),
    .CLK(clknet_leaf_104_clk_regs));
 sg13g2_dfrbpq_1 _09971_ (.RESET_B(net1276),
    .D(_00110_),
    .Q(\rf_ram.RAM[17][23] ),
    .CLK(clknet_leaf_22_clk_regs));
 sg13g2_dfrbpq_1 _09972_ (.RESET_B(net1275),
    .D(_00111_),
    .Q(\rf_ram.RAM[17][24] ),
    .CLK(clknet_leaf_71_clk_regs));
 sg13g2_dfrbpq_1 _09973_ (.RESET_B(net1274),
    .D(_00112_),
    .Q(\rf_ram.RAM[17][25] ),
    .CLK(clknet_leaf_56_clk_regs));
 sg13g2_dfrbpq_1 _09974_ (.RESET_B(net1273),
    .D(_00113_),
    .Q(\rf_ram.RAM[17][26] ),
    .CLK(clknet_leaf_56_clk_regs));
 sg13g2_dfrbpq_1 _09975_ (.RESET_B(net1272),
    .D(_00114_),
    .Q(\rf_ram.RAM[17][27] ),
    .CLK(clknet_leaf_45_clk_regs));
 sg13g2_dfrbpq_1 _09976_ (.RESET_B(net1271),
    .D(_00115_),
    .Q(\rf_ram.RAM[17][28] ),
    .CLK(clknet_leaf_28_clk_regs));
 sg13g2_dfrbpq_1 _09977_ (.RESET_B(net1270),
    .D(_00116_),
    .Q(\rf_ram.RAM[17][29] ),
    .CLK(clknet_leaf_170_clk_regs));
 sg13g2_dfrbpq_1 _09978_ (.RESET_B(net1269),
    .D(_00117_),
    .Q(\rf_ram.RAM[17][30] ),
    .CLK(clknet_leaf_162_clk_regs));
 sg13g2_dfrbpq_1 _09979_ (.RESET_B(net1268),
    .D(_00118_),
    .Q(\rf_ram.RAM[17][31] ),
    .CLK(clknet_leaf_170_clk_regs));
 sg13g2_dfrbpq_1 _09980_ (.RESET_B(net1267),
    .D(_00119_),
    .Q(\rf_ram.RAM[18][0] ),
    .CLK(clknet_leaf_19_clk_regs));
 sg13g2_dfrbpq_1 _09981_ (.RESET_B(net1266),
    .D(_00120_),
    .Q(\rf_ram.RAM[18][1] ),
    .CLK(clknet_leaf_54_clk_regs));
 sg13g2_dfrbpq_1 _09982_ (.RESET_B(net1265),
    .D(_00121_),
    .Q(\rf_ram.RAM[18][2] ),
    .CLK(clknet_leaf_68_clk_regs));
 sg13g2_dfrbpq_1 _09983_ (.RESET_B(net1264),
    .D(_00122_),
    .Q(\rf_ram.RAM[18][3] ),
    .CLK(clknet_leaf_87_clk_regs));
 sg13g2_dfrbpq_1 _09984_ (.RESET_B(net1263),
    .D(_00123_),
    .Q(\rf_ram.RAM[18][4] ),
    .CLK(clknet_leaf_87_clk_regs));
 sg13g2_dfrbpq_1 _09985_ (.RESET_B(net1262),
    .D(_00124_),
    .Q(\rf_ram.RAM[18][5] ),
    .CLK(clknet_leaf_88_clk_regs));
 sg13g2_dfrbpq_1 _09986_ (.RESET_B(net1261),
    .D(_00125_),
    .Q(\rf_ram.RAM[18][6] ),
    .CLK(clknet_leaf_92_clk_regs));
 sg13g2_dfrbpq_1 _09987_ (.RESET_B(net1260),
    .D(_00126_),
    .Q(\rf_ram.RAM[18][7] ),
    .CLK(clknet_leaf_95_clk_regs));
 sg13g2_dfrbpq_1 _09988_ (.RESET_B(net1259),
    .D(_00127_),
    .Q(\rf_ram.RAM[18][8] ),
    .CLK(clknet_leaf_115_clk_regs));
 sg13g2_dfrbpq_1 _09989_ (.RESET_B(net1258),
    .D(_00128_),
    .Q(\rf_ram.RAM[18][9] ),
    .CLK(clknet_leaf_126_clk_regs));
 sg13g2_dfrbpq_1 _09990_ (.RESET_B(net1257),
    .D(_00129_),
    .Q(\rf_ram.RAM[18][10] ),
    .CLK(clknet_leaf_118_clk_regs));
 sg13g2_dfrbpq_1 _09991_ (.RESET_B(net1256),
    .D(_00130_),
    .Q(\rf_ram.RAM[18][11] ),
    .CLK(clknet_leaf_134_clk_regs));
 sg13g2_dfrbpq_1 _09992_ (.RESET_B(net1255),
    .D(_00131_),
    .Q(\rf_ram.RAM[18][12] ),
    .CLK(clknet_leaf_126_clk_regs));
 sg13g2_dfrbpq_1 _09993_ (.RESET_B(net1254),
    .D(_00132_),
    .Q(\rf_ram.RAM[18][13] ),
    .CLK(clknet_leaf_144_clk_regs));
 sg13g2_dfrbpq_1 _09994_ (.RESET_B(net1253),
    .D(_00133_),
    .Q(\rf_ram.RAM[18][14] ),
    .CLK(clknet_leaf_159_clk_regs));
 sg13g2_dfrbpq_1 _09995_ (.RESET_B(net1252),
    .D(_00134_),
    .Q(\rf_ram.RAM[18][15] ),
    .CLK(clknet_leaf_144_clk_regs));
 sg13g2_dfrbpq_1 _09996_ (.RESET_B(net1251),
    .D(_00135_),
    .Q(\rf_ram.RAM[18][16] ),
    .CLK(clknet_leaf_104_clk_regs));
 sg13g2_dfrbpq_1 _09997_ (.RESET_B(net1250),
    .D(_00136_),
    .Q(\rf_ram.RAM[18][17] ),
    .CLK(clknet_leaf_138_clk_regs));
 sg13g2_dfrbpq_1 _09998_ (.RESET_B(net1249),
    .D(_00137_),
    .Q(\rf_ram.RAM[18][18] ),
    .CLK(clknet_leaf_137_clk_regs));
 sg13g2_dfrbpq_1 _09999_ (.RESET_B(net1248),
    .D(_00138_),
    .Q(\rf_ram.RAM[18][19] ),
    .CLK(clknet_leaf_160_clk_regs));
 sg13g2_dfrbpq_1 _10000_ (.RESET_B(net1247),
    .D(_00139_),
    .Q(\rf_ram.RAM[18][20] ),
    .CLK(clknet_leaf_149_clk_regs));
 sg13g2_dfrbpq_1 _10001_ (.RESET_B(net1246),
    .D(_00140_),
    .Q(\rf_ram.RAM[18][21] ),
    .CLK(clknet_leaf_62_clk_regs));
 sg13g2_dfrbpq_1 _10002_ (.RESET_B(net1245),
    .D(_00141_),
    .Q(\rf_ram.RAM[18][22] ),
    .CLK(clknet_leaf_104_clk_regs));
 sg13g2_dfrbpq_1 _10003_ (.RESET_B(net1244),
    .D(_00142_),
    .Q(\rf_ram.RAM[18][23] ),
    .CLK(clknet_leaf_22_clk_regs));
 sg13g2_dfrbpq_1 _10004_ (.RESET_B(net1243),
    .D(_00143_),
    .Q(\rf_ram.RAM[18][24] ),
    .CLK(clknet_leaf_71_clk_regs));
 sg13g2_dfrbpq_1 _10005_ (.RESET_B(net1242),
    .D(_00144_),
    .Q(\rf_ram.RAM[18][25] ),
    .CLK(clknet_leaf_56_clk_regs));
 sg13g2_dfrbpq_1 _10006_ (.RESET_B(net1241),
    .D(_00145_),
    .Q(\rf_ram.RAM[18][26] ),
    .CLK(clknet_leaf_56_clk_regs));
 sg13g2_dfrbpq_1 _10007_ (.RESET_B(net1240),
    .D(_00146_),
    .Q(\rf_ram.RAM[18][27] ),
    .CLK(clknet_leaf_46_clk_regs));
 sg13g2_dfrbpq_1 _10008_ (.RESET_B(net1239),
    .D(_00147_),
    .Q(\rf_ram.RAM[18][28] ),
    .CLK(clknet_leaf_24_clk_regs));
 sg13g2_dfrbpq_1 _10009_ (.RESET_B(net1238),
    .D(_00148_),
    .Q(\rf_ram.RAM[18][29] ),
    .CLK(clknet_leaf_170_clk_regs));
 sg13g2_dfrbpq_1 _10010_ (.RESET_B(net1237),
    .D(_00149_),
    .Q(\rf_ram.RAM[18][30] ),
    .CLK(clknet_leaf_163_clk_regs));
 sg13g2_dfrbpq_1 _10011_ (.RESET_B(net1236),
    .D(_00150_),
    .Q(\rf_ram.RAM[18][31] ),
    .CLK(clknet_leaf_169_clk_regs));
 sg13g2_dfrbpq_1 _10012_ (.RESET_B(net1235),
    .D(net2741),
    .Q(\rf_ram.RAM[1][0] ),
    .CLK(clknet_leaf_14_clk_regs));
 sg13g2_dfrbpq_1 _10013_ (.RESET_B(net1234),
    .D(_00152_),
    .Q(\rf_ram.RAM[1][1] ),
    .CLK(clknet_leaf_56_clk_regs));
 sg13g2_dfrbpq_1 _10014_ (.RESET_B(net1233),
    .D(_00153_),
    .Q(\rf_ram.RAM[1][2] ),
    .CLK(clknet_leaf_76_clk_regs));
 sg13g2_dfrbpq_1 _10015_ (.RESET_B(net1232),
    .D(_00154_),
    .Q(\rf_ram.RAM[1][3] ),
    .CLK(clknet_leaf_68_clk_regs));
 sg13g2_dfrbpq_1 _10016_ (.RESET_B(net1231),
    .D(_00155_),
    .Q(\rf_ram.RAM[1][4] ),
    .CLK(clknet_leaf_82_clk_regs));
 sg13g2_dfrbpq_1 _10017_ (.RESET_B(net1230),
    .D(_00156_),
    .Q(\rf_ram.RAM[1][5] ),
    .CLK(clknet_leaf_83_clk_regs));
 sg13g2_dfrbpq_1 _10018_ (.RESET_B(net1229),
    .D(_00157_),
    .Q(\rf_ram.RAM[1][6] ),
    .CLK(clknet_leaf_90_clk_regs));
 sg13g2_dfrbpq_1 _10019_ (.RESET_B(net1228),
    .D(_00158_),
    .Q(\rf_ram.RAM[1][7] ),
    .CLK(clknet_leaf_100_clk_regs));
 sg13g2_dfrbpq_1 _10020_ (.RESET_B(net1227),
    .D(_00159_),
    .Q(\rf_ram.RAM[1][8] ),
    .CLK(clknet_leaf_112_clk_regs));
 sg13g2_dfrbpq_1 _10021_ (.RESET_B(net1226),
    .D(_00160_),
    .Q(\rf_ram.RAM[1][9] ),
    .CLK(clknet_leaf_130_clk_regs));
 sg13g2_dfrbpq_1 _10022_ (.RESET_B(net1225),
    .D(_00161_),
    .Q(\rf_ram.RAM[1][10] ),
    .CLK(clknet_leaf_121_clk_regs));
 sg13g2_dfrbpq_1 _10023_ (.RESET_B(net1224),
    .D(_00162_),
    .Q(\rf_ram.RAM[1][11] ),
    .CLK(clknet_leaf_129_clk_regs));
 sg13g2_dfrbpq_1 _10024_ (.RESET_B(net1223),
    .D(_00163_),
    .Q(\rf_ram.RAM[1][12] ),
    .CLK(clknet_leaf_128_clk_regs));
 sg13g2_dfrbpq_1 _10025_ (.RESET_B(net1222),
    .D(_00164_),
    .Q(\rf_ram.RAM[1][13] ),
    .CLK(clknet_leaf_121_clk_regs));
 sg13g2_dfrbpq_1 _10026_ (.RESET_B(net1221),
    .D(_00165_),
    .Q(\rf_ram.RAM[1][14] ),
    .CLK(clknet_leaf_161_clk_regs));
 sg13g2_dfrbpq_1 _10027_ (.RESET_B(net1188),
    .D(_00166_),
    .Q(\rf_ram.RAM[1][15] ),
    .CLK(clknet_leaf_148_clk_regs));
 sg13g2_dfrbpq_1 _10028_ (.RESET_B(net1187),
    .D(_00167_),
    .Q(\rf_ram.RAM[1][16] ),
    .CLK(clknet_leaf_102_clk_regs));
 sg13g2_dfrbpq_1 _10029_ (.RESET_B(net1185),
    .D(_00168_),
    .Q(\rf_ram.RAM[1][17] ),
    .CLK(clknet_leaf_137_clk_regs));
 sg13g2_dfrbpq_1 _10030_ (.RESET_B(net1184),
    .D(_00169_),
    .Q(\rf_ram.RAM[1][18] ),
    .CLK(clknet_leaf_136_clk_regs));
 sg13g2_dfrbpq_1 _10031_ (.RESET_B(net1183),
    .D(_00170_),
    .Q(\rf_ram.RAM[1][19] ),
    .CLK(clknet_leaf_156_clk_regs));
 sg13g2_dfrbpq_1 _10032_ (.RESET_B(net1181),
    .D(_00171_),
    .Q(\rf_ram.RAM[1][20] ),
    .CLK(clknet_leaf_20_clk_regs));
 sg13g2_dfrbpq_1 _10033_ (.RESET_B(net1180),
    .D(_00172_),
    .Q(\rf_ram.RAM[1][21] ),
    .CLK(clknet_leaf_61_clk_regs));
 sg13g2_dfrbpq_1 _10034_ (.RESET_B(net1179),
    .D(_00173_),
    .Q(\rf_ram.RAM[1][22] ),
    .CLK(clknet_leaf_64_clk_regs));
 sg13g2_dfrbpq_1 _10035_ (.RESET_B(net1178),
    .D(_00174_),
    .Q(\rf_ram.RAM[1][23] ),
    .CLK(clknet_leaf_17_clk_regs));
 sg13g2_dfrbpq_1 _10036_ (.RESET_B(net1177),
    .D(_00175_),
    .Q(\rf_ram.RAM[1][24] ),
    .CLK(clknet_leaf_74_clk_regs));
 sg13g2_dfrbpq_1 _10037_ (.RESET_B(net1176),
    .D(_00176_),
    .Q(\rf_ram.RAM[1][25] ),
    .CLK(clknet_leaf_46_clk_regs));
 sg13g2_dfrbpq_1 _10038_ (.RESET_B(net1175),
    .D(_00177_),
    .Q(\rf_ram.RAM[1][26] ),
    .CLK(clknet_leaf_57_clk_regs));
 sg13g2_dfrbpq_1 _10039_ (.RESET_B(net1174),
    .D(_00178_),
    .Q(\rf_ram.RAM[1][27] ),
    .CLK(clknet_leaf_45_clk_regs));
 sg13g2_dfrbpq_1 _10040_ (.RESET_B(net1173),
    .D(_00179_),
    .Q(\rf_ram.RAM[1][28] ),
    .CLK(clknet_leaf_28_clk_regs));
 sg13g2_dfrbpq_1 _10041_ (.RESET_B(net1172),
    .D(_00180_),
    .Q(\rf_ram.RAM[1][29] ),
    .CLK(clknet_leaf_170_clk_regs));
 sg13g2_dfrbpq_1 _10042_ (.RESET_B(net1171),
    .D(_00181_),
    .Q(\rf_ram.RAM[1][30] ),
    .CLK(clknet_leaf_163_clk_regs));
 sg13g2_dfrbpq_1 _10043_ (.RESET_B(net1170),
    .D(_00182_),
    .Q(\rf_ram.RAM[1][31] ),
    .CLK(clknet_leaf_3_clk_regs));
 sg13g2_dfrbpq_1 _10044_ (.RESET_B(net1169),
    .D(net1576),
    .Q(\rf_ram.RAM[20][0] ),
    .CLK(clknet_leaf_16_clk_regs));
 sg13g2_dfrbpq_1 _10045_ (.RESET_B(net1168),
    .D(_00184_),
    .Q(\rf_ram.RAM[20][1] ),
    .CLK(clknet_leaf_51_clk_regs));
 sg13g2_dfrbpq_1 _10046_ (.RESET_B(net1167),
    .D(_00185_),
    .Q(\rf_ram.RAM[20][2] ),
    .CLK(clknet_leaf_76_clk_regs));
 sg13g2_dfrbpq_1 _10047_ (.RESET_B(net1166),
    .D(_00186_),
    .Q(\rf_ram.RAM[20][3] ),
    .CLK(clknet_leaf_81_clk_regs));
 sg13g2_dfrbpq_1 _10048_ (.RESET_B(net1165),
    .D(_00187_),
    .Q(\rf_ram.RAM[20][4] ),
    .CLK(clknet_leaf_76_clk_regs));
 sg13g2_dfrbpq_1 _10049_ (.RESET_B(net1164),
    .D(_00188_),
    .Q(\rf_ram.RAM[20][5] ),
    .CLK(clknet_leaf_84_clk_regs));
 sg13g2_dfrbpq_1 _10050_ (.RESET_B(net1163),
    .D(_00189_),
    .Q(\rf_ram.RAM[20][6] ),
    .CLK(clknet_leaf_90_clk_regs));
 sg13g2_dfrbpq_1 _10051_ (.RESET_B(net1162),
    .D(_00190_),
    .Q(\rf_ram.RAM[20][7] ),
    .CLK(clknet_leaf_96_clk_regs));
 sg13g2_dfrbpq_1 _10052_ (.RESET_B(net1161),
    .D(_00191_),
    .Q(\rf_ram.RAM[20][8] ),
    .CLK(clknet_leaf_116_clk_regs));
 sg13g2_dfrbpq_1 _10053_ (.RESET_B(net1160),
    .D(_00192_),
    .Q(\rf_ram.RAM[20][9] ),
    .CLK(clknet_leaf_121_clk_regs));
 sg13g2_dfrbpq_1 _10054_ (.RESET_B(net1159),
    .D(_00193_),
    .Q(\rf_ram.RAM[20][10] ),
    .CLK(clknet_leaf_119_clk_regs));
 sg13g2_dfrbpq_1 _10055_ (.RESET_B(net1158),
    .D(_00194_),
    .Q(\rf_ram.RAM[20][11] ),
    .CLK(clknet_leaf_132_clk_regs));
 sg13g2_dfrbpq_1 _10056_ (.RESET_B(net1157),
    .D(_00195_),
    .Q(\rf_ram.RAM[20][12] ),
    .CLK(clknet_leaf_123_clk_regs));
 sg13g2_dfrbpq_1 _10057_ (.RESET_B(net1156),
    .D(_00196_),
    .Q(\rf_ram.RAM[20][13] ),
    .CLK(clknet_leaf_110_clk_regs));
 sg13g2_dfrbpq_1 _10058_ (.RESET_B(net1155),
    .D(_00197_),
    .Q(\rf_ram.RAM[20][14] ),
    .CLK(clknet_leaf_140_clk_regs));
 sg13g2_dfrbpq_1 _10059_ (.RESET_B(net1154),
    .D(_00198_),
    .Q(\rf_ram.RAM[20][15] ),
    .CLK(clknet_leaf_147_clk_regs));
 sg13g2_dfrbpq_1 _10060_ (.RESET_B(net1153),
    .D(_00199_),
    .Q(\rf_ram.RAM[20][16] ),
    .CLK(clknet_leaf_67_clk_regs));
 sg13g2_dfrbpq_1 _10061_ (.RESET_B(net1152),
    .D(_00200_),
    .Q(\rf_ram.RAM[20][17] ),
    .CLK(clknet_leaf_142_clk_regs));
 sg13g2_dfrbpq_1 _10062_ (.RESET_B(net1151),
    .D(_00201_),
    .Q(\rf_ram.RAM[20][18] ),
    .CLK(clknet_leaf_139_clk_regs));
 sg13g2_dfrbpq_1 _10063_ (.RESET_B(net1150),
    .D(_00202_),
    .Q(\rf_ram.RAM[20][19] ),
    .CLK(clknet_leaf_152_clk_regs));
 sg13g2_dfrbpq_1 _10064_ (.RESET_B(net1149),
    .D(_00203_),
    .Q(\rf_ram.RAM[20][20] ),
    .CLK(clknet_leaf_151_clk_regs));
 sg13g2_dfrbpq_1 _10065_ (.RESET_B(net1088),
    .D(_00204_),
    .Q(\rf_ram.RAM[20][21] ),
    .CLK(clknet_leaf_60_clk_regs));
 sg13g2_dfrbpq_1 _10066_ (.RESET_B(net1087),
    .D(_00205_),
    .Q(\rf_ram.RAM[20][22] ),
    .CLK(clknet_leaf_66_clk_regs));
 sg13g2_dfrbpq_1 _10067_ (.RESET_B(net1086),
    .D(_00206_),
    .Q(\rf_ram.RAM[20][23] ),
    .CLK(clknet_leaf_25_clk_regs));
 sg13g2_dfrbpq_1 _10068_ (.RESET_B(net1085),
    .D(_00207_),
    .Q(\rf_ram.RAM[20][24] ),
    .CLK(clknet_leaf_73_clk_regs));
 sg13g2_dfrbpq_1 _10069_ (.RESET_B(net1084),
    .D(_00208_),
    .Q(\rf_ram.RAM[20][25] ),
    .CLK(clknet_leaf_49_clk_regs));
 sg13g2_dfrbpq_1 _10070_ (.RESET_B(net1083),
    .D(_00209_),
    .Q(\rf_ram.RAM[20][26] ),
    .CLK(clknet_leaf_49_clk_regs));
 sg13g2_dfrbpq_1 _10071_ (.RESET_B(net1082),
    .D(_00210_),
    .Q(\rf_ram.RAM[20][27] ),
    .CLK(clknet_leaf_43_clk_regs));
 sg13g2_dfrbpq_1 _10072_ (.RESET_B(net1081),
    .D(_00211_),
    .Q(\rf_ram.RAM[20][28] ),
    .CLK(clknet_leaf_26_clk_regs));
 sg13g2_dfrbpq_1 _10073_ (.RESET_B(net1080),
    .D(_00212_),
    .Q(\rf_ram.RAM[20][29] ),
    .CLK(clknet_leaf_4_clk_regs));
 sg13g2_dfrbpq_1 _10074_ (.RESET_B(net1079),
    .D(_00213_),
    .Q(\rf_ram.RAM[20][30] ),
    .CLK(clknet_leaf_165_clk_regs));
 sg13g2_dfrbpq_1 _10075_ (.RESET_B(net1078),
    .D(_00214_),
    .Q(\rf_ram.RAM[20][31] ),
    .CLK(clknet_leaf_4_clk_regs));
 sg13g2_dfrbpq_1 _10076_ (.RESET_B(net1077),
    .D(net3272),
    .Q(\rf_ram.RAM[21][0] ),
    .CLK(clknet_leaf_16_clk_regs));
 sg13g2_dfrbpq_1 _10077_ (.RESET_B(net1076),
    .D(_00216_),
    .Q(\rf_ram.RAM[21][1] ),
    .CLK(clknet_leaf_51_clk_regs));
 sg13g2_dfrbpq_1 _10078_ (.RESET_B(net1075),
    .D(_00217_),
    .Q(\rf_ram.RAM[21][2] ),
    .CLK(clknet_leaf_75_clk_regs));
 sg13g2_dfrbpq_1 _10079_ (.RESET_B(net1074),
    .D(_00218_),
    .Q(\rf_ram.RAM[21][3] ),
    .CLK(clknet_leaf_83_clk_regs));
 sg13g2_dfrbpq_1 _10080_ (.RESET_B(net1073),
    .D(_00219_),
    .Q(\rf_ram.RAM[21][4] ),
    .CLK(clknet_leaf_76_clk_regs));
 sg13g2_dfrbpq_1 _10081_ (.RESET_B(net1072),
    .D(_00220_),
    .Q(\rf_ram.RAM[21][5] ),
    .CLK(clknet_leaf_84_clk_regs));
 sg13g2_dfrbpq_1 _10082_ (.RESET_B(net1071),
    .D(_00221_),
    .Q(\rf_ram.RAM[21][6] ),
    .CLK(clknet_leaf_90_clk_regs));
 sg13g2_dfrbpq_1 _10083_ (.RESET_B(net1070),
    .D(_00222_),
    .Q(\rf_ram.RAM[21][7] ),
    .CLK(clknet_leaf_95_clk_regs));
 sg13g2_dfrbpq_1 _10084_ (.RESET_B(net1069),
    .D(_00223_),
    .Q(\rf_ram.RAM[21][8] ),
    .CLK(clknet_leaf_112_clk_regs));
 sg13g2_dfrbpq_1 _10085_ (.RESET_B(net1068),
    .D(_00224_),
    .Q(\rf_ram.RAM[21][9] ),
    .CLK(clknet_leaf_122_clk_regs));
 sg13g2_dfrbpq_1 _10086_ (.RESET_B(net1067),
    .D(_00225_),
    .Q(\rf_ram.RAM[21][10] ),
    .CLK(clknet_leaf_119_clk_regs));
 sg13g2_dfrbpq_1 _10087_ (.RESET_B(net1066),
    .D(_00226_),
    .Q(\rf_ram.RAM[21][11] ),
    .CLK(clknet_leaf_134_clk_regs));
 sg13g2_dfrbpq_1 _10088_ (.RESET_B(net1065),
    .D(_00227_),
    .Q(\rf_ram.RAM[21][12] ),
    .CLK(clknet_leaf_118_clk_regs));
 sg13g2_dfrbpq_1 _10089_ (.RESET_B(net1064),
    .D(_00228_),
    .Q(\rf_ram.RAM[21][13] ),
    .CLK(clknet_leaf_108_clk_regs));
 sg13g2_dfrbpq_1 _10090_ (.RESET_B(net1063),
    .D(_00229_),
    .Q(\rf_ram.RAM[21][14] ),
    .CLK(clknet_leaf_156_clk_regs));
 sg13g2_dfrbpq_1 _10091_ (.RESET_B(net1062),
    .D(_00230_),
    .Q(\rf_ram.RAM[21][15] ),
    .CLK(clknet_leaf_147_clk_regs));
 sg13g2_dfrbpq_1 _10092_ (.RESET_B(net1061),
    .D(_00231_),
    .Q(\rf_ram.RAM[21][16] ),
    .CLK(clknet_leaf_67_clk_regs));
 sg13g2_dfrbpq_1 _10093_ (.RESET_B(net1060),
    .D(_00232_),
    .Q(\rf_ram.RAM[21][17] ),
    .CLK(clknet_leaf_142_clk_regs));
 sg13g2_dfrbpq_1 _10094_ (.RESET_B(net1059),
    .D(_00233_),
    .Q(\rf_ram.RAM[21][18] ),
    .CLK(clknet_leaf_137_clk_regs));
 sg13g2_dfrbpq_1 _10095_ (.RESET_B(net1058),
    .D(_00234_),
    .Q(\rf_ram.RAM[21][19] ),
    .CLK(clknet_leaf_156_clk_regs));
 sg13g2_dfrbpq_1 _10096_ (.RESET_B(net1057),
    .D(_00235_),
    .Q(\rf_ram.RAM[21][20] ),
    .CLK(clknet_leaf_150_clk_regs));
 sg13g2_dfrbpq_1 _10097_ (.RESET_B(net1056),
    .D(_00236_),
    .Q(\rf_ram.RAM[21][21] ),
    .CLK(clknet_leaf_60_clk_regs));
 sg13g2_dfrbpq_1 _10098_ (.RESET_B(net1055),
    .D(_00237_),
    .Q(\rf_ram.RAM[21][22] ),
    .CLK(clknet_leaf_66_clk_regs));
 sg13g2_dfrbpq_1 _10099_ (.RESET_B(net1054),
    .D(_00238_),
    .Q(\rf_ram.RAM[21][23] ),
    .CLK(clknet_leaf_26_clk_regs));
 sg13g2_dfrbpq_1 _10100_ (.RESET_B(net1053),
    .D(_00239_),
    .Q(\rf_ram.RAM[21][24] ),
    .CLK(clknet_leaf_75_clk_regs));
 sg13g2_dfrbpq_1 _10101_ (.RESET_B(net1052),
    .D(_00240_),
    .Q(\rf_ram.RAM[21][25] ),
    .CLK(clknet_leaf_48_clk_regs));
 sg13g2_dfrbpq_1 _10102_ (.RESET_B(net1051),
    .D(_00241_),
    .Q(\rf_ram.RAM[21][26] ),
    .CLK(clknet_leaf_48_clk_regs));
 sg13g2_dfrbpq_1 _10103_ (.RESET_B(net1050),
    .D(_00242_),
    .Q(\rf_ram.RAM[21][27] ),
    .CLK(clknet_leaf_42_clk_regs));
 sg13g2_dfrbpq_1 _10104_ (.RESET_B(net1049),
    .D(_00243_),
    .Q(\rf_ram.RAM[21][28] ),
    .CLK(clknet_leaf_27_clk_regs));
 sg13g2_dfrbpq_1 _10105_ (.RESET_B(net1048),
    .D(_00244_),
    .Q(\rf_ram.RAM[21][29] ),
    .CLK(clknet_leaf_4_clk_regs));
 sg13g2_dfrbpq_1 _10106_ (.RESET_B(net1047),
    .D(_00245_),
    .Q(\rf_ram.RAM[21][30] ),
    .CLK(clknet_leaf_165_clk_regs));
 sg13g2_dfrbpq_1 _10107_ (.RESET_B(net1046),
    .D(_00246_),
    .Q(\rf_ram.RAM[21][31] ),
    .CLK(clknet_leaf_5_clk_regs));
 sg13g2_dfrbpq_1 _10108_ (.RESET_B(net1045),
    .D(net1697),
    .Q(\rf_ram.RAM[22][0] ),
    .CLK(clknet_leaf_16_clk_regs));
 sg13g2_dfrbpq_1 _10109_ (.RESET_B(net1044),
    .D(_00248_),
    .Q(\rf_ram.RAM[22][1] ),
    .CLK(clknet_leaf_51_clk_regs));
 sg13g2_dfrbpq_1 _10110_ (.RESET_B(net1043),
    .D(_00249_),
    .Q(\rf_ram.RAM[22][2] ),
    .CLK(clknet_leaf_75_clk_regs));
 sg13g2_dfrbpq_1 _10111_ (.RESET_B(net1042),
    .D(_00250_),
    .Q(\rf_ram.RAM[22][3] ),
    .CLK(clknet_leaf_83_clk_regs));
 sg13g2_dfrbpq_1 _10112_ (.RESET_B(net1041),
    .D(_00251_),
    .Q(\rf_ram.RAM[22][4] ),
    .CLK(clknet_leaf_76_clk_regs));
 sg13g2_dfrbpq_1 _10113_ (.RESET_B(net1040),
    .D(_00252_),
    .Q(\rf_ram.RAM[22][5] ),
    .CLK(clknet_leaf_83_clk_regs));
 sg13g2_dfrbpq_1 _10114_ (.RESET_B(net1039),
    .D(_00253_),
    .Q(\rf_ram.RAM[22][6] ),
    .CLK(clknet_leaf_90_clk_regs));
 sg13g2_dfrbpq_1 _10115_ (.RESET_B(net1038),
    .D(_00254_),
    .Q(\rf_ram.RAM[22][7] ),
    .CLK(clknet_leaf_115_clk_regs));
 sg13g2_dfrbpq_1 _10116_ (.RESET_B(net1037),
    .D(_00255_),
    .Q(\rf_ram.RAM[22][8] ),
    .CLK(clknet_leaf_112_clk_regs));
 sg13g2_dfrbpq_1 _10117_ (.RESET_B(net1036),
    .D(_00256_),
    .Q(\rf_ram.RAM[22][9] ),
    .CLK(clknet_leaf_121_clk_regs));
 sg13g2_dfrbpq_1 _10118_ (.RESET_B(net1035),
    .D(_00257_),
    .Q(\rf_ram.RAM[22][10] ),
    .CLK(clknet_leaf_117_clk_regs));
 sg13g2_dfrbpq_1 _10119_ (.RESET_B(net1034),
    .D(_00258_),
    .Q(\rf_ram.RAM[22][11] ),
    .CLK(clknet_leaf_129_clk_regs));
 sg13g2_dfrbpq_1 _10120_ (.RESET_B(net1033),
    .D(_00259_),
    .Q(\rf_ram.RAM[22][12] ),
    .CLK(clknet_leaf_123_clk_regs));
 sg13g2_dfrbpq_1 _10121_ (.RESET_B(net1032),
    .D(_00260_),
    .Q(\rf_ram.RAM[22][13] ),
    .CLK(clknet_leaf_110_clk_regs));
 sg13g2_dfrbpq_1 _10122_ (.RESET_B(net1031),
    .D(_00261_),
    .Q(\rf_ram.RAM[22][14] ),
    .CLK(clknet_leaf_157_clk_regs));
 sg13g2_dfrbpq_1 _10123_ (.RESET_B(net1030),
    .D(_00262_),
    .Q(\rf_ram.RAM[22][15] ),
    .CLK(clknet_leaf_147_clk_regs));
 sg13g2_dfrbpq_1 _10124_ (.RESET_B(net1029),
    .D(_00263_),
    .Q(\rf_ram.RAM[22][16] ),
    .CLK(clknet_leaf_67_clk_regs));
 sg13g2_dfrbpq_1 _10125_ (.RESET_B(net1028),
    .D(_00264_),
    .Q(\rf_ram.RAM[22][17] ),
    .CLK(clknet_leaf_142_clk_regs));
 sg13g2_dfrbpq_1 _10126_ (.RESET_B(net1027),
    .D(_00265_),
    .Q(\rf_ram.RAM[22][18] ),
    .CLK(clknet_leaf_136_clk_regs));
 sg13g2_dfrbpq_1 _10127_ (.RESET_B(net1026),
    .D(_00266_),
    .Q(\rf_ram.RAM[22][19] ),
    .CLK(clknet_leaf_156_clk_regs));
 sg13g2_dfrbpq_1 _10128_ (.RESET_B(net1025),
    .D(_00267_),
    .Q(\rf_ram.RAM[22][20] ),
    .CLK(clknet_leaf_150_clk_regs));
 sg13g2_dfrbpq_1 _10129_ (.RESET_B(net1024),
    .D(_00268_),
    .Q(\rf_ram.RAM[22][21] ),
    .CLK(clknet_leaf_59_clk_regs));
 sg13g2_dfrbpq_1 _10130_ (.RESET_B(net1023),
    .D(_00269_),
    .Q(\rf_ram.RAM[22][22] ),
    .CLK(clknet_leaf_66_clk_regs));
 sg13g2_dfrbpq_1 _10131_ (.RESET_B(net1022),
    .D(_00270_),
    .Q(\rf_ram.RAM[22][23] ),
    .CLK(clknet_leaf_25_clk_regs));
 sg13g2_dfrbpq_1 _10132_ (.RESET_B(net1021),
    .D(_00271_),
    .Q(\rf_ram.RAM[22][24] ),
    .CLK(clknet_leaf_74_clk_regs));
 sg13g2_dfrbpq_1 _10133_ (.RESET_B(net1020),
    .D(_00272_),
    .Q(\rf_ram.RAM[22][25] ),
    .CLK(clknet_leaf_48_clk_regs));
 sg13g2_dfrbpq_1 _10134_ (.RESET_B(net1019),
    .D(_00273_),
    .Q(\rf_ram.RAM[22][26] ),
    .CLK(clknet_leaf_48_clk_regs));
 sg13g2_dfrbpq_1 _10135_ (.RESET_B(net1018),
    .D(_00274_),
    .Q(\rf_ram.RAM[22][27] ),
    .CLK(clknet_leaf_43_clk_regs));
 sg13g2_dfrbpq_1 _10136_ (.RESET_B(net1017),
    .D(_00275_),
    .Q(\rf_ram.RAM[22][28] ),
    .CLK(clknet_leaf_26_clk_regs));
 sg13g2_dfrbpq_1 _10137_ (.RESET_B(net1016),
    .D(_00276_),
    .Q(\rf_ram.RAM[22][29] ),
    .CLK(clknet_leaf_4_clk_regs));
 sg13g2_dfrbpq_1 _10138_ (.RESET_B(net1015),
    .D(_00277_),
    .Q(\rf_ram.RAM[22][30] ),
    .CLK(clknet_leaf_154_clk_regs));
 sg13g2_dfrbpq_1 _10139_ (.RESET_B(net1014),
    .D(_00278_),
    .Q(\rf_ram.RAM[22][31] ),
    .CLK(clknet_leaf_5_clk_regs));
 sg13g2_dfrbpq_1 _10140_ (.RESET_B(net1013),
    .D(_00279_),
    .Q(\rf_ram.RAM[23][0] ),
    .CLK(clknet_leaf_15_clk_regs));
 sg13g2_dfrbpq_1 _10141_ (.RESET_B(net1012),
    .D(_00280_),
    .Q(\rf_ram.RAM[23][1] ),
    .CLK(clknet_leaf_51_clk_regs));
 sg13g2_dfrbpq_1 _10142_ (.RESET_B(net1011),
    .D(_00281_),
    .Q(\rf_ram.RAM[23][2] ),
    .CLK(clknet_leaf_76_clk_regs));
 sg13g2_dfrbpq_1 _10143_ (.RESET_B(net1010),
    .D(_00282_),
    .Q(\rf_ram.RAM[23][3] ),
    .CLK(clknet_leaf_81_clk_regs));
 sg13g2_dfrbpq_1 _10144_ (.RESET_B(net1009),
    .D(_00283_),
    .Q(\rf_ram.RAM[23][4] ),
    .CLK(clknet_leaf_77_clk_regs));
 sg13g2_dfrbpq_1 _10145_ (.RESET_B(net1008),
    .D(_00284_),
    .Q(\rf_ram.RAM[23][5] ),
    .CLK(clknet_leaf_84_clk_regs));
 sg13g2_dfrbpq_1 _10146_ (.RESET_B(net1007),
    .D(_00285_),
    .Q(\rf_ram.RAM[23][6] ),
    .CLK(clknet_leaf_91_clk_regs));
 sg13g2_dfrbpq_1 _10147_ (.RESET_B(net1006),
    .D(_00286_),
    .Q(\rf_ram.RAM[23][7] ),
    .CLK(clknet_leaf_115_clk_regs));
 sg13g2_dfrbpq_1 _10148_ (.RESET_B(net1005),
    .D(_00287_),
    .Q(\rf_ram.RAM[23][8] ),
    .CLK(clknet_leaf_114_clk_regs));
 sg13g2_dfrbpq_1 _10149_ (.RESET_B(net1004),
    .D(_00288_),
    .Q(\rf_ram.RAM[23][9] ),
    .CLK(clknet_leaf_122_clk_regs));
 sg13g2_dfrbpq_1 _10150_ (.RESET_B(net1003),
    .D(_00289_),
    .Q(\rf_ram.RAM[23][10] ),
    .CLK(clknet_leaf_119_clk_regs));
 sg13g2_dfrbpq_1 _10151_ (.RESET_B(net1002),
    .D(_00290_),
    .Q(\rf_ram.RAM[23][11] ),
    .CLK(clknet_leaf_134_clk_regs));
 sg13g2_dfrbpq_1 _10152_ (.RESET_B(net1001),
    .D(_00291_),
    .Q(\rf_ram.RAM[23][12] ),
    .CLK(clknet_leaf_122_clk_regs));
 sg13g2_dfrbpq_1 _10153_ (.RESET_B(net1000),
    .D(_00292_),
    .Q(\rf_ram.RAM[23][13] ),
    .CLK(clknet_leaf_111_clk_regs));
 sg13g2_dfrbpq_1 _10154_ (.RESET_B(net999),
    .D(_00293_),
    .Q(\rf_ram.RAM[23][14] ),
    .CLK(clknet_leaf_140_clk_regs));
 sg13g2_dfrbpq_1 _10155_ (.RESET_B(net998),
    .D(_00294_),
    .Q(\rf_ram.RAM[23][15] ),
    .CLK(clknet_leaf_147_clk_regs));
 sg13g2_dfrbpq_1 _10156_ (.RESET_B(net997),
    .D(_00295_),
    .Q(\rf_ram.RAM[23][16] ),
    .CLK(clknet_leaf_67_clk_regs));
 sg13g2_dfrbpq_1 _10157_ (.RESET_B(net996),
    .D(_00296_),
    .Q(\rf_ram.RAM[23][17] ),
    .CLK(clknet_leaf_140_clk_regs));
 sg13g2_dfrbpq_1 _10158_ (.RESET_B(net995),
    .D(_00297_),
    .Q(\rf_ram.RAM[23][18] ),
    .CLK(clknet_leaf_139_clk_regs));
 sg13g2_dfrbpq_1 _10159_ (.RESET_B(net994),
    .D(_00298_),
    .Q(\rf_ram.RAM[23][19] ),
    .CLK(clknet_leaf_156_clk_regs));
 sg13g2_dfrbpq_1 _10160_ (.RESET_B(net993),
    .D(_00299_),
    .Q(\rf_ram.RAM[23][20] ),
    .CLK(clknet_leaf_151_clk_regs));
 sg13g2_dfrbpq_1 _10161_ (.RESET_B(net992),
    .D(_00300_),
    .Q(\rf_ram.RAM[23][21] ),
    .CLK(clknet_leaf_61_clk_regs));
 sg13g2_dfrbpq_1 _10162_ (.RESET_B(net991),
    .D(_00301_),
    .Q(\rf_ram.RAM[23][22] ),
    .CLK(clknet_leaf_66_clk_regs));
 sg13g2_dfrbpq_1 _10163_ (.RESET_B(net990),
    .D(_00302_),
    .Q(\rf_ram.RAM[23][23] ),
    .CLK(clknet_leaf_26_clk_regs));
 sg13g2_dfrbpq_1 _10164_ (.RESET_B(net989),
    .D(_00303_),
    .Q(\rf_ram.RAM[23][24] ),
    .CLK(clknet_leaf_73_clk_regs));
 sg13g2_dfrbpq_1 _10165_ (.RESET_B(net988),
    .D(_00304_),
    .Q(\rf_ram.RAM[23][25] ),
    .CLK(clknet_leaf_49_clk_regs));
 sg13g2_dfrbpq_1 _10166_ (.RESET_B(net987),
    .D(_00305_),
    .Q(\rf_ram.RAM[23][26] ),
    .CLK(clknet_leaf_49_clk_regs));
 sg13g2_dfrbpq_1 _10167_ (.RESET_B(net986),
    .D(_00306_),
    .Q(\rf_ram.RAM[23][27] ),
    .CLK(clknet_leaf_43_clk_regs));
 sg13g2_dfrbpq_1 _10168_ (.RESET_B(net985),
    .D(_00307_),
    .Q(\rf_ram.RAM[23][28] ),
    .CLK(clknet_leaf_35_clk_regs));
 sg13g2_dfrbpq_1 _10169_ (.RESET_B(net984),
    .D(_00308_),
    .Q(\rf_ram.RAM[23][29] ),
    .CLK(clknet_leaf_4_clk_regs));
 sg13g2_dfrbpq_1 _10170_ (.RESET_B(net983),
    .D(_00309_),
    .Q(\rf_ram.RAM[23][30] ),
    .CLK(clknet_leaf_165_clk_regs));
 sg13g2_dfrbpq_1 _10171_ (.RESET_B(net982),
    .D(_00310_),
    .Q(\rf_ram.RAM[23][31] ),
    .CLK(clknet_leaf_4_clk_regs));
 sg13g2_dfrbpq_2 _10172_ (.RESET_B(net981),
    .D(_00311_),
    .Q(\cpu.rf_ram_if.rcnt[0] ),
    .CLK(clknet_leaf_36_clk_regs));
 sg13g2_dfrbpq_1 _10173_ (.RESET_B(net980),
    .D(net3263),
    .Q(\cpu.rf_ram_if.rcnt[2] ),
    .CLK(clknet_leaf_45_clk_regs));
 sg13g2_dfrbpq_1 _10174_ (.RESET_B(net979),
    .D(_00313_),
    .Q(\cpu.rf_ram_if.rcnt[3] ),
    .CLK(clknet_leaf_45_clk_regs));
 sg13g2_dfrbpq_1 _10175_ (.RESET_B(net978),
    .D(_00314_),
    .Q(\cpu.rf_ram_if.rcnt[4] ),
    .CLK(clknet_leaf_44_clk_regs));
 sg13g2_dfrbpq_2 _10176_ (.RESET_B(net977),
    .D(_00315_),
    .Q(\cpu.arbiter.i_wb_mem_rdt[16] ),
    .CLK(clknet_leaf_11_clk_regs));
 sg13g2_dfrbpq_2 _10177_ (.RESET_B(net976),
    .D(net3495),
    .Q(\cpu.arbiter.i_wb_mem_rdt[17] ),
    .CLK(clknet_leaf_6_clk_regs));
 sg13g2_dfrbpq_2 _10178_ (.RESET_B(net975),
    .D(net3486),
    .Q(\cpu.arbiter.i_wb_mem_rdt[18] ),
    .CLK(clknet_leaf_6_clk_regs));
 sg13g2_dfrbpq_2 _10179_ (.RESET_B(net974),
    .D(net3566),
    .Q(\cpu.arbiter.i_wb_mem_rdt[19] ),
    .CLK(clknet_leaf_3_clk_regs));
 sg13g2_dfrbpq_2 _10180_ (.RESET_B(net973),
    .D(_00319_),
    .Q(\cpu.arbiter.i_wb_mem_rdt[20] ),
    .CLK(clknet_leaf_5_clk_regs));
 sg13g2_dfrbpq_2 _10181_ (.RESET_B(net972),
    .D(net3559),
    .Q(\cpu.arbiter.i_wb_mem_rdt[21] ),
    .CLK(clknet_leaf_6_clk_regs));
 sg13g2_dfrbpq_2 _10182_ (.RESET_B(net971),
    .D(_00321_),
    .Q(\cpu.arbiter.i_wb_mem_rdt[22] ),
    .CLK(clknet_leaf_6_clk_regs));
 sg13g2_dfrbpq_2 _10183_ (.RESET_B(net970),
    .D(net3682),
    .Q(\cpu.arbiter.i_wb_mem_rdt[23] ),
    .CLK(clknet_leaf_9_clk_regs));
 sg13g2_dfrbpq_2 _10184_ (.RESET_B(net969),
    .D(_00323_),
    .Q(\cpu.arbiter.i_wb_mem_rdt[24] ),
    .CLK(clknet_leaf_9_clk_regs));
 sg13g2_dfrbpq_2 _10185_ (.RESET_B(net968),
    .D(net3585),
    .Q(\cpu.arbiter.i_wb_mem_rdt[25] ),
    .CLK(clknet_leaf_3_clk_regs));
 sg13g2_dfrbpq_2 _10186_ (.RESET_B(net967),
    .D(net3557),
    .Q(\cpu.arbiter.i_wb_mem_rdt[26] ),
    .CLK(clknet_leaf_1_clk_regs));
 sg13g2_dfrbpq_2 _10187_ (.RESET_B(net966),
    .D(net3537),
    .Q(\cpu.arbiter.i_wb_mem_rdt[27] ),
    .CLK(clknet_leaf_3_clk_regs));
 sg13g2_dfrbpq_2 _10188_ (.RESET_B(net965),
    .D(net3603),
    .Q(\cpu.arbiter.i_wb_mem_rdt[28] ),
    .CLK(clknet_leaf_3_clk_regs));
 sg13g2_dfrbpq_2 _10189_ (.RESET_B(net964),
    .D(net3614),
    .Q(\cpu.arbiter.i_wb_mem_rdt[29] ),
    .CLK(clknet_leaf_7_clk_regs));
 sg13g2_dfrbpq_2 _10190_ (.RESET_B(net963),
    .D(net3593),
    .Q(\cpu.arbiter.i_wb_mem_rdt[30] ),
    .CLK(clknet_leaf_11_clk_regs));
 sg13g2_dfrbpq_2 _10191_ (.RESET_B(net962),
    .D(net3689),
    .Q(\cpu.arbiter.i_wb_mem_rdt[31] ),
    .CLK(clknet_leaf_29_clk_regs));
 sg13g2_dfrbpq_1 _10192_ (.RESET_B(net961),
    .D(_00331_),
    .Q(\cpu.i_wb_ext_rdt[0] ),
    .CLK(clknet_leaf_42_clk_regs));
 sg13g2_dfrbpq_1 _10193_ (.RESET_B(net960),
    .D(_00332_),
    .Q(\cpu.i_wb_ext_rdt[1] ),
    .CLK(clknet_leaf_42_clk_regs));
 sg13g2_dfrbpq_1 _10194_ (.RESET_B(net959),
    .D(_00333_),
    .Q(\cpu.i_wb_ext_rdt[2] ),
    .CLK(clknet_leaf_42_clk_regs));
 sg13g2_dfrbpq_1 _10195_ (.RESET_B(net958),
    .D(_00334_),
    .Q(\cpu.i_wb_ext_rdt[3] ),
    .CLK(clknet_leaf_42_clk_regs));
 sg13g2_dfrbpq_1 _10196_ (.RESET_B(net957),
    .D(_00335_),
    .Q(\cpu.i_wb_ext_rdt[4] ),
    .CLK(clknet_leaf_39_clk_regs));
 sg13g2_dfrbpq_1 _10197_ (.RESET_B(net956),
    .D(_00336_),
    .Q(\cpu.i_wb_ext_rdt[5] ),
    .CLK(clknet_leaf_39_clk_regs));
 sg13g2_dfrbpq_1 _10198_ (.RESET_B(net955),
    .D(_00337_),
    .Q(\cpu.i_wb_ext_rdt[6] ),
    .CLK(clknet_leaf_40_clk_regs));
 sg13g2_dfrbpq_1 _10199_ (.RESET_B(net954),
    .D(_00338_),
    .Q(\cpu.i_wb_ext_rdt[7] ),
    .CLK(clknet_leaf_39_clk_regs));
 sg13g2_dfrbpq_1 _10200_ (.RESET_B(net953),
    .D(net2811),
    .Q(\rf_ram.RAM[31][0] ),
    .CLK(clknet_leaf_153_clk_regs));
 sg13g2_dfrbpq_1 _10201_ (.RESET_B(net952),
    .D(_00340_),
    .Q(\rf_ram.RAM[31][1] ),
    .CLK(clknet_leaf_52_clk_regs));
 sg13g2_dfrbpq_1 _10202_ (.RESET_B(net951),
    .D(_00341_),
    .Q(\rf_ram.RAM[31][2] ),
    .CLK(clknet_leaf_67_clk_regs));
 sg13g2_dfrbpq_1 _10203_ (.RESET_B(net950),
    .D(_00342_),
    .Q(\rf_ram.RAM[31][3] ),
    .CLK(clknet_leaf_89_clk_regs));
 sg13g2_dfrbpq_1 _10204_ (.RESET_B(net949),
    .D(_00343_),
    .Q(\rf_ram.RAM[31][4] ),
    .CLK(clknet_leaf_86_clk_regs));
 sg13g2_dfrbpq_1 _10205_ (.RESET_B(net948),
    .D(_00344_),
    .Q(\rf_ram.RAM[31][5] ),
    .CLK(clknet_leaf_92_clk_regs));
 sg13g2_dfrbpq_1 _10206_ (.RESET_B(net947),
    .D(_00345_),
    .Q(\rf_ram.RAM[31][6] ),
    .CLK(clknet_leaf_93_clk_regs));
 sg13g2_dfrbpq_1 _10207_ (.RESET_B(net946),
    .D(_00346_),
    .Q(\rf_ram.RAM[31][7] ),
    .CLK(clknet_leaf_93_clk_regs));
 sg13g2_dfrbpq_1 _10208_ (.RESET_B(net945),
    .D(_00347_),
    .Q(\rf_ram.RAM[31][8] ),
    .CLK(clknet_leaf_116_clk_regs));
 sg13g2_dfrbpq_1 _10209_ (.RESET_B(net944),
    .D(_00348_),
    .Q(\rf_ram.RAM[31][9] ),
    .CLK(clknet_leaf_124_clk_regs));
 sg13g2_dfrbpq_1 _10210_ (.RESET_B(net943),
    .D(_00349_),
    .Q(\rf_ram.RAM[31][10] ),
    .CLK(clknet_leaf_117_clk_regs));
 sg13g2_dfrbpq_1 _10211_ (.RESET_B(net942),
    .D(_00350_),
    .Q(\rf_ram.RAM[31][11] ),
    .CLK(clknet_leaf_134_clk_regs));
 sg13g2_dfrbpq_1 _10212_ (.RESET_B(net941),
    .D(_00351_),
    .Q(\rf_ram.RAM[31][12] ),
    .CLK(clknet_leaf_123_clk_regs));
 sg13g2_dfrbpq_1 _10213_ (.RESET_B(net940),
    .D(_00352_),
    .Q(\rf_ram.RAM[31][13] ),
    .CLK(clknet_leaf_101_clk_regs));
 sg13g2_dfrbpq_1 _10214_ (.RESET_B(net939),
    .D(_00353_),
    .Q(\rf_ram.RAM[31][14] ),
    .CLK(clknet_leaf_140_clk_regs));
 sg13g2_dfrbpq_1 _10215_ (.RESET_B(net938),
    .D(_00354_),
    .Q(\rf_ram.RAM[31][15] ),
    .CLK(clknet_leaf_109_clk_regs));
 sg13g2_dfrbpq_1 _10216_ (.RESET_B(net937),
    .D(_00355_),
    .Q(\rf_ram.RAM[31][16] ),
    .CLK(clknet_leaf_109_clk_regs));
 sg13g2_dfrbpq_1 _10217_ (.RESET_B(net936),
    .D(_00356_),
    .Q(\rf_ram.RAM[31][17] ),
    .CLK(clknet_leaf_138_clk_regs));
 sg13g2_dfrbpq_1 _10218_ (.RESET_B(net935),
    .D(_00357_),
    .Q(\rf_ram.RAM[31][18] ),
    .CLK(clknet_leaf_136_clk_regs));
 sg13g2_dfrbpq_1 _10219_ (.RESET_B(net934),
    .D(_00358_),
    .Q(\rf_ram.RAM[31][19] ),
    .CLK(clknet_leaf_154_clk_regs));
 sg13g2_dfrbpq_1 _10220_ (.RESET_B(net933),
    .D(_00359_),
    .Q(\rf_ram.RAM[31][20] ),
    .CLK(clknet_leaf_152_clk_regs));
 sg13g2_dfrbpq_1 _10221_ (.RESET_B(net932),
    .D(_00360_),
    .Q(\rf_ram.RAM[31][21] ),
    .CLK(clknet_leaf_65_clk_regs));
 sg13g2_dfrbpq_1 _10222_ (.RESET_B(net931),
    .D(_00361_),
    .Q(\rf_ram.RAM[31][22] ),
    .CLK(clknet_leaf_67_clk_regs));
 sg13g2_dfrbpq_1 _10223_ (.RESET_B(net930),
    .D(_00362_),
    .Q(\rf_ram.RAM[31][23] ),
    .CLK(clknet_leaf_59_clk_regs));
 sg13g2_dfrbpq_1 _10224_ (.RESET_B(net929),
    .D(_00363_),
    .Q(\rf_ram.RAM[31][24] ),
    .CLK(clknet_leaf_73_clk_regs));
 sg13g2_dfrbpq_1 _10225_ (.RESET_B(net928),
    .D(_00364_),
    .Q(\rf_ram.RAM[31][25] ),
    .CLK(clknet_leaf_50_clk_regs));
 sg13g2_dfrbpq_1 _10226_ (.RESET_B(net927),
    .D(_00365_),
    .Q(\rf_ram.RAM[31][26] ),
    .CLK(clknet_leaf_51_clk_regs));
 sg13g2_dfrbpq_1 _10227_ (.RESET_B(net926),
    .D(_00366_),
    .Q(\rf_ram.RAM[31][27] ),
    .CLK(clknet_leaf_43_clk_regs));
 sg13g2_dfrbpq_1 _10228_ (.RESET_B(net925),
    .D(_00367_),
    .Q(\rf_ram.RAM[31][28] ),
    .CLK(clknet_leaf_26_clk_regs));
 sg13g2_dfrbpq_1 _10229_ (.RESET_B(net924),
    .D(_00368_),
    .Q(\rf_ram.RAM[31][29] ),
    .CLK(clknet_leaf_154_clk_regs));
 sg13g2_dfrbpq_1 _10230_ (.RESET_B(net923),
    .D(_00369_),
    .Q(\rf_ram.RAM[31][30] ),
    .CLK(clknet_leaf_163_clk_regs));
 sg13g2_dfrbpq_1 _10231_ (.RESET_B(net922),
    .D(_00370_),
    .Q(\rf_ram.RAM[31][31] ),
    .CLK(clknet_leaf_168_clk_regs));
 sg13g2_dfrbpq_1 _10232_ (.RESET_B(net921),
    .D(net3282),
    .Q(\rf_ram.RAM[29][0] ),
    .CLK(clknet_leaf_154_clk_regs));
 sg13g2_dfrbpq_1 _10233_ (.RESET_B(net920),
    .D(_00372_),
    .Q(\rf_ram.RAM[29][1] ),
    .CLK(clknet_leaf_52_clk_regs));
 sg13g2_dfrbpq_1 _10234_ (.RESET_B(net919),
    .D(_00373_),
    .Q(\rf_ram.RAM[29][2] ),
    .CLK(clknet_leaf_68_clk_regs));
 sg13g2_dfrbpq_1 _10235_ (.RESET_B(net918),
    .D(_00374_),
    .Q(\rf_ram.RAM[29][3] ),
    .CLK(clknet_leaf_86_clk_regs));
 sg13g2_dfrbpq_1 _10236_ (.RESET_B(net917),
    .D(_00375_),
    .Q(\rf_ram.RAM[29][4] ),
    .CLK(clknet_leaf_87_clk_regs));
 sg13g2_dfrbpq_1 _10237_ (.RESET_B(net916),
    .D(_00376_),
    .Q(\rf_ram.RAM[29][5] ),
    .CLK(clknet_leaf_92_clk_regs));
 sg13g2_dfrbpq_1 _10238_ (.RESET_B(net915),
    .D(_00377_),
    .Q(\rf_ram.RAM[29][6] ),
    .CLK(clknet_leaf_94_clk_regs));
 sg13g2_dfrbpq_1 _10239_ (.RESET_B(net914),
    .D(_00378_),
    .Q(\rf_ram.RAM[29][7] ),
    .CLK(clknet_leaf_95_clk_regs));
 sg13g2_dfrbpq_1 _10240_ (.RESET_B(net913),
    .D(_00379_),
    .Q(\rf_ram.RAM[29][8] ),
    .CLK(clknet_leaf_116_clk_regs));
 sg13g2_dfrbpq_1 _10241_ (.RESET_B(net912),
    .D(_00380_),
    .Q(\rf_ram.RAM[29][9] ),
    .CLK(clknet_leaf_124_clk_regs));
 sg13g2_dfrbpq_1 _10242_ (.RESET_B(net911),
    .D(_00381_),
    .Q(\rf_ram.RAM[29][10] ),
    .CLK(clknet_leaf_118_clk_regs));
 sg13g2_dfrbpq_1 _10243_ (.RESET_B(net910),
    .D(_00382_),
    .Q(\rf_ram.RAM[29][11] ),
    .CLK(clknet_leaf_135_clk_regs));
 sg13g2_dfrbpq_1 _10244_ (.RESET_B(net909),
    .D(_00383_),
    .Q(\rf_ram.RAM[29][12] ),
    .CLK(clknet_leaf_123_clk_regs));
 sg13g2_dfrbpq_1 _10245_ (.RESET_B(net908),
    .D(_00384_),
    .Q(\rf_ram.RAM[29][13] ),
    .CLK(clknet_leaf_90_clk_regs));
 sg13g2_dfrbpq_1 _10246_ (.RESET_B(net907),
    .D(_00385_),
    .Q(\rf_ram.RAM[29][14] ),
    .CLK(clknet_leaf_140_clk_regs));
 sg13g2_dfrbpq_1 _10247_ (.RESET_B(net906),
    .D(_00386_),
    .Q(\rf_ram.RAM[29][15] ),
    .CLK(clknet_leaf_109_clk_regs));
 sg13g2_dfrbpq_1 _10248_ (.RESET_B(net905),
    .D(_00387_),
    .Q(\rf_ram.RAM[29][16] ),
    .CLK(clknet_leaf_107_clk_regs));
 sg13g2_dfrbpq_1 _10249_ (.RESET_B(net904),
    .D(_00388_),
    .Q(\rf_ram.RAM[29][17] ),
    .CLK(clknet_leaf_139_clk_regs));
 sg13g2_dfrbpq_1 _10250_ (.RESET_B(net903),
    .D(_00389_),
    .Q(\rf_ram.RAM[29][18] ),
    .CLK(clknet_leaf_135_clk_regs));
 sg13g2_dfrbpq_1 _10251_ (.RESET_B(net902),
    .D(_00390_),
    .Q(\rf_ram.RAM[29][19] ),
    .CLK(clknet_leaf_155_clk_regs));
 sg13g2_dfrbpq_1 _10252_ (.RESET_B(net901),
    .D(_00391_),
    .Q(\rf_ram.RAM[29][20] ),
    .CLK(clknet_leaf_151_clk_regs));
 sg13g2_dfrbpq_1 _10253_ (.RESET_B(net900),
    .D(_00392_),
    .Q(\rf_ram.RAM[29][21] ),
    .CLK(clknet_leaf_65_clk_regs));
 sg13g2_dfrbpq_1 _10254_ (.RESET_B(net899),
    .D(_00393_),
    .Q(\rf_ram.RAM[29][22] ),
    .CLK(clknet_leaf_102_clk_regs));
 sg13g2_dfrbpq_1 _10255_ (.RESET_B(net898),
    .D(_00394_),
    .Q(\rf_ram.RAM[29][23] ),
    .CLK(clknet_leaf_59_clk_regs));
 sg13g2_dfrbpq_1 _10256_ (.RESET_B(net897),
    .D(_00395_),
    .Q(\rf_ram.RAM[29][24] ),
    .CLK(clknet_leaf_73_clk_regs));
 sg13g2_dfrbpq_1 _10257_ (.RESET_B(net896),
    .D(_00396_),
    .Q(\rf_ram.RAM[29][25] ),
    .CLK(clknet_leaf_50_clk_regs));
 sg13g2_dfrbpq_1 _10258_ (.RESET_B(net895),
    .D(_00397_),
    .Q(\rf_ram.RAM[29][26] ),
    .CLK(clknet_leaf_50_clk_regs));
 sg13g2_dfrbpq_1 _10259_ (.RESET_B(net894),
    .D(_00398_),
    .Q(\rf_ram.RAM[29][27] ),
    .CLK(clknet_leaf_43_clk_regs));
 sg13g2_dfrbpq_1 _10260_ (.RESET_B(net893),
    .D(_00399_),
    .Q(\rf_ram.RAM[29][28] ),
    .CLK(clknet_leaf_25_clk_regs));
 sg13g2_dfrbpq_1 _10261_ (.RESET_B(net892),
    .D(_00400_),
    .Q(\rf_ram.RAM[29][29] ),
    .CLK(clknet_leaf_154_clk_regs));
 sg13g2_dfrbpq_1 _10262_ (.RESET_B(net891),
    .D(_00401_),
    .Q(\rf_ram.RAM[29][30] ),
    .CLK(clknet_leaf_163_clk_regs));
 sg13g2_dfrbpq_1 _10263_ (.RESET_B(net890),
    .D(_00402_),
    .Q(\rf_ram.RAM[29][31] ),
    .CLK(clknet_leaf_168_clk_regs));
 sg13g2_dfrbpq_1 _10264_ (.RESET_B(net889),
    .D(net3393),
    .Q(\cpu.arbiter.i_wb_cpu_dbus_adr[2] ),
    .CLK(clknet_leaf_38_clk_regs));
 sg13g2_dfrbpq_1 _10265_ (.RESET_B(net888),
    .D(net3677),
    .Q(\cpu.arbiter.i_wb_cpu_dbus_adr[3] ),
    .CLK(clknet_leaf_38_clk_regs));
 sg13g2_dfrbpq_1 _10266_ (.RESET_B(net887),
    .D(_00405_),
    .Q(\cpu.arbiter.i_wb_cpu_dbus_adr[4] ),
    .CLK(clknet_leaf_39_clk_regs));
 sg13g2_dfrbpq_1 _10267_ (.RESET_B(net886),
    .D(_00406_),
    .Q(\cpu.arbiter.i_wb_cpu_dbus_adr[5] ),
    .CLK(clknet_leaf_39_clk_regs));
 sg13g2_dfrbpq_1 _10268_ (.RESET_B(net885),
    .D(net3655),
    .Q(\cpu.arbiter.i_wb_cpu_dbus_adr[6] ),
    .CLK(clknet_leaf_38_clk_regs));
 sg13g2_dfrbpq_1 _10269_ (.RESET_B(net884),
    .D(net3665),
    .Q(\cpu.arbiter.i_wb_cpu_dbus_adr[7] ),
    .CLK(clknet_leaf_37_clk_regs));
 sg13g2_dfrbpq_1 _10270_ (.RESET_B(net883),
    .D(_00409_),
    .Q(\cpu.arbiter.i_wb_cpu_dbus_adr[8] ),
    .CLK(clknet_leaf_37_clk_regs));
 sg13g2_dfrbpq_2 _10271_ (.RESET_B(net882),
    .D(_00410_),
    .Q(\cpu.arbiter.i_wb_cpu_dbus_adr[9] ),
    .CLK(clknet_leaf_30_clk_regs));
 sg13g2_dfrbpq_1 _10272_ (.RESET_B(net881),
    .D(net3663),
    .Q(\cpu.arbiter.i_wb_cpu_dbus_adr[10] ),
    .CLK(clknet_leaf_10_clk_regs));
 sg13g2_dfrbpq_1 _10273_ (.RESET_B(net880),
    .D(_00412_),
    .Q(\cpu.arbiter.i_wb_cpu_dbus_adr[11] ),
    .CLK(clknet_leaf_10_clk_regs));
 sg13g2_dfrbpq_1 _10274_ (.RESET_B(net879),
    .D(_00413_),
    .Q(\cpu.arbiter.i_wb_cpu_dbus_adr[12] ),
    .CLK(clknet_leaf_8_clk_regs));
 sg13g2_dfrbpq_1 _10275_ (.RESET_B(net878),
    .D(net3672),
    .Q(\cpu.arbiter.i_wb_cpu_dbus_adr[13] ),
    .CLK(clknet_leaf_8_clk_regs));
 sg13g2_dfrbpq_1 _10276_ (.RESET_B(net877),
    .D(_00415_),
    .Q(\cpu.arbiter.i_wb_cpu_dbus_adr[14] ),
    .CLK(clknet_leaf_8_clk_regs));
 sg13g2_dfrbpq_1 _10277_ (.RESET_B(net876),
    .D(net3529),
    .Q(\cpu.arbiter.i_wb_cpu_dbus_adr[15] ),
    .CLK(clknet_leaf_7_clk_regs));
 sg13g2_dfrbpq_1 _10278_ (.RESET_B(net875),
    .D(net3515),
    .Q(\cpu.arbiter.i_wb_cpu_dbus_adr[16] ),
    .CLK(clknet_leaf_7_clk_regs));
 sg13g2_dfrbpq_1 _10279_ (.RESET_B(net874),
    .D(_00418_),
    .Q(\cpu.arbiter.i_wb_cpu_dbus_adr[17] ),
    .CLK(clknet_leaf_2_clk_regs));
 sg13g2_dfrbpq_1 _10280_ (.RESET_B(net873),
    .D(_00419_),
    .Q(\cpu.arbiter.i_wb_cpu_dbus_adr[18] ),
    .CLK(clknet_leaf_2_clk_regs));
 sg13g2_dfrbpq_1 _10281_ (.RESET_B(net872),
    .D(_00420_),
    .Q(\cpu.arbiter.i_wb_cpu_dbus_adr[19] ),
    .CLK(clknet_leaf_2_clk_regs));
 sg13g2_dfrbpq_1 _10282_ (.RESET_B(net871),
    .D(_00421_),
    .Q(\cpu.arbiter.i_wb_cpu_dbus_adr[20] ),
    .CLK(clknet_leaf_7_clk_regs));
 sg13g2_dfrbpq_1 _10283_ (.RESET_B(net870),
    .D(_00422_),
    .Q(\cpu.arbiter.i_wb_cpu_dbus_adr[21] ),
    .CLK(clknet_leaf_0_clk_regs));
 sg13g2_dfrbpq_1 _10284_ (.RESET_B(net869),
    .D(net3562),
    .Q(\cpu.arbiter.i_wb_cpu_dbus_adr[22] ),
    .CLK(clknet_leaf_171_clk_regs));
 sg13g2_dfrbpq_1 _10285_ (.RESET_B(net868),
    .D(net3507),
    .Q(\cpu.arbiter.i_wb_cpu_dbus_adr[23] ),
    .CLK(clknet_leaf_171_clk_regs));
 sg13g2_dfrbpq_1 _10286_ (.RESET_B(net867),
    .D(_00425_),
    .Q(\cpu.arbiter.i_wb_cpu_dbus_adr[24] ),
    .CLK(clknet_leaf_171_clk_regs));
 sg13g2_dfrbpq_1 _10287_ (.RESET_B(net866),
    .D(_00426_),
    .Q(\cpu.arbiter.i_wb_cpu_dbus_adr[25] ),
    .CLK(clknet_leaf_171_clk_regs));
 sg13g2_dfrbpq_1 _10288_ (.RESET_B(net865),
    .D(_00427_),
    .Q(\cpu.arbiter.i_wb_cpu_dbus_adr[26] ),
    .CLK(clknet_leaf_171_clk_regs));
 sg13g2_dfrbpq_1 _10289_ (.RESET_B(net864),
    .D(net3555),
    .Q(\cpu.arbiter.i_wb_cpu_dbus_adr[27] ),
    .CLK(clknet_leaf_171_clk_regs));
 sg13g2_dfrbpq_1 _10290_ (.RESET_B(net863),
    .D(net3509),
    .Q(\cpu.arbiter.i_wb_cpu_dbus_adr[28] ),
    .CLK(clknet_leaf_171_clk_regs));
 sg13g2_dfrbpq_1 _10291_ (.RESET_B(net862),
    .D(_00430_),
    .Q(\cpu.arbiter.i_wb_cpu_dbus_adr[29] ),
    .CLK(clknet_leaf_172_clk_regs));
 sg13g2_dfrbpq_2 _10292_ (.RESET_B(net861),
    .D(_00431_),
    .Q(\cpu.arbiter.i_wb_cpu_dbus_adr[30] ),
    .CLK(clknet_leaf_39_clk_regs));
 sg13g2_dfrbpq_2 _10293_ (.RESET_B(net1089),
    .D(net3745),
    .Q(\cpu.arbiter.i_wb_cpu_dbus_adr[31] ),
    .CLK(clknet_leaf_33_clk_regs));
 sg13g2_dfrbpq_2 _10294_ (.RESET_B(net1090),
    .D(net3647),
    .Q(\cpu.rf_ram_if.rdata1[0] ),
    .CLK(clknet_leaf_63_clk_regs));
 sg13g2_dfrbpq_1 _10295_ (.RESET_B(net1091),
    .D(_00042_),
    .Q(\cpu.rf_ram_if.rdata1[1] ),
    .CLK(clknet_leaf_104_clk_regs));
 sg13g2_dfrbpq_1 _10296_ (.RESET_B(net1092),
    .D(net3539),
    .Q(\cpu.rf_ram_if.rdata1[2] ),
    .CLK(clknet_leaf_98_clk_regs));
 sg13g2_dfrbpq_1 _10297_ (.RESET_B(net1093),
    .D(net3358),
    .Q(\cpu.rf_ram_if.rdata1[3] ),
    .CLK(clknet_leaf_96_clk_regs));
 sg13g2_dfrbpq_1 _10298_ (.RESET_B(net1094),
    .D(net3409),
    .Q(\cpu.rf_ram_if.rdata1[4] ),
    .CLK(clknet_leaf_97_clk_regs));
 sg13g2_dfrbpq_1 _10299_ (.RESET_B(net1095),
    .D(net3366),
    .Q(\cpu.rf_ram_if.rdata1[5] ),
    .CLK(clknet_leaf_97_clk_regs));
 sg13g2_dfrbpq_1 _10300_ (.RESET_B(net1096),
    .D(net3445),
    .Q(\cpu.rf_ram_if.rdata1[6] ),
    .CLK(clknet_leaf_97_clk_regs));
 sg13g2_dfrbpq_1 _10301_ (.RESET_B(net1097),
    .D(net3483),
    .Q(\cpu.rf_ram_if.rdata1[7] ),
    .CLK(clknet_leaf_97_clk_regs));
 sg13g2_dfrbpq_1 _10302_ (.RESET_B(net1098),
    .D(net3471),
    .Q(\cpu.rf_ram_if.rdata1[8] ),
    .CLK(clknet_leaf_114_clk_regs));
 sg13g2_dfrbpq_1 _10303_ (.RESET_B(net1099),
    .D(net3356),
    .Q(\cpu.rf_ram_if.rdata1[9] ),
    .CLK(clknet_leaf_119_clk_regs));
 sg13g2_dfrbpq_1 _10304_ (.RESET_B(net1100),
    .D(net3379),
    .Q(\cpu.rf_ram_if.rdata1[10] ),
    .CLK(clknet_leaf_120_clk_regs));
 sg13g2_dfrbpq_1 _10305_ (.RESET_B(net1101),
    .D(net3431),
    .Q(\cpu.rf_ram_if.rdata1[11] ),
    .CLK(clknet_leaf_111_clk_regs));
 sg13g2_dfrbpq_1 _10306_ (.RESET_B(net1102),
    .D(net3352),
    .Q(\cpu.rf_ram_if.rdata1[12] ),
    .CLK(clknet_leaf_111_clk_regs));
 sg13g2_dfrbpq_1 _10307_ (.RESET_B(net1103),
    .D(net3524),
    .Q(\cpu.rf_ram_if.rdata1[13] ),
    .CLK(clknet_leaf_110_clk_regs));
 sg13g2_dfrbpq_1 _10308_ (.RESET_B(net1104),
    .D(net3397),
    .Q(\cpu.rf_ram_if.rdata1[14] ),
    .CLK(clknet_leaf_145_clk_regs));
 sg13g2_dfrbpq_1 _10309_ (.RESET_B(net1105),
    .D(net3354),
    .Q(\cpu.rf_ram_if.rdata1[15] ),
    .CLK(clknet_leaf_145_clk_regs));
 sg13g2_dfrbpq_1 _10310_ (.RESET_B(net1106),
    .D(net3370),
    .Q(\cpu.rf_ram_if.rdata1[16] ),
    .CLK(clknet_leaf_145_clk_regs));
 sg13g2_dfrbpq_1 _10311_ (.RESET_B(net1107),
    .D(net3339),
    .Q(\cpu.rf_ram_if.rdata1[17] ),
    .CLK(clknet_leaf_145_clk_regs));
 sg13g2_dfrbpq_1 _10312_ (.RESET_B(net1108),
    .D(net3513),
    .Q(\cpu.rf_ram_if.rdata1[18] ),
    .CLK(clknet_leaf_146_clk_regs));
 sg13g2_dfrbpq_1 _10313_ (.RESET_B(net1109),
    .D(net3503),
    .Q(\cpu.rf_ram_if.rdata1[19] ),
    .CLK(clknet_leaf_149_clk_regs));
 sg13g2_dfrbpq_1 _10314_ (.RESET_B(net1110),
    .D(net3305),
    .Q(\cpu.rf_ram_if.rdata1[20] ),
    .CLK(clknet_leaf_63_clk_regs));
 sg13g2_dfrbpq_1 _10315_ (.RESET_B(net1111),
    .D(net3402),
    .Q(\cpu.rf_ram_if.rdata1[21] ),
    .CLK(clknet_leaf_62_clk_regs));
 sg13g2_dfrbpq_1 _10316_ (.RESET_B(net1112),
    .D(net3605),
    .Q(\cpu.rf_ram_if.rdata1[22] ),
    .CLK(clknet_leaf_21_clk_regs));
 sg13g2_dfrbpq_1 _10317_ (.RESET_B(net1113),
    .D(net3372),
    .Q(\cpu.rf_ram_if.rdata1[23] ),
    .CLK(clknet_leaf_23_clk_regs));
 sg13g2_dfrbpq_1 _10318_ (.RESET_B(net1114),
    .D(net3406),
    .Q(\cpu.rf_ram_if.rdata1[24] ),
    .CLK(clknet_leaf_23_clk_regs));
 sg13g2_dfrbpq_1 _10319_ (.RESET_B(net1115),
    .D(net3447),
    .Q(\cpu.rf_ram_if.rdata1[25] ),
    .CLK(clknet_leaf_23_clk_regs));
 sg13g2_dfrbpq_1 _10320_ (.RESET_B(net1116),
    .D(net3469),
    .Q(\cpu.rf_ram_if.rdata1[26] ),
    .CLK(clknet_leaf_18_clk_regs));
 sg13g2_dfrbpq_1 _10321_ (.RESET_B(net1117),
    .D(net3425),
    .Q(\cpu.rf_ram_if.rdata1[27] ),
    .CLK(clknet_leaf_13_clk_regs));
 sg13g2_dfrbpq_1 _10322_ (.RESET_B(net1118),
    .D(net3413),
    .Q(\cpu.rf_ram_if.rdata1[28] ),
    .CLK(clknet_leaf_13_clk_regs));
 sg13g2_dfrbpq_1 _10323_ (.RESET_B(net1119),
    .D(net3415),
    .Q(\cpu.rf_ram_if.rdata1[29] ),
    .CLK(clknet_leaf_13_clk_regs));
 sg13g2_dfrbpq_2 _10324_ (.RESET_B(net1120),
    .D(net3645),
    .Q(\cpu.cpu.alu.i_rs1 [0]),
    .CLK(clknet_leaf_29_clk_regs));
 sg13g2_dfrbpq_2 _10325_ (.RESET_B(net1121),
    .D(net3657),
    .Q(\cpu.rf_ram_if.rdata0[1] ),
    .CLK(clknet_leaf_63_clk_regs));
 sg13g2_dfrbpq_1 _10326_ (.RESET_B(net1122),
    .D(net3575),
    .Q(\cpu.rf_ram_if.rdata0[2] ),
    .CLK(clknet_leaf_103_clk_regs));
 sg13g2_dfrbpq_1 _10327_ (.RESET_B(net1123),
    .D(net3499),
    .Q(\cpu.rf_ram_if.rdata0[3] ),
    .CLK(clknet_leaf_98_clk_regs));
 sg13g2_dfrbpq_1 _10328_ (.RESET_B(net1124),
    .D(net3360),
    .Q(\cpu.rf_ram_if.rdata0[4] ),
    .CLK(clknet_leaf_97_clk_regs));
 sg13g2_dfrbpq_1 _10329_ (.RESET_B(net1125),
    .D(net3376),
    .Q(\cpu.rf_ram_if.rdata0[5] ),
    .CLK(clknet_leaf_97_clk_regs));
 sg13g2_dfrbpq_1 _10330_ (.RESET_B(net1126),
    .D(net3328),
    .Q(\cpu.rf_ram_if.rdata0[6] ),
    .CLK(clknet_leaf_97_clk_regs));
 sg13g2_dfrbpq_1 _10331_ (.RESET_B(net1127),
    .D(net3505),
    .Q(\cpu.rf_ram_if.rdata0[7] ),
    .CLK(clknet_leaf_113_clk_regs));
 sg13g2_dfrbpq_1 _10332_ (.RESET_B(net1128),
    .D(net3453),
    .Q(\cpu.rf_ram_if.rdata0[8] ),
    .CLK(clknet_leaf_115_clk_regs));
 sg13g2_dfrbpq_1 _10333_ (.RESET_B(net1129),
    .D(net3423),
    .Q(\cpu.rf_ram_if.rdata0[9] ),
    .CLK(clknet_leaf_114_clk_regs));
 sg13g2_dfrbpq_1 _10334_ (.RESET_B(net1130),
    .D(net3395),
    .Q(\cpu.rf_ram_if.rdata0[10] ),
    .CLK(clknet_leaf_119_clk_regs));
 sg13g2_dfrbpq_1 _10335_ (.RESET_B(net1131),
    .D(net3449),
    .Q(\cpu.rf_ram_if.rdata0[11] ),
    .CLK(clknet_leaf_120_clk_regs));
 sg13g2_dfrbpq_1 _10336_ (.RESET_B(net1132),
    .D(net3417),
    .Q(\cpu.rf_ram_if.rdata0[12] ),
    .CLK(clknet_leaf_111_clk_regs));
 sg13g2_dfrbpq_1 _10337_ (.RESET_B(net1133),
    .D(net3331),
    .Q(\cpu.rf_ram_if.rdata0[13] ),
    .CLK(clknet_leaf_111_clk_regs));
 sg13g2_dfrbpq_1 _10338_ (.RESET_B(net1134),
    .D(net3531),
    .Q(\cpu.rf_ram_if.rdata0[14] ),
    .CLK(clknet_leaf_110_clk_regs));
 sg13g2_dfrbpq_1 _10339_ (.RESET_B(net1135),
    .D(net3467),
    .Q(\cpu.rf_ram_if.rdata0[15] ),
    .CLK(clknet_leaf_145_clk_regs));
 sg13g2_dfrbpq_1 _10340_ (.RESET_B(net1136),
    .D(net3385),
    .Q(\cpu.rf_ram_if.rdata0[16] ),
    .CLK(clknet_leaf_146_clk_regs));
 sg13g2_dfrbpq_1 _10341_ (.RESET_B(net1137),
    .D(net3348),
    .Q(\cpu.rf_ram_if.rdata0[17] ),
    .CLK(clknet_leaf_146_clk_regs));
 sg13g2_dfrbpq_1 _10342_ (.RESET_B(net1138),
    .D(net3350),
    .Q(\cpu.rf_ram_if.rdata0[18] ),
    .CLK(clknet_leaf_146_clk_regs));
 sg13g2_dfrbpq_1 _10343_ (.RESET_B(net1139),
    .D(net3526),
    .Q(\cpu.rf_ram_if.rdata0[19] ),
    .CLK(clknet_leaf_146_clk_regs));
 sg13g2_dfrbpq_1 _10344_ (.RESET_B(net1140),
    .D(net1405),
    .Q(\cpu.rf_ram_if.rdata0[20] ),
    .CLK(clknet_leaf_149_clk_regs));
 sg13g2_dfrbpq_1 _10345_ (.RESET_B(net1141),
    .D(net3761),
    .Q(\cpu.rf_ram_if.rdata0[21] ),
    .CLK(clknet_5_18__leaf_clk_regs));
 sg13g2_dfrbpq_1 _10346_ (.RESET_B(net1142),
    .D(net3428),
    .Q(\cpu.rf_ram_if.rdata0[22] ),
    .CLK(clknet_leaf_62_clk_regs));
 sg13g2_dfrbpq_1 _10347_ (.RESET_B(net1143),
    .D(net3573),
    .Q(\cpu.rf_ram_if.rdata0[23] ),
    .CLK(clknet_leaf_21_clk_regs));
 sg13g2_dfrbpq_1 _10348_ (.RESET_B(net1144),
    .D(net3333),
    .Q(\cpu.rf_ram_if.rdata0[24] ),
    .CLK(clknet_leaf_23_clk_regs));
 sg13g2_dfrbpq_1 _10349_ (.RESET_B(net1145),
    .D(net3411),
    .Q(\cpu.rf_ram_if.rdata0[25] ),
    .CLK(clknet_leaf_23_clk_regs));
 sg13g2_dfrbpq_1 _10350_ (.RESET_B(net1146),
    .D(net3460),
    .Q(\cpu.rf_ram_if.rdata0[26] ),
    .CLK(clknet_leaf_23_clk_regs));
 sg13g2_dfrbpq_1 _10351_ (.RESET_B(net1147),
    .D(net3443),
    .Q(\cpu.rf_ram_if.rdata0[27] ),
    .CLK(clknet_leaf_18_clk_regs));
 sg13g2_dfrbpq_1 _10352_ (.RESET_B(net1148),
    .D(net3346),
    .Q(\cpu.rf_ram_if.rdata0[28] ),
    .CLK(clknet_leaf_13_clk_regs));
 sg13g2_dfrbpq_1 _10353_ (.RESET_B(net1182),
    .D(net3390),
    .Q(\cpu.rf_ram_if.rdata0[29] ),
    .CLK(clknet_leaf_13_clk_regs));
 sg13g2_dfrbpq_1 _10354_ (.RESET_B(net860),
    .D(net3404),
    .Q(\cpu.rf_ram_if.rdata0[30] ),
    .CLK(clknet_leaf_13_clk_regs));
 sg13g2_dfrbpq_1 _10355_ (.RESET_B(net859),
    .D(_00433_),
    .Q(\cpu.i_rf_rdata[0] ),
    .CLK(clknet_leaf_18_clk_regs));
 sg13g2_dfrbpq_1 _10356_ (.RESET_B(net858),
    .D(_00434_),
    .Q(\cpu.i_rf_rdata[1] ),
    .CLK(clknet_leaf_71_clk_regs));
 sg13g2_dfrbpq_1 _10357_ (.RESET_B(net857),
    .D(_00435_),
    .Q(\cpu.i_rf_rdata[2] ),
    .CLK(clknet_leaf_104_clk_regs));
 sg13g2_dfrbpq_1 _10358_ (.RESET_B(net856),
    .D(net3797),
    .Q(\cpu.i_rf_rdata[3] ),
    .CLK(clknet_leaf_91_clk_regs));
 sg13g2_dfrbpq_1 _10359_ (.RESET_B(net855),
    .D(net3787),
    .Q(\cpu.i_rf_rdata[4] ),
    .CLK(clknet_leaf_91_clk_regs));
 sg13g2_dfrbpq_1 _10360_ (.RESET_B(net854),
    .D(_00438_),
    .Q(\cpu.i_rf_rdata[5] ),
    .CLK(clknet_leaf_100_clk_regs));
 sg13g2_dfrbpq_1 _10361_ (.RESET_B(net853),
    .D(_00439_),
    .Q(\cpu.i_rf_rdata[6] ),
    .CLK(clknet_leaf_100_clk_regs));
 sg13g2_dfrbpq_1 _10362_ (.RESET_B(net852),
    .D(_00440_),
    .Q(\cpu.i_rf_rdata[7] ),
    .CLK(clknet_leaf_97_clk_regs));
 sg13g2_dfrbpq_1 _10363_ (.RESET_B(net851),
    .D(_00441_),
    .Q(\cpu.i_rf_rdata[8] ),
    .CLK(clknet_leaf_115_clk_regs));
 sg13g2_dfrbpq_1 _10364_ (.RESET_B(net850),
    .D(net3802),
    .Q(\cpu.i_rf_rdata[9] ),
    .CLK(clknet_leaf_111_clk_regs));
 sg13g2_dfrbpq_1 _10365_ (.RESET_B(net849),
    .D(_00443_),
    .Q(\cpu.i_rf_rdata[10] ),
    .CLK(clknet_leaf_119_clk_regs));
 sg13g2_dfrbpq_1 _10366_ (.RESET_B(net848),
    .D(_00444_),
    .Q(\cpu.i_rf_rdata[11] ),
    .CLK(clknet_leaf_131_clk_regs));
 sg13g2_dfrbpq_1 _10367_ (.RESET_B(net847),
    .D(_00445_),
    .Q(\cpu.i_rf_rdata[12] ),
    .CLK(clknet_leaf_121_clk_regs));
 sg13g2_dfrbpq_1 _10368_ (.RESET_B(net846),
    .D(_00446_),
    .Q(\cpu.i_rf_rdata[13] ),
    .CLK(clknet_leaf_110_clk_regs));
 sg13g2_dfrbpq_1 _10369_ (.RESET_B(net845),
    .D(_00447_),
    .Q(\cpu.i_rf_rdata[14] ),
    .CLK(clknet_leaf_143_clk_regs));
 sg13g2_dfrbpq_1 _10370_ (.RESET_B(net844),
    .D(_00448_),
    .Q(\cpu.i_rf_rdata[15] ),
    .CLK(clknet_leaf_145_clk_regs));
 sg13g2_dfrbpq_1 _10371_ (.RESET_B(net843),
    .D(net3784),
    .Q(\cpu.i_rf_rdata[16] ),
    .CLK(clknet_leaf_107_clk_regs));
 sg13g2_dfrbpq_1 _10372_ (.RESET_B(net842),
    .D(_00450_),
    .Q(\cpu.i_rf_rdata[17] ),
    .CLK(clknet_leaf_141_clk_regs));
 sg13g2_dfrbpq_1 _10373_ (.RESET_B(net841),
    .D(net3792),
    .Q(\cpu.i_rf_rdata[18] ),
    .CLK(clknet_leaf_146_clk_regs));
 sg13g2_dfrbpq_1 _10374_ (.RESET_B(net840),
    .D(net3809),
    .Q(\cpu.i_rf_rdata[19] ),
    .CLK(clknet_leaf_146_clk_regs));
 sg13g2_dfrbpq_1 _10375_ (.RESET_B(net839),
    .D(_00453_),
    .Q(\cpu.i_rf_rdata[20] ),
    .CLK(clknet_leaf_149_clk_regs));
 sg13g2_dfrbpq_1 _10376_ (.RESET_B(net838),
    .D(_00454_),
    .Q(\cpu.i_rf_rdata[21] ),
    .CLK(clknet_leaf_63_clk_regs));
 sg13g2_dfrbpq_1 _10377_ (.RESET_B(net837),
    .D(_00455_),
    .Q(\cpu.i_rf_rdata[22] ),
    .CLK(clknet_leaf_63_clk_regs));
 sg13g2_dfrbpq_1 _10378_ (.RESET_B(net836),
    .D(_00456_),
    .Q(\cpu.i_rf_rdata[23] ),
    .CLK(clknet_leaf_19_clk_regs));
 sg13g2_dfrbpq_2 _10379_ (.RESET_B(net835),
    .D(_00457_),
    .Q(\cpu.i_rf_rdata[24] ),
    .CLK(clknet_leaf_71_clk_regs));
 sg13g2_dfrbpq_2 _10380_ (.RESET_B(net834),
    .D(_00458_),
    .Q(\cpu.i_rf_rdata[25] ),
    .CLK(clknet_leaf_47_clk_regs));
 sg13g2_dfrbpq_1 _10381_ (.RESET_B(net833),
    .D(net3795),
    .Q(\cpu.i_rf_rdata[26] ),
    .CLK(clknet_leaf_24_clk_regs));
 sg13g2_dfrbpq_2 _10382_ (.RESET_B(net832),
    .D(_00460_),
    .Q(\cpu.i_rf_rdata[27] ),
    .CLK(clknet_leaf_45_clk_regs));
 sg13g2_dfrbpq_1 _10383_ (.RESET_B(net831),
    .D(_00461_),
    .Q(\cpu.i_rf_rdata[28] ),
    .CLK(clknet_leaf_28_clk_regs));
 sg13g2_dfrbpq_1 _10384_ (.RESET_B(net830),
    .D(_00462_),
    .Q(\cpu.i_rf_rdata[29] ),
    .CLK(clknet_leaf_15_clk_regs));
 sg13g2_dfrbpq_1 _10385_ (.RESET_B(net829),
    .D(_00463_),
    .Q(\cpu.i_rf_rdata[30] ),
    .CLK(clknet_leaf_15_clk_regs));
 sg13g2_dfrbpq_1 _10386_ (.RESET_B(net828),
    .D(net3806),
    .Q(\cpu.i_rf_rdata[31] ),
    .CLK(clknet_leaf_14_clk_regs));
 sg13g2_dfrbpq_1 _10387_ (.RESET_B(net1186),
    .D(_00465_),
    .Q(\cpu.cpu.state.ibus_cyc ),
    .CLK(clknet_leaf_33_clk_regs));
 sg13g2_dfrbpq_1 _10388_ (.RESET_B(net827),
    .D(net2583),
    .Q(\cpu.rf_ram_if.gen_wtrig_ratio_neq_2.wtrig0_r ),
    .CLK(clknet_leaf_22_clk_regs));
 sg13g2_dfrbpq_1 _10389_ (.RESET_B(net826),
    .D(_00466_),
    .Q(\cpu.rf_ram_if.rdata1[30] ),
    .CLK(clknet_leaf_14_clk_regs));
 sg13g2_dfrbpq_1 _10390_ (.RESET_B(net825),
    .D(_00467_),
    .Q(\cpu.rf_ram_if.rdata0[31] ),
    .CLK(clknet_leaf_14_clk_regs));
 sg13g2_dfrbpq_1 _10391_ (.RESET_B(net1189),
    .D(_00468_),
    .Q(\cpu.rf_ram_if.rgnt ),
    .CLK(clknet_leaf_31_clk_regs));
 sg13g2_dfrbpq_2 _10392_ (.RESET_B(net824),
    .D(\cpu.rf_ram_if.rtrig0 ),
    .Q(\cpu.rf_ram_if.rtrig1 ),
    .CLK(clknet_leaf_28_clk_regs));
 sg13g2_dfrbpq_1 _10393_ (.RESET_B(net823),
    .D(_00469_),
    .Q(\cpu.rf_ram_if.rgate ),
    .CLK(clknet_leaf_36_clk_regs));
 sg13g2_dfrbpq_2 _10394_ (.RESET_B(net1190),
    .D(_00470_),
    .Q(\cpu.rf_ram_if.rcnt[1] ),
    .CLK(clknet_leaf_35_clk_regs));
 sg13g2_dfrbpq_1 _10395_ (.RESET_B(net1191),
    .D(net1410),
    .Q(\cpu.rf_ram_if.wdata0_r[0] ),
    .CLK(clknet_leaf_22_clk_regs));
 sg13g2_dfrbpq_2 _10396_ (.RESET_B(net1192),
    .D(net1412),
    .Q(\cpu.rf_ram_if.wdata0_r[1] ),
    .CLK(clknet_leaf_71_clk_regs));
 sg13g2_dfrbpq_2 _10397_ (.RESET_B(net1193),
    .D(net1387),
    .Q(\cpu.rf_ram_if.wdata0_r[2] ),
    .CLK(clknet_leaf_80_clk_regs));
 sg13g2_dfrbpq_1 _10398_ (.RESET_B(net1194),
    .D(net1400),
    .Q(\cpu.rf_ram_if.wdata0_r[3] ),
    .CLK(clknet_leaf_80_clk_regs));
 sg13g2_dfrbpq_1 _10399_ (.RESET_B(net1195),
    .D(net1393),
    .Q(\cpu.rf_ram_if.wdata0_r[4] ),
    .CLK(clknet_leaf_81_clk_regs));
 sg13g2_dfrbpq_1 _10400_ (.RESET_B(net1196),
    .D(net1408),
    .Q(\cpu.rf_ram_if.wdata0_r[5] ),
    .CLK(clknet_leaf_81_clk_regs));
 sg13g2_dfrbpq_1 _10401_ (.RESET_B(net1197),
    .D(net1397),
    .Q(\cpu.rf_ram_if.wdata0_r[6] ),
    .CLK(clknet_leaf_99_clk_regs));
 sg13g2_dfrbpq_1 _10402_ (.RESET_B(net1198),
    .D(net1402),
    .Q(\cpu.rf_ram_if.wdata0_r[7] ),
    .CLK(clknet_leaf_99_clk_regs));
 sg13g2_dfrbpq_1 _10403_ (.RESET_B(net1199),
    .D(net1409),
    .Q(\cpu.rf_ram_if.wdata0_r[8] ),
    .CLK(clknet_leaf_114_clk_regs));
 sg13g2_dfrbpq_1 _10404_ (.RESET_B(net1200),
    .D(net1392),
    .Q(\cpu.rf_ram_if.wdata0_r[9] ),
    .CLK(clknet_leaf_121_clk_regs));
 sg13g2_dfrbpq_1 _10405_ (.RESET_B(net1201),
    .D(net1381),
    .Q(\cpu.rf_ram_if.wdata0_r[10] ),
    .CLK(clknet_leaf_121_clk_regs));
 sg13g2_dfrbpq_1 _10406_ (.RESET_B(net1202),
    .D(net1401),
    .Q(\cpu.rf_ram_if.wdata0_r[11] ),
    .CLK(clknet_leaf_132_clk_regs));
 sg13g2_dfrbpq_1 _10407_ (.RESET_B(net1203),
    .D(net1396),
    .Q(\cpu.rf_ram_if.wdata0_r[12] ),
    .CLK(clknet_leaf_132_clk_regs));
 sg13g2_dfrbpq_1 _10408_ (.RESET_B(net1204),
    .D(net1389),
    .Q(\cpu.rf_ram_if.wdata0_r[13] ),
    .CLK(clknet_leaf_143_clk_regs));
 sg13g2_dfrbpq_1 _10409_ (.RESET_B(net1205),
    .D(net1385),
    .Q(\cpu.rf_ram_if.wdata0_r[14] ),
    .CLK(clknet_leaf_142_clk_regs));
 sg13g2_dfrbpq_1 _10410_ (.RESET_B(net1206),
    .D(net1394),
    .Q(\cpu.rf_ram_if.wdata0_r[15] ),
    .CLK(clknet_leaf_141_clk_regs));
 sg13g2_dfrbpq_1 _10411_ (.RESET_B(net1207),
    .D(net1398),
    .Q(\cpu.rf_ram_if.wdata0_r[16] ),
    .CLK(clknet_leaf_141_clk_regs));
 sg13g2_dfrbpq_1 _10412_ (.RESET_B(net1208),
    .D(net1388),
    .Q(\cpu.rf_ram_if.wdata0_r[17] ),
    .CLK(clknet_leaf_141_clk_regs));
 sg13g2_dfrbpq_1 _10413_ (.RESET_B(net1209),
    .D(net1390),
    .Q(\cpu.rf_ram_if.wdata0_r[18] ),
    .CLK(clknet_leaf_141_clk_regs));
 sg13g2_dfrbpq_1 _10414_ (.RESET_B(net1210),
    .D(net1413),
    .Q(\cpu.rf_ram_if.wdata0_r[19] ),
    .CLK(clknet_leaf_146_clk_regs));
 sg13g2_dfrbpq_2 _10415_ (.RESET_B(net1211),
    .D(net1403),
    .Q(\cpu.rf_ram_if.wdata0_r[20] ),
    .CLK(clknet_leaf_64_clk_regs));
 sg13g2_dfrbpq_1 _10416_ (.RESET_B(net1212),
    .D(net1383),
    .Q(\cpu.rf_ram_if.wdata0_r[21] ),
    .CLK(clknet_leaf_65_clk_regs));
 sg13g2_dfrbpq_1 _10417_ (.RESET_B(net1213),
    .D(net1399),
    .Q(\cpu.rf_ram_if.wdata0_r[22] ),
    .CLK(clknet_leaf_65_clk_regs));
 sg13g2_dfrbpq_1 _10418_ (.RESET_B(net1214),
    .D(net1391),
    .Q(\cpu.rf_ram_if.wdata0_r[23] ),
    .CLK(clknet_leaf_65_clk_regs));
 sg13g2_dfrbpq_1 _10419_ (.RESET_B(net1215),
    .D(net1407),
    .Q(\cpu.rf_ram_if.wdata0_r[24] ),
    .CLK(clknet_leaf_65_clk_regs));
 sg13g2_dfrbpq_1 _10420_ (.RESET_B(net1216),
    .D(net1411),
    .Q(\cpu.rf_ram_if.wdata0_r[25] ),
    .CLK(clknet_leaf_58_clk_regs));
 sg13g2_dfrbpq_1 _10421_ (.RESET_B(net1217),
    .D(net1382),
    .Q(\cpu.rf_ram_if.wdata0_r[26] ),
    .CLK(clknet_leaf_35_clk_regs));
 sg13g2_dfrbpq_1 _10422_ (.RESET_B(net1218),
    .D(net1406),
    .Q(\cpu.rf_ram_if.wdata0_r[27] ),
    .CLK(clknet_leaf_35_clk_regs));
 sg13g2_dfrbpq_2 _10423_ (.RESET_B(net1219),
    .D(net1395),
    .Q(\cpu.rf_ram_if.wdata0_r[28] ),
    .CLK(clknet_leaf_15_clk_regs));
 sg13g2_dfrbpq_1 _10424_ (.RESET_B(net1220),
    .D(net1386),
    .Q(\cpu.rf_ram_if.wdata0_r[29] ),
    .CLK(clknet_leaf_15_clk_regs));
 sg13g2_dfrbpq_1 _10425_ (.RESET_B(net1290),
    .D(net1384),
    .Q(\cpu.rf_ram_if.wdata0_r[30] ),
    .CLK(clknet_leaf_6_clk_regs));
 sg13g2_dfrbpq_1 _10426_ (.RESET_B(net821),
    .D(\cpu.cpu.o_wdata0 [0]),
    .Q(\cpu.rf_ram_if.wdata0_r[31] ),
    .CLK(clknet_leaf_6_clk_regs));
 sg13g2_dfrbpq_1 _10427_ (.RESET_B(net820),
    .D(net2350),
    .Q(\cpu.rf_ram_if.rreq_r ),
    .CLK(clknet_leaf_31_clk_regs));
 sg13g2_dfrbpq_2 _10428_ (.RESET_B(net819),
    .D(net3607),
    .Q(\cpu.rf_ram_if.wen0_r ),
    .CLK(clknet_leaf_34_clk_regs));
 sg13g2_dfrbpq_1 _10429_ (.RESET_B(net818),
    .D(net2995),
    .Q(\cpu.cpu.mem_if.signbit ),
    .CLK(clknet_leaf_34_clk_regs));
 sg13g2_dfrbpq_2 _10430_ (.RESET_B(net817),
    .D(net3493),
    .Q(\cpu.cpu.state.o_cnt[2] ),
    .CLK(clknet_leaf_31_clk_regs));
 sg13g2_dfrbpq_2 _10431_ (.RESET_B(net816),
    .D(net3699),
    .Q(\cpu.cpu.bufreg2.i_bytecnt[0] ),
    .CLK(clknet_leaf_32_clk_regs));
 sg13g2_dfrbpq_2 _10432_ (.RESET_B(net815),
    .D(net3758),
    .Q(\cpu.cpu.bufreg2.i_bytecnt[1] ),
    .CLK(clknet_leaf_32_clk_regs));
 sg13g2_dfrbpq_1 _10433_ (.RESET_B(net814),
    .D(_00477_),
    .Q(\cpu.cpu.ctrl.i_jump ),
    .CLK(clknet_leaf_32_clk_regs));
 sg13g2_dfrbpq_2 _10434_ (.RESET_B(net812),
    .D(_00478_),
    .Q(\cpu.cpu.state.init_done ),
    .CLK(clknet_leaf_32_clk_regs));
 sg13g2_dfrbpq_2 _10435_ (.RESET_B(net810),
    .D(_00479_),
    .Q(\cpu.cpu.state.cnt_r[0] ),
    .CLK(clknet_leaf_31_clk_regs));
 sg13g2_dfrbpq_2 _10436_ (.RESET_B(net809),
    .D(_00480_),
    .Q(\cpu.cpu.state.cnt_r[1] ),
    .CLK(clknet_leaf_31_clk_regs));
 sg13g2_dfrbpq_2 _10437_ (.RESET_B(net808),
    .D(_00481_),
    .Q(\cpu.cpu.state.cnt_r[2] ),
    .CLK(clknet_leaf_31_clk_regs));
 sg13g2_dfrbpq_2 _10438_ (.RESET_B(net807),
    .D(_00482_),
    .Q(\cpu.cpu.state.cnt_r[3] ),
    .CLK(clknet_leaf_31_clk_regs));
 sg13g2_dfrbpq_2 _10439_ (.RESET_B(net806),
    .D(_00483_),
    .Q(\cpu.arbiter.i_wb_cpu_dbus_dat[0] ),
    .CLK(clknet_leaf_40_clk_regs));
 sg13g2_dfrbpq_2 _10440_ (.RESET_B(net805),
    .D(_00484_),
    .Q(\cpu.arbiter.i_wb_cpu_dbus_dat[1] ),
    .CLK(clknet_leaf_41_clk_regs));
 sg13g2_dfrbpq_2 _10441_ (.RESET_B(net804),
    .D(net3577),
    .Q(\cpu.arbiter.i_wb_cpu_dbus_dat[2] ),
    .CLK(clknet_leaf_41_clk_regs));
 sg13g2_dfrbpq_2 _10442_ (.RESET_B(net803),
    .D(_00486_),
    .Q(\cpu.arbiter.i_wb_cpu_dbus_dat[3] ),
    .CLK(clknet_leaf_40_clk_regs));
 sg13g2_dfrbpq_1 _10443_ (.RESET_B(net802),
    .D(net3636),
    .Q(\cpu.arbiter.i_wb_cpu_dbus_dat[4] ),
    .CLK(clknet_leaf_40_clk_regs));
 sg13g2_dfrbpq_1 _10444_ (.RESET_B(net801),
    .D(net3687),
    .Q(\cpu.arbiter.i_wb_cpu_dbus_dat[5] ),
    .CLK(clknet_leaf_40_clk_regs));
 sg13g2_dfrbpq_1 _10445_ (.RESET_B(net800),
    .D(net3633),
    .Q(\cpu.arbiter.i_wb_cpu_dbus_dat[6] ),
    .CLK(clknet_leaf_40_clk_regs));
 sg13g2_dfrbpq_1 _10446_ (.RESET_B(net799),
    .D(net3649),
    .Q(\cpu.arbiter.i_wb_cpu_dbus_dat[7] ),
    .CLK(clknet_leaf_40_clk_regs));
 sg13g2_dfrbpq_2 _10447_ (.RESET_B(net798),
    .D(_00491_),
    .Q(\cpu.arbiter.i_wb_cpu_dbus_dat[8] ),
    .CLK(clknet_leaf_31_clk_regs));
 sg13g2_dfrbpq_1 _10448_ (.RESET_B(net797),
    .D(net3553),
    .Q(\cpu.arbiter.i_wb_cpu_dbus_dat[9] ),
    .CLK(clknet_leaf_30_clk_regs));
 sg13g2_dfrbpq_1 _10449_ (.RESET_B(net796),
    .D(net3547),
    .Q(\cpu.arbiter.i_wb_cpu_dbus_dat[10] ),
    .CLK(clknet_leaf_11_clk_regs));
 sg13g2_dfrbpq_1 _10450_ (.RESET_B(net795),
    .D(net3611),
    .Q(\cpu.arbiter.i_wb_cpu_dbus_dat[11] ),
    .CLK(clknet_leaf_10_clk_regs));
 sg13g2_dfrbpq_1 _10451_ (.RESET_B(net794),
    .D(net3549),
    .Q(\cpu.arbiter.i_wb_cpu_dbus_dat[12] ),
    .CLK(clknet_leaf_10_clk_regs));
 sg13g2_dfrbpq_1 _10452_ (.RESET_B(net793),
    .D(net3618),
    .Q(\cpu.arbiter.i_wb_cpu_dbus_dat[13] ),
    .CLK(clknet_leaf_8_clk_regs));
 sg13g2_dfrbpq_1 _10453_ (.RESET_B(net792),
    .D(_00497_),
    .Q(\cpu.arbiter.i_wb_cpu_dbus_dat[14] ),
    .CLK(clknet_leaf_8_clk_regs));
 sg13g2_dfrbpq_1 _10454_ (.RESET_B(net791),
    .D(net3599),
    .Q(\cpu.arbiter.i_wb_cpu_dbus_dat[15] ),
    .CLK(clknet_leaf_9_clk_regs));
 sg13g2_dfrbpq_2 _10455_ (.RESET_B(net790),
    .D(_00499_),
    .Q(\cpu.arbiter.i_wb_cpu_dbus_dat[16] ),
    .CLK(clknet_leaf_9_clk_regs));
 sg13g2_dfrbpq_1 _10456_ (.RESET_B(net789),
    .D(net3589),
    .Q(\cpu.arbiter.i_wb_cpu_dbus_dat[17] ),
    .CLK(clknet_leaf_9_clk_regs));
 sg13g2_dfrbpq_1 _10457_ (.RESET_B(net788),
    .D(_00501_),
    .Q(\cpu.arbiter.i_wb_cpu_dbus_dat[18] ),
    .CLK(clknet_leaf_7_clk_regs));
 sg13g2_dfrbpq_1 _10458_ (.RESET_B(net787),
    .D(net3581),
    .Q(\cpu.arbiter.i_wb_cpu_dbus_dat[19] ),
    .CLK(clknet_leaf_3_clk_regs));
 sg13g2_dfrbpq_1 _10459_ (.RESET_B(net786),
    .D(net3522),
    .Q(\cpu.arbiter.i_wb_cpu_dbus_dat[20] ),
    .CLK(clknet_leaf_3_clk_regs));
 sg13g2_dfrbpq_1 _10460_ (.RESET_B(net785),
    .D(net3520),
    .Q(\cpu.arbiter.i_wb_cpu_dbus_dat[21] ),
    .CLK(clknet_leaf_7_clk_regs));
 sg13g2_dfrbpq_1 _10461_ (.RESET_B(net784),
    .D(net3551),
    .Q(\cpu.arbiter.i_wb_cpu_dbus_dat[22] ),
    .CLK(clknet_leaf_7_clk_regs));
 sg13g2_dfrbpq_1 _10462_ (.RESET_B(net783),
    .D(net3651),
    .Q(\cpu.arbiter.i_wb_cpu_dbus_dat[23] ),
    .CLK(clknet_leaf_9_clk_regs));
 sg13g2_dfrbpq_2 _10463_ (.RESET_B(net782),
    .D(_00507_),
    .Q(\cpu.cpu.decode.opcode[0] ),
    .CLK(clknet_leaf_42_clk_regs));
 sg13g2_dfrbpq_2 _10464_ (.RESET_B(net781),
    .D(_00508_),
    .Q(\cpu.cpu.decode.opcode[1] ),
    .CLK(clknet_leaf_41_clk_regs));
 sg13g2_dfrbpq_2 _10465_ (.RESET_B(net780),
    .D(_00509_),
    .Q(\cpu.cpu.decode.opcode[2] ),
    .CLK(clknet_leaf_34_clk_regs));
 sg13g2_dfrbpq_1 _10466_ (.RESET_B(net779),
    .D(_00510_),
    .Q(\cpu.arbiter.i_wb_cpu_dbus_we ),
    .CLK(clknet_leaf_44_clk_regs));
 sg13g2_dfrbpq_1 _10467_ (.RESET_B(net778),
    .D(_00511_),
    .Q(\cpu.cpu.branch_op ),
    .CLK(clknet_leaf_44_clk_regs));
 sg13g2_dfrbpq_2 _10468_ (.RESET_B(net777),
    .D(_00512_),
    .Q(\cpu.cpu.bne_or_bge ),
    .CLK(clknet_leaf_34_clk_regs));
 sg13g2_dfrbpq_1 _10469_ (.RESET_B(net776),
    .D(_00513_),
    .Q(\cpu.cpu.decode.co_mem_word ),
    .CLK(clknet_leaf_36_clk_regs));
 sg13g2_dfrbpq_2 _10470_ (.RESET_B(net775),
    .D(_00514_),
    .Q(\cpu.cpu.bufreg.i_right_shift_op ),
    .CLK(clknet_leaf_30_clk_regs));
 sg13g2_dfrbpq_1 _10471_ (.RESET_B(net774),
    .D(net3517),
    .Q(\cpu.cpu.decode.co_ebreak ),
    .CLK(clknet_leaf_29_clk_regs));
 sg13g2_dfrbpq_2 _10472_ (.RESET_B(net773),
    .D(_00516_),
    .Q(\cpu.cpu.immdec.gen_immdec_w_eq_1.imm24_20[0] ),
    .CLK(clknet_leaf_12_clk_regs));
 sg13g2_dfrbpq_1 _10473_ (.RESET_B(net772),
    .D(net3708),
    .Q(\cpu.cpu.immdec.gen_immdec_w_eq_1.imm24_20[1] ),
    .CLK(clknet_leaf_15_clk_regs));
 sg13g2_dfrbpq_1 _10474_ (.RESET_B(net771),
    .D(_00518_),
    .Q(\cpu.cpu.immdec.gen_immdec_w_eq_1.imm24_20[2] ),
    .CLK(clknet_leaf_14_clk_regs));
 sg13g2_dfrbpq_1 _10475_ (.RESET_B(net770),
    .D(_00519_),
    .Q(\cpu.cpu.immdec.gen_immdec_w_eq_1.imm24_20[3] ),
    .CLK(clknet_leaf_12_clk_regs));
 sg13g2_dfrbpq_1 _10476_ (.RESET_B(net769),
    .D(_00520_),
    .Q(\cpu.cpu.immdec.gen_immdec_w_eq_1.imm24_20[4] ),
    .CLK(clknet_leaf_12_clk_regs));
 sg13g2_dfrbpq_2 _10477_ (.RESET_B(net768),
    .D(_00521_),
    .Q(\cpu.cpu.immdec.gen_immdec_w_eq_1.imm30_25[0] ),
    .CLK(clknet_leaf_4_clk_regs));
 sg13g2_dfrbpq_1 _10478_ (.RESET_B(net767),
    .D(net3399),
    .Q(\cpu.cpu.immdec.gen_immdec_w_eq_1.imm30_25[1] ),
    .CLK(clknet_leaf_1_clk_regs));
 sg13g2_dfrbpq_1 _10479_ (.RESET_B(net766),
    .D(net3363),
    .Q(\cpu.cpu.immdec.gen_immdec_w_eq_1.imm30_25[2] ),
    .CLK(clknet_leaf_171_clk_regs));
 sg13g2_dfrbpq_1 _10480_ (.RESET_B(net765),
    .D(net3374),
    .Q(\cpu.cpu.immdec.gen_immdec_w_eq_1.imm30_25[3] ),
    .CLK(clknet_leaf_0_clk_regs));
 sg13g2_dfrbpq_1 _10481_ (.RESET_B(net764),
    .D(net3458),
    .Q(\cpu.cpu.immdec.gen_immdec_w_eq_1.imm30_25[4] ),
    .CLK(clknet_leaf_1_clk_regs));
 sg13g2_dfrbpq_1 _10482_ (.RESET_B(net763),
    .D(net3421),
    .Q(\cpu.cpu.immdec.gen_immdec_w_eq_1.imm30_25[5] ),
    .CLK(clknet_leaf_11_clk_regs));
 sg13g2_dfrbpq_1 _10483_ (.RESET_B(net762),
    .D(net3255),
    .Q(\cpu.cpu.immdec.gen_immdec_w_eq_1.imm7 ),
    .CLK(clknet_leaf_27_clk_regs));
 sg13g2_dfrbpq_1 _10484_ (.RESET_B(net761),
    .D(net3511),
    .Q(\cpu.cpu.immdec.gen_immdec_w_eq_1.imm19_12_20[0] ),
    .CLK(clknet_leaf_29_clk_regs));
 sg13g2_dfrbpq_1 _10485_ (.RESET_B(net760),
    .D(net3441),
    .Q(\cpu.cpu.immdec.gen_immdec_w_eq_1.imm19_12_20[1] ),
    .CLK(clknet_leaf_12_clk_regs));
 sg13g2_dfrbpq_1 _10486_ (.RESET_B(net759),
    .D(net3488),
    .Q(\cpu.cpu.immdec.gen_immdec_w_eq_1.imm19_12_20[2] ),
    .CLK(clknet_leaf_12_clk_regs));
 sg13g2_dfrbpq_1 _10487_ (.RESET_B(net758),
    .D(net3436),
    .Q(\cpu.cpu.immdec.gen_immdec_w_eq_1.imm19_12_20[3] ),
    .CLK(clknet_leaf_11_clk_regs));
 sg13g2_dfrbpq_1 _10488_ (.RESET_B(net757),
    .D(net3419),
    .Q(\cpu.cpu.csr_imm [0]),
    .CLK(clknet_leaf_12_clk_regs));
 sg13g2_dfrbpq_1 _10489_ (.RESET_B(net756),
    .D(_00533_),
    .Q(\cpu.cpu.immdec.gen_immdec_w_eq_1.imm19_12_20[5] ),
    .CLK(clknet_leaf_12_clk_regs));
 sg13g2_dfrbpq_1 _10490_ (.RESET_B(net755),
    .D(_00534_),
    .Q(\cpu.cpu.immdec.gen_immdec_w_eq_1.imm19_12_20[6] ),
    .CLK(clknet_leaf_12_clk_regs));
 sg13g2_dfrbpq_2 _10491_ (.RESET_B(net754),
    .D(net3579),
    .Q(\cpu.cpu.immdec.gen_immdec_w_eq_1.imm19_12_20[7] ),
    .CLK(clknet_leaf_6_clk_regs));
 sg13g2_dfrbpq_1 _10492_ (.RESET_B(net753),
    .D(net3625),
    .Q(\cpu.cpu.immdec.gen_immdec_w_eq_1.imm19_12_20[8] ),
    .CLK(clknet_leaf_6_clk_regs));
 sg13g2_dfrbpq_1 _10493_ (.RESET_B(net752),
    .D(net3641),
    .Q(\cpu.cpu.immdec.gen_immdec_w_eq_1.imm31 ),
    .CLK(clknet_leaf_29_clk_regs));
 sg13g2_dfrbpq_2 _10494_ (.RESET_B(net751),
    .D(net3733),
    .Q(\cpu.cpu.bufreg.i_sh_signed ),
    .CLK(clknet_leaf_30_clk_regs));
 sg13g2_dfrbpq_1 _10495_ (.RESET_B(net1333),
    .D(_00539_),
    .Q(\cpu.cpu.alu.cmp_r ),
    .CLK(clknet_leaf_34_clk_regs));
 sg13g2_dfrbpq_1 _10496_ (.RESET_B(net750),
    .D(_00062_),
    .Q(\cpu.cpu.bufreg.c_r [0]),
    .CLK(clknet_leaf_29_clk_regs));
 sg13g2_dfrbpq_2 _10497_ (.RESET_B(net749),
    .D(_00540_),
    .Q(\cpu.arbiter.i_wb_cpu_dbus_dat[24] ),
    .CLK(clknet_leaf_0_clk_regs));
 sg13g2_dfrbpq_2 _10498_ (.RESET_B(net748),
    .D(net3735),
    .Q(\cpu.arbiter.i_wb_cpu_dbus_dat[25] ),
    .CLK(clknet_leaf_1_clk_regs));
 sg13g2_dfrbpq_2 _10499_ (.RESET_B(net747),
    .D(_00542_),
    .Q(\cpu.arbiter.i_wb_cpu_dbus_dat[26] ),
    .CLK(clknet_leaf_2_clk_regs));
 sg13g2_dfrbpq_2 _10500_ (.RESET_B(net746),
    .D(net3675),
    .Q(\cpu.arbiter.i_wb_cpu_dbus_dat[27] ),
    .CLK(clknet_leaf_2_clk_regs));
 sg13g2_dfrbpq_2 _10501_ (.RESET_B(net745),
    .D(net3740),
    .Q(\cpu.arbiter.i_wb_cpu_dbus_dat[28] ),
    .CLK(clknet_leaf_2_clk_regs));
 sg13g2_dfrbpq_1 _10502_ (.RESET_B(net744),
    .D(net3743),
    .Q(\cpu.arbiter.i_wb_cpu_dbus_dat[29] ),
    .CLK(clknet_leaf_7_clk_regs));
 sg13g2_dfrbpq_1 _10503_ (.RESET_B(net743),
    .D(net3451),
    .Q(\cpu.arbiter.i_wb_cpu_dbus_dat[30] ),
    .CLK(clknet_leaf_30_clk_regs));
 sg13g2_dfrbpq_1 _10504_ (.RESET_B(net742),
    .D(net3465),
    .Q(\cpu.arbiter.i_wb_cpu_dbus_dat[31] ),
    .CLK(clknet_leaf_30_clk_regs));
 sg13g2_dfrbpq_2 _10505_ (.RESET_B(net741),
    .D(net3748),
    .Q(\cpu.cpu.bufreg.data[0] ),
    .CLK(clknet_leaf_33_clk_regs));
 sg13g2_dfrbpq_2 _10506_ (.RESET_B(net740),
    .D(_00549_),
    .Q(\cpu.cpu.bufreg.data[1] ),
    .CLK(clknet_leaf_33_clk_regs));
 sg13g2_dfrbpq_1 _10507_ (.RESET_B(net739),
    .D(net3145),
    .Q(\rf_ram.RAM[10][0] ),
    .CLK(clknet_leaf_16_clk_regs));
 sg13g2_dfrbpq_1 _10508_ (.RESET_B(net738),
    .D(_00551_),
    .Q(\rf_ram.RAM[10][1] ),
    .CLK(clknet_leaf_54_clk_regs));
 sg13g2_dfrbpq_1 _10509_ (.RESET_B(net737),
    .D(_00552_),
    .Q(\rf_ram.RAM[10][2] ),
    .CLK(clknet_leaf_78_clk_regs));
 sg13g2_dfrbpq_1 _10510_ (.RESET_B(net736),
    .D(_00553_),
    .Q(\rf_ram.RAM[10][3] ),
    .CLK(clknet_leaf_79_clk_regs));
 sg13g2_dfrbpq_1 _10511_ (.RESET_B(net735),
    .D(_00554_),
    .Q(\rf_ram.RAM[10][4] ),
    .CLK(clknet_leaf_80_clk_regs));
 sg13g2_dfrbpq_1 _10512_ (.RESET_B(net734),
    .D(_00555_),
    .Q(\rf_ram.RAM[10][5] ),
    .CLK(clknet_leaf_80_clk_regs));
 sg13g2_dfrbpq_1 _10513_ (.RESET_B(net733),
    .D(_00556_),
    .Q(\rf_ram.RAM[10][6] ),
    .CLK(clknet_leaf_100_clk_regs));
 sg13g2_dfrbpq_1 _10514_ (.RESET_B(net732),
    .D(_00557_),
    .Q(\rf_ram.RAM[10][7] ),
    .CLK(clknet_leaf_98_clk_regs));
 sg13g2_dfrbpq_1 _10515_ (.RESET_B(net731),
    .D(_00558_),
    .Q(\rf_ram.RAM[10][8] ),
    .CLK(clknet_leaf_113_clk_regs));
 sg13g2_dfrbpq_1 _10516_ (.RESET_B(net730),
    .D(_00559_),
    .Q(\rf_ram.RAM[10][9] ),
    .CLK(clknet_leaf_122_clk_regs));
 sg13g2_dfrbpq_1 _10517_ (.RESET_B(net729),
    .D(_00560_),
    .Q(\rf_ram.RAM[10][10] ),
    .CLK(clknet_leaf_112_clk_regs));
 sg13g2_dfrbpq_1 _10518_ (.RESET_B(net728),
    .D(_00561_),
    .Q(\rf_ram.RAM[10][11] ),
    .CLK(clknet_leaf_130_clk_regs));
 sg13g2_dfrbpq_1 _10519_ (.RESET_B(net727),
    .D(_00562_),
    .Q(\rf_ram.RAM[10][12] ),
    .CLK(clknet_leaf_130_clk_regs));
 sg13g2_dfrbpq_1 _10520_ (.RESET_B(net726),
    .D(_00563_),
    .Q(\rf_ram.RAM[10][13] ),
    .CLK(clknet_leaf_98_clk_regs));
 sg13g2_dfrbpq_1 _10521_ (.RESET_B(net725),
    .D(_00564_),
    .Q(\rf_ram.RAM[10][14] ),
    .CLK(clknet_leaf_158_clk_regs));
 sg13g2_dfrbpq_1 _10522_ (.RESET_B(net724),
    .D(_00565_),
    .Q(\rf_ram.RAM[10][15] ),
    .CLK(clknet_leaf_109_clk_regs));
 sg13g2_dfrbpq_1 _10523_ (.RESET_B(net723),
    .D(_00566_),
    .Q(\rf_ram.RAM[10][16] ),
    .CLK(clknet_leaf_68_clk_regs));
 sg13g2_dfrbpq_1 _10524_ (.RESET_B(net722),
    .D(_00567_),
    .Q(\rf_ram.RAM[10][17] ),
    .CLK(clknet_leaf_137_clk_regs));
 sg13g2_dfrbpq_1 _10525_ (.RESET_B(net721),
    .D(_00568_),
    .Q(\rf_ram.RAM[10][18] ),
    .CLK(clknet_leaf_136_clk_regs));
 sg13g2_dfrbpq_1 _10526_ (.RESET_B(net720),
    .D(_00569_),
    .Q(\rf_ram.RAM[10][19] ),
    .CLK(clknet_leaf_161_clk_regs));
 sg13g2_dfrbpq_1 _10527_ (.RESET_B(net719),
    .D(_00570_),
    .Q(\rf_ram.RAM[10][20] ),
    .CLK(clknet_leaf_152_clk_regs));
 sg13g2_dfrbpq_1 _10528_ (.RESET_B(net718),
    .D(_00571_),
    .Q(\rf_ram.RAM[10][21] ),
    .CLK(clknet_leaf_61_clk_regs));
 sg13g2_dfrbpq_1 _10529_ (.RESET_B(net717),
    .D(_00572_),
    .Q(\rf_ram.RAM[10][22] ),
    .CLK(clknet_leaf_105_clk_regs));
 sg13g2_dfrbpq_1 _10530_ (.RESET_B(net716),
    .D(_00573_),
    .Q(\rf_ram.RAM[10][23] ),
    .CLK(clknet_leaf_21_clk_regs));
 sg13g2_dfrbpq_1 _10531_ (.RESET_B(net715),
    .D(_00574_),
    .Q(\rf_ram.RAM[10][24] ),
    .CLK(clknet_leaf_72_clk_regs));
 sg13g2_dfrbpq_1 _10532_ (.RESET_B(net714),
    .D(_00575_),
    .Q(\rf_ram.RAM[10][25] ),
    .CLK(clknet_leaf_57_clk_regs));
 sg13g2_dfrbpq_1 _10533_ (.RESET_B(net713),
    .D(_00576_),
    .Q(\rf_ram.RAM[10][26] ),
    .CLK(clknet_leaf_58_clk_regs));
 sg13g2_dfrbpq_1 _10534_ (.RESET_B(net712),
    .D(_00577_),
    .Q(\rf_ram.RAM[10][27] ),
    .CLK(clknet_leaf_35_clk_regs));
 sg13g2_dfrbpq_1 _10535_ (.RESET_B(net711),
    .D(_00578_),
    .Q(\rf_ram.RAM[10][28] ),
    .CLK(clknet_leaf_28_clk_regs));
 sg13g2_dfrbpq_1 _10536_ (.RESET_B(net710),
    .D(_00579_),
    .Q(\rf_ram.RAM[10][29] ),
    .CLK(clknet_leaf_5_clk_regs));
 sg13g2_dfrbpq_1 _10537_ (.RESET_B(net709),
    .D(_00580_),
    .Q(\rf_ram.RAM[10][30] ),
    .CLK(clknet_leaf_164_clk_regs));
 sg13g2_dfrbpq_1 _10538_ (.RESET_B(net1334),
    .D(_00581_),
    .Q(\rf_ram.RAM[10][31] ),
    .CLK(clknet_leaf_167_clk_regs));
 sg13g2_dfrbpq_1 _10539_ (.RESET_B(net1367),
    .D(_00064_),
    .Q(\cpu.cpu.ctrl.pc_plus_offset_cy_r_w [0]),
    .CLK(clknet_leaf_34_clk_regs));
 sg13g2_dfrbpq_1 _10540_ (.RESET_B(net708),
    .D(net3434),
    .Q(\cpu.cpu.ctrl.pc_plus_4_cy_r_w [0]),
    .CLK(clknet_leaf_32_clk_regs));
 sg13g2_dfrbpq_2 _10541_ (.RESET_B(net707),
    .D(_00582_),
    .Q(\cpu.cpu.ctrl.pc [0]),
    .CLK(clknet_leaf_32_clk_regs));
 sg13g2_dfrbpq_1 _10542_ (.RESET_B(net705),
    .D(_00583_),
    .Q(\cpu.arbiter.i_wb_cpu_ibus_adr[1] ),
    .CLK(clknet_leaf_33_clk_regs));
 sg13g2_dfrbpq_1 _10543_ (.RESET_B(net703),
    .D(_00584_),
    .Q(\cpu.arbiter.i_wb_cpu_ibus_adr[2] ),
    .CLK(clknet_leaf_37_clk_regs));
 sg13g2_dfrbpq_1 _10544_ (.RESET_B(net701),
    .D(_00585_),
    .Q(\cpu.arbiter.i_wb_cpu_ibus_adr[3] ),
    .CLK(clknet_leaf_38_clk_regs));
 sg13g2_dfrbpq_1 _10545_ (.RESET_B(net699),
    .D(_00586_),
    .Q(\cpu.arbiter.i_wb_cpu_ibus_adr[4] ),
    .CLK(clknet_leaf_37_clk_regs));
 sg13g2_dfrbpq_1 _10546_ (.RESET_B(net697),
    .D(_00587_),
    .Q(\cpu.arbiter.i_wb_cpu_ibus_adr[5] ),
    .CLK(clknet_leaf_38_clk_regs));
 sg13g2_dfrbpq_1 _10547_ (.RESET_B(net695),
    .D(_00588_),
    .Q(\cpu.arbiter.i_wb_cpu_ibus_adr[6] ),
    .CLK(clknet_leaf_33_clk_regs));
 sg13g2_dfrbpq_1 _10548_ (.RESET_B(net693),
    .D(_00589_),
    .Q(\cpu.arbiter.i_wb_cpu_ibus_adr[7] ),
    .CLK(clknet_leaf_33_clk_regs));
 sg13g2_dfrbpq_1 _10549_ (.RESET_B(net691),
    .D(_00590_),
    .Q(\cpu.arbiter.i_wb_cpu_ibus_adr[8] ),
    .CLK(clknet_leaf_32_clk_regs));
 sg13g2_dfrbpq_1 _10550_ (.RESET_B(net689),
    .D(_00591_),
    .Q(\cpu.arbiter.i_wb_cpu_ibus_adr[9] ),
    .CLK(clknet_leaf_32_clk_regs));
 sg13g2_dfrbpq_2 _10551_ (.RESET_B(net687),
    .D(_00592_),
    .Q(\cpu.arbiter.i_wb_cpu_ibus_adr[10] ),
    .CLK(clknet_leaf_10_clk_regs));
 sg13g2_dfrbpq_1 _10552_ (.RESET_B(net685),
    .D(_00593_),
    .Q(\cpu.arbiter.i_wb_cpu_ibus_adr[11] ),
    .CLK(clknet_leaf_10_clk_regs));
 sg13g2_dfrbpq_1 _10553_ (.RESET_B(net683),
    .D(_00594_),
    .Q(\cpu.arbiter.i_wb_cpu_ibus_adr[12] ),
    .CLK(clknet_leaf_10_clk_regs));
 sg13g2_dfrbpq_1 _10554_ (.RESET_B(net681),
    .D(_00595_),
    .Q(\cpu.arbiter.i_wb_cpu_ibus_adr[13] ),
    .CLK(clknet_leaf_8_clk_regs));
 sg13g2_dfrbpq_1 _10555_ (.RESET_B(net679),
    .D(_00596_),
    .Q(\cpu.arbiter.i_wb_cpu_ibus_adr[14] ),
    .CLK(clknet_leaf_8_clk_regs));
 sg13g2_dfrbpq_2 _10556_ (.RESET_B(net677),
    .D(_00597_),
    .Q(\cpu.arbiter.i_wb_cpu_ibus_adr[15] ),
    .CLK(clknet_leaf_2_clk_regs));
 sg13g2_dfrbpq_1 _10557_ (.RESET_B(net516),
    .D(_00598_),
    .Q(\cpu.arbiter.i_wb_cpu_ibus_adr[16] ),
    .CLK(clknet_leaf_2_clk_regs));
 sg13g2_dfrbpq_1 _10558_ (.RESET_B(net512),
    .D(_00599_),
    .Q(\cpu.arbiter.i_wb_cpu_ibus_adr[17] ),
    .CLK(clknet_leaf_1_clk_regs));
 sg13g2_dfrbpq_1 _10559_ (.RESET_B(net822),
    .D(_00600_),
    .Q(\cpu.arbiter.i_wb_cpu_ibus_adr[18] ),
    .CLK(clknet_leaf_1_clk_regs));
 sg13g2_dfrbpq_1 _10560_ (.RESET_B(net811),
    .D(_00601_),
    .Q(\cpu.arbiter.i_wb_cpu_ibus_adr[19] ),
    .CLK(clknet_leaf_1_clk_regs));
 sg13g2_dfrbpq_1 _10561_ (.RESET_B(net704),
    .D(_00602_),
    .Q(\cpu.arbiter.i_wb_cpu_ibus_adr[20] ),
    .CLK(clknet_leaf_0_clk_regs));
 sg13g2_dfrbpq_1 _10562_ (.RESET_B(net700),
    .D(_00603_),
    .Q(\cpu.arbiter.i_wb_cpu_ibus_adr[21] ),
    .CLK(clknet_leaf_172_clk_regs));
 sg13g2_dfrbpq_1 _10563_ (.RESET_B(net696),
    .D(_00604_),
    .Q(\cpu.arbiter.i_wb_cpu_ibus_adr[22] ),
    .CLK(clknet_leaf_0_clk_regs));
 sg13g2_dfrbpq_1 _10564_ (.RESET_B(net692),
    .D(_00605_),
    .Q(\cpu.arbiter.i_wb_cpu_ibus_adr[23] ),
    .CLK(clknet_leaf_0_clk_regs));
 sg13g2_dfrbpq_1 _10565_ (.RESET_B(net688),
    .D(_00606_),
    .Q(\cpu.arbiter.i_wb_cpu_ibus_adr[24] ),
    .CLK(clknet_leaf_0_clk_regs));
 sg13g2_dfrbpq_1 _10566_ (.RESET_B(net684),
    .D(_00607_),
    .Q(\cpu.arbiter.i_wb_cpu_ibus_adr[25] ),
    .CLK(clknet_leaf_0_clk_regs));
 sg13g2_dfrbpq_1 _10567_ (.RESET_B(net680),
    .D(_00608_),
    .Q(\cpu.arbiter.i_wb_cpu_ibus_adr[26] ),
    .CLK(clknet_leaf_1_clk_regs));
 sg13g2_dfrbpq_1 _10568_ (.RESET_B(net676),
    .D(_00609_),
    .Q(\cpu.arbiter.i_wb_cpu_ibus_adr[27] ),
    .CLK(clknet_leaf_172_clk_regs));
 sg13g2_dfrbpq_1 _10569_ (.RESET_B(net510),
    .D(_00610_),
    .Q(\cpu.arbiter.i_wb_cpu_ibus_adr[28] ),
    .CLK(clknet_leaf_172_clk_regs));
 sg13g2_dfrbpq_1 _10570_ (.RESET_B(net706),
    .D(_00611_),
    .Q(\cpu.arbiter.i_wb_cpu_ibus_adr[29] ),
    .CLK(clknet_leaf_172_clk_regs));
 sg13g2_dfrbpq_1 _10571_ (.RESET_B(net698),
    .D(_00612_),
    .Q(\cpu.arbiter.i_wb_cpu_ibus_adr[30] ),
    .CLK(clknet_leaf_172_clk_regs));
 sg13g2_dfrbpq_1 _10572_ (.RESET_B(net686),
    .D(_00613_),
    .Q(\cpu.arbiter.i_wb_cpu_ibus_adr[31] ),
    .CLK(clknet_leaf_172_clk_regs));
 sg13g2_dfrbpq_1 _10573_ (.RESET_B(net690),
    .D(net3766),
    .Q(\cpu.cpu.alu.add_cy_r [0]),
    .CLK(clknet_leaf_34_clk_regs));
 sg13g2_dfrbpq_2 _10574_ (.RESET_B(net682),
    .D(net3478),
    .Q(\cpu.cpu.immdec.gen_immdec_w_eq_1.imm11_7[0] ),
    .CLK(clknet_leaf_27_clk_regs));
 sg13g2_dfrbpq_2 _10575_ (.RESET_B(net678),
    .D(net3583),
    .Q(\cpu.cpu.immdec.gen_immdec_w_eq_1.imm11_7[1] ),
    .CLK(clknet_leaf_29_clk_regs));
 sg13g2_dfrbpq_2 _10576_ (.RESET_B(net514),
    .D(net3711),
    .Q(\cpu.cpu.immdec.gen_immdec_w_eq_1.imm11_7[2] ),
    .CLK(clknet_leaf_29_clk_regs));
 sg13g2_dfrbpq_2 _10577_ (.RESET_B(net813),
    .D(_00617_),
    .Q(\cpu.cpu.immdec.gen_immdec_w_eq_1.imm11_7[3] ),
    .CLK(clknet_leaf_13_clk_regs));
 sg13g2_dfrbpq_2 _10578_ (.RESET_B(net702),
    .D(_00618_),
    .Q(\cpu.cpu.immdec.gen_immdec_w_eq_1.imm11_7[4] ),
    .CLK(clknet_leaf_13_clk_regs));
 sg13g2_dfrbpq_1 _10579_ (.RESET_B(net694),
    .D(_00619_),
    .Q(\ram_spi_if.spi_mosi ),
    .CLK(net1380));
 sg13g2_tiehi _09876__19 (.L_HI(net19));
 sg13g2_tiehi _09875__20 (.L_HI(net20));
 sg13g2_tiehi _09874__21 (.L_HI(net21));
 sg13g2_tiehi _09873__22 (.L_HI(net22));
 sg13g2_tiehi _09872__23 (.L_HI(net23));
 sg13g2_tiehi _09871__24 (.L_HI(net24));
 sg13g2_tiehi _09870__25 (.L_HI(net25));
 sg13g2_tiehi _09869__26 (.L_HI(net26));
 sg13g2_tiehi _09868__27 (.L_HI(net27));
 sg13g2_tiehi _09867__28 (.L_HI(net28));
 sg13g2_tiehi _09866__29 (.L_HI(net29));
 sg13g2_tiehi _09865__30 (.L_HI(net30));
 sg13g2_tiehi _09864__31 (.L_HI(net31));
 sg13g2_tiehi _09863__32 (.L_HI(net32));
 sg13g2_tiehi _09862__33 (.L_HI(net33));
 sg13g2_tiehi _09861__34 (.L_HI(net34));
 sg13g2_tiehi _09860__35 (.L_HI(net35));
 sg13g2_tiehi _09859__36 (.L_HI(net36));
 sg13g2_tiehi _09858__37 (.L_HI(net37));
 sg13g2_tiehi _09857__38 (.L_HI(net38));
 sg13g2_tiehi _09856__39 (.L_HI(net39));
 sg13g2_tiehi _09855__40 (.L_HI(net40));
 sg13g2_tiehi _09854__41 (.L_HI(net41));
 sg13g2_tiehi _09853__42 (.L_HI(net42));
 sg13g2_tiehi _09852__43 (.L_HI(net43));
 sg13g2_tiehi _09851__44 (.L_HI(net44));
 sg13g2_tiehi _09850__45 (.L_HI(net45));
 sg13g2_tiehi _09849__46 (.L_HI(net46));
 sg13g2_tiehi _09848__47 (.L_HI(net47));
 sg13g2_tiehi _09847__48 (.L_HI(net48));
 sg13g2_tiehi _09846__49 (.L_HI(net49));
 sg13g2_tiehi _09845__50 (.L_HI(net50));
 sg13g2_tiehi _09844__51 (.L_HI(net51));
 sg13g2_tiehi _09843__52 (.L_HI(net52));
 sg13g2_tiehi _09842__53 (.L_HI(net53));
 sg13g2_tiehi _09841__54 (.L_HI(net54));
 sg13g2_tiehi _09840__55 (.L_HI(net55));
 sg13g2_tiehi _09839__56 (.L_HI(net56));
 sg13g2_tiehi _09838__57 (.L_HI(net57));
 sg13g2_tiehi _09837__58 (.L_HI(net58));
 sg13g2_tiehi _09836__59 (.L_HI(net59));
 sg13g2_tiehi _09835__60 (.L_HI(net60));
 sg13g2_tiehi _09834__61 (.L_HI(net61));
 sg13g2_tiehi _09833__62 (.L_HI(net62));
 sg13g2_tiehi _09832__63 (.L_HI(net63));
 sg13g2_tiehi _09831__64 (.L_HI(net64));
 sg13g2_tiehi _09830__65 (.L_HI(net65));
 sg13g2_tiehi _09829__66 (.L_HI(net66));
 sg13g2_tiehi _09828__67 (.L_HI(net67));
 sg13g2_tiehi _09827__68 (.L_HI(net68));
 sg13g2_tiehi _09826__69 (.L_HI(net69));
 sg13g2_tiehi _09825__70 (.L_HI(net70));
 sg13g2_tiehi _09824__71 (.L_HI(net71));
 sg13g2_tiehi _09823__72 (.L_HI(net72));
 sg13g2_tiehi _09822__73 (.L_HI(net73));
 sg13g2_tiehi _09821__74 (.L_HI(net74));
 sg13g2_tiehi _09820__75 (.L_HI(net75));
 sg13g2_tiehi _09819__76 (.L_HI(net76));
 sg13g2_tiehi _09818__77 (.L_HI(net77));
 sg13g2_tiehi _09817__78 (.L_HI(net78));
 sg13g2_tiehi _09816__79 (.L_HI(net79));
 sg13g2_tiehi _09815__80 (.L_HI(net80));
 sg13g2_tiehi _09814__81 (.L_HI(net81));
 sg13g2_tiehi _09214__82 (.L_HI(net82));
 sg13g2_tiehi _09277__83 (.L_HI(net83));
 sg13g2_tiehi _09813__84 (.L_HI(net84));
 sg13g2_tiehi _09812__85 (.L_HI(net85));
 sg13g2_tiehi _09811__86 (.L_HI(net86));
 sg13g2_tiehi _09810__87 (.L_HI(net87));
 sg13g2_tiehi _09809__88 (.L_HI(net88));
 sg13g2_tiehi _09808__89 (.L_HI(net89));
 sg13g2_tiehi _09807__90 (.L_HI(net90));
 sg13g2_tiehi _09806__91 (.L_HI(net91));
 sg13g2_tiehi _09805__92 (.L_HI(net92));
 sg13g2_tiehi _09804__93 (.L_HI(net93));
 sg13g2_tiehi _09803__94 (.L_HI(net94));
 sg13g2_tiehi _09802__95 (.L_HI(net95));
 sg13g2_tiehi _09801__96 (.L_HI(net96));
 sg13g2_tiehi _09800__97 (.L_HI(net97));
 sg13g2_tiehi _09799__98 (.L_HI(net98));
 sg13g2_tiehi _09798__99 (.L_HI(net99));
 sg13g2_tiehi _09797__100 (.L_HI(net100));
 sg13g2_tiehi _09796__101 (.L_HI(net101));
 sg13g2_tiehi _09795__102 (.L_HI(net102));
 sg13g2_tiehi _09794__103 (.L_HI(net103));
 sg13g2_tiehi _09793__104 (.L_HI(net104));
 sg13g2_tiehi _09792__105 (.L_HI(net105));
 sg13g2_tiehi _09791__106 (.L_HI(net106));
 sg13g2_tiehi _09790__107 (.L_HI(net107));
 sg13g2_tiehi _09789__108 (.L_HI(net108));
 sg13g2_tiehi _09788__109 (.L_HI(net109));
 sg13g2_tiehi _09787__110 (.L_HI(net110));
 sg13g2_tiehi _09786__111 (.L_HI(net111));
 sg13g2_tiehi _09785__112 (.L_HI(net112));
 sg13g2_tiehi _09784__113 (.L_HI(net113));
 sg13g2_tiehi _09783__114 (.L_HI(net114));
 sg13g2_tiehi _09782__115 (.L_HI(net115));
 sg13g2_tiehi _09781__116 (.L_HI(net116));
 sg13g2_tiehi _09780__117 (.L_HI(net117));
 sg13g2_tiehi _09779__118 (.L_HI(net118));
 sg13g2_tiehi _09778__119 (.L_HI(net119));
 sg13g2_tiehi _09777__120 (.L_HI(net120));
 sg13g2_tiehi _09776__121 (.L_HI(net121));
 sg13g2_tiehi _09775__122 (.L_HI(net122));
 sg13g2_tiehi _09774__123 (.L_HI(net123));
 sg13g2_tiehi _09773__124 (.L_HI(net124));
 sg13g2_tiehi _09772__125 (.L_HI(net125));
 sg13g2_tiehi _09771__126 (.L_HI(net126));
 sg13g2_tiehi _09770__127 (.L_HI(net127));
 sg13g2_tiehi _09769__128 (.L_HI(net128));
 sg13g2_tiehi _09768__129 (.L_HI(net129));
 sg13g2_tiehi _09767__130 (.L_HI(net130));
 sg13g2_tiehi _09766__131 (.L_HI(net131));
 sg13g2_tiehi _09765__132 (.L_HI(net132));
 sg13g2_tiehi _09764__133 (.L_HI(net133));
 sg13g2_tiehi _09763__134 (.L_HI(net134));
 sg13g2_tiehi _09762__135 (.L_HI(net135));
 sg13g2_tiehi _09761__136 (.L_HI(net136));
 sg13g2_tiehi _09760__137 (.L_HI(net137));
 sg13g2_tiehi _09759__138 (.L_HI(net138));
 sg13g2_tiehi _09758__139 (.L_HI(net139));
 sg13g2_tiehi _09757__140 (.L_HI(net140));
 sg13g2_tiehi _09756__141 (.L_HI(net141));
 sg13g2_tiehi _09755__142 (.L_HI(net142));
 sg13g2_tiehi _09754__143 (.L_HI(net143));
 sg13g2_tiehi _09753__144 (.L_HI(net144));
 sg13g2_tiehi _09752__145 (.L_HI(net145));
 sg13g2_tiehi _09751__146 (.L_HI(net146));
 sg13g2_tiehi _09750__147 (.L_HI(net147));
 sg13g2_tiehi _09749__148 (.L_HI(net148));
 sg13g2_tiehi _09748__149 (.L_HI(net149));
 sg13g2_tiehi _09747__150 (.L_HI(net150));
 sg13g2_tiehi _09746__151 (.L_HI(net151));
 sg13g2_tiehi _09745__152 (.L_HI(net152));
 sg13g2_tiehi _09744__153 (.L_HI(net153));
 sg13g2_tiehi _09743__154 (.L_HI(net154));
 sg13g2_tiehi _09742__155 (.L_HI(net155));
 sg13g2_tiehi _09741__156 (.L_HI(net156));
 sg13g2_tiehi _09740__157 (.L_HI(net157));
 sg13g2_tiehi _09739__158 (.L_HI(net158));
 sg13g2_tiehi _09738__159 (.L_HI(net159));
 sg13g2_tiehi _09737__160 (.L_HI(net160));
 sg13g2_tiehi _09736__161 (.L_HI(net161));
 sg13g2_tiehi _09735__162 (.L_HI(net162));
 sg13g2_tiehi _09734__163 (.L_HI(net163));
 sg13g2_tiehi _09733__164 (.L_HI(net164));
 sg13g2_tiehi _09732__165 (.L_HI(net165));
 sg13g2_tiehi _09731__166 (.L_HI(net166));
 sg13g2_tiehi _09730__167 (.L_HI(net167));
 sg13g2_tiehi _09729__168 (.L_HI(net168));
 sg13g2_tiehi _09728__169 (.L_HI(net169));
 sg13g2_tiehi _09727__170 (.L_HI(net170));
 sg13g2_tiehi _09726__171 (.L_HI(net171));
 sg13g2_tiehi _09725__172 (.L_HI(net172));
 sg13g2_tiehi _09724__173 (.L_HI(net173));
 sg13g2_tiehi _09723__174 (.L_HI(net174));
 sg13g2_tiehi _09722__175 (.L_HI(net175));
 sg13g2_tiehi _09721__176 (.L_HI(net176));
 sg13g2_tiehi _09720__177 (.L_HI(net177));
 sg13g2_tiehi _09719__178 (.L_HI(net178));
 sg13g2_tiehi _09718__179 (.L_HI(net179));
 sg13g2_tiehi _09717__180 (.L_HI(net180));
 sg13g2_tiehi _09716__181 (.L_HI(net181));
 sg13g2_tiehi _09715__182 (.L_HI(net182));
 sg13g2_tiehi _09714__183 (.L_HI(net183));
 sg13g2_tiehi _09713__184 (.L_HI(net184));
 sg13g2_tiehi _09712__185 (.L_HI(net185));
 sg13g2_tiehi _09711__186 (.L_HI(net186));
 sg13g2_tiehi _09710__187 (.L_HI(net187));
 sg13g2_tiehi _09709__188 (.L_HI(net188));
 sg13g2_tiehi _09708__189 (.L_HI(net189));
 sg13g2_tiehi _09707__190 (.L_HI(net190));
 sg13g2_tiehi _09706__191 (.L_HI(net191));
 sg13g2_tiehi _09705__192 (.L_HI(net192));
 sg13g2_tiehi _09704__193 (.L_HI(net193));
 sg13g2_tiehi _09703__194 (.L_HI(net194));
 sg13g2_tiehi _09702__195 (.L_HI(net195));
 sg13g2_tiehi _09701__196 (.L_HI(net196));
 sg13g2_tiehi _09700__197 (.L_HI(net197));
 sg13g2_tiehi _09699__198 (.L_HI(net198));
 sg13g2_tiehi _09698__199 (.L_HI(net199));
 sg13g2_tiehi _09697__200 (.L_HI(net200));
 sg13g2_tiehi _09696__201 (.L_HI(net201));
 sg13g2_tiehi _09695__202 (.L_HI(net202));
 sg13g2_tiehi _09694__203 (.L_HI(net203));
 sg13g2_tiehi _09693__204 (.L_HI(net204));
 sg13g2_tiehi _09692__205 (.L_HI(net205));
 sg13g2_tiehi _09691__206 (.L_HI(net206));
 sg13g2_tiehi _09690__207 (.L_HI(net207));
 sg13g2_tiehi _09689__208 (.L_HI(net208));
 sg13g2_tiehi _09688__209 (.L_HI(net209));
 sg13g2_tiehi _09687__210 (.L_HI(net210));
 sg13g2_tiehi _09686__211 (.L_HI(net211));
 sg13g2_tiehi _09685__212 (.L_HI(net212));
 sg13g2_tiehi _09684__213 (.L_HI(net213));
 sg13g2_tiehi _09683__214 (.L_HI(net214));
 sg13g2_tiehi _09682__215 (.L_HI(net215));
 sg13g2_tiehi _09681__216 (.L_HI(net216));
 sg13g2_tiehi _09680__217 (.L_HI(net217));
 sg13g2_tiehi _09679__218 (.L_HI(net218));
 sg13g2_tiehi _09678__219 (.L_HI(net219));
 sg13g2_tiehi _09677__220 (.L_HI(net220));
 sg13g2_tiehi _09676__221 (.L_HI(net221));
 sg13g2_tiehi _09675__222 (.L_HI(net222));
 sg13g2_tiehi _09674__223 (.L_HI(net223));
 sg13g2_tiehi _09673__224 (.L_HI(net224));
 sg13g2_tiehi _09672__225 (.L_HI(net225));
 sg13g2_tiehi _09671__226 (.L_HI(net226));
 sg13g2_tiehi _09670__227 (.L_HI(net227));
 sg13g2_tiehi _09669__228 (.L_HI(net228));
 sg13g2_tiehi _09668__229 (.L_HI(net229));
 sg13g2_tiehi _09667__230 (.L_HI(net230));
 sg13g2_tiehi _09666__231 (.L_HI(net231));
 sg13g2_tiehi _09665__232 (.L_HI(net232));
 sg13g2_tiehi _09664__233 (.L_HI(net233));
 sg13g2_tiehi _09663__234 (.L_HI(net234));
 sg13g2_tiehi _09662__235 (.L_HI(net235));
 sg13g2_tiehi _09661__236 (.L_HI(net236));
 sg13g2_tiehi _09660__237 (.L_HI(net237));
 sg13g2_tiehi _09659__238 (.L_HI(net238));
 sg13g2_tiehi _09658__239 (.L_HI(net239));
 sg13g2_tiehi _09657__240 (.L_HI(net240));
 sg13g2_tiehi _09656__241 (.L_HI(net241));
 sg13g2_tiehi _09655__242 (.L_HI(net242));
 sg13g2_tiehi _09654__243 (.L_HI(net243));
 sg13g2_tiehi _09653__244 (.L_HI(net244));
 sg13g2_tiehi _09652__245 (.L_HI(net245));
 sg13g2_tiehi _09651__246 (.L_HI(net246));
 sg13g2_tiehi _09650__247 (.L_HI(net247));
 sg13g2_tiehi _09649__248 (.L_HI(net248));
 sg13g2_tiehi _09648__249 (.L_HI(net249));
 sg13g2_tiehi _09647__250 (.L_HI(net250));
 sg13g2_tiehi _09646__251 (.L_HI(net251));
 sg13g2_tiehi _09645__252 (.L_HI(net252));
 sg13g2_tiehi _09644__253 (.L_HI(net253));
 sg13g2_tiehi _09643__254 (.L_HI(net254));
 sg13g2_tiehi _09642__255 (.L_HI(net255));
 sg13g2_tiehi _09641__256 (.L_HI(net256));
 sg13g2_tiehi _09640__257 (.L_HI(net257));
 sg13g2_tiehi _09639__258 (.L_HI(net258));
 sg13g2_tiehi _09638__259 (.L_HI(net259));
 sg13g2_tiehi _09637__260 (.L_HI(net260));
 sg13g2_tiehi _09636__261 (.L_HI(net261));
 sg13g2_tiehi _09635__262 (.L_HI(net262));
 sg13g2_tiehi _09634__263 (.L_HI(net263));
 sg13g2_tiehi _09633__264 (.L_HI(net264));
 sg13g2_tiehi _09632__265 (.L_HI(net265));
 sg13g2_tiehi _09631__266 (.L_HI(net266));
 sg13g2_tiehi _09630__267 (.L_HI(net267));
 sg13g2_tiehi _09629__268 (.L_HI(net268));
 sg13g2_tiehi _09628__269 (.L_HI(net269));
 sg13g2_tiehi _09627__270 (.L_HI(net270));
 sg13g2_tiehi _09626__271 (.L_HI(net271));
 sg13g2_tiehi _09625__272 (.L_HI(net272));
 sg13g2_tiehi _09624__273 (.L_HI(net273));
 sg13g2_tiehi _09623__274 (.L_HI(net274));
 sg13g2_tiehi _09622__275 (.L_HI(net275));
 sg13g2_tiehi _09621__276 (.L_HI(net276));
 sg13g2_tiehi _09620__277 (.L_HI(net277));
 sg13g2_tiehi _09619__278 (.L_HI(net278));
 sg13g2_tiehi _09618__279 (.L_HI(net279));
 sg13g2_tiehi _09617__280 (.L_HI(net280));
 sg13g2_tiehi _09616__281 (.L_HI(net281));
 sg13g2_tiehi _09615__282 (.L_HI(net282));
 sg13g2_tiehi _09614__283 (.L_HI(net283));
 sg13g2_tiehi _09613__284 (.L_HI(net284));
 sg13g2_tiehi _09612__285 (.L_HI(net285));
 sg13g2_tiehi _09611__286 (.L_HI(net286));
 sg13g2_tiehi _09610__287 (.L_HI(net287));
 sg13g2_tiehi _09609__288 (.L_HI(net288));
 sg13g2_tiehi _09608__289 (.L_HI(net289));
 sg13g2_tiehi _09607__290 (.L_HI(net290));
 sg13g2_tiehi _09606__291 (.L_HI(net291));
 sg13g2_tiehi _09605__292 (.L_HI(net292));
 sg13g2_tiehi _09604__293 (.L_HI(net293));
 sg13g2_tiehi _09603__294 (.L_HI(net294));
 sg13g2_tiehi _09602__295 (.L_HI(net295));
 sg13g2_tiehi _09601__296 (.L_HI(net296));
 sg13g2_tiehi _09600__297 (.L_HI(net297));
 sg13g2_tiehi _09599__298 (.L_HI(net298));
 sg13g2_tiehi _09598__299 (.L_HI(net299));
 sg13g2_tiehi _09597__300 (.L_HI(net300));
 sg13g2_tiehi _09596__301 (.L_HI(net301));
 sg13g2_tiehi _09595__302 (.L_HI(net302));
 sg13g2_tiehi _09594__303 (.L_HI(net303));
 sg13g2_tiehi _09593__304 (.L_HI(net304));
 sg13g2_tiehi _09592__305 (.L_HI(net305));
 sg13g2_tiehi _09591__306 (.L_HI(net306));
 sg13g2_tiehi _09590__307 (.L_HI(net307));
 sg13g2_tiehi _09589__308 (.L_HI(net308));
 sg13g2_tiehi _09588__309 (.L_HI(net309));
 sg13g2_tiehi _09587__310 (.L_HI(net310));
 sg13g2_tiehi _09586__311 (.L_HI(net311));
 sg13g2_tiehi _09585__312 (.L_HI(net312));
 sg13g2_tiehi _09584__313 (.L_HI(net313));
 sg13g2_tiehi _09583__314 (.L_HI(net314));
 sg13g2_tiehi _09582__315 (.L_HI(net315));
 sg13g2_tiehi _09581__316 (.L_HI(net316));
 sg13g2_tiehi _09580__317 (.L_HI(net317));
 sg13g2_tiehi _09579__318 (.L_HI(net318));
 sg13g2_tiehi _09578__319 (.L_HI(net319));
 sg13g2_tiehi _09577__320 (.L_HI(net320));
 sg13g2_tiehi _09576__321 (.L_HI(net321));
 sg13g2_tiehi _09575__322 (.L_HI(net322));
 sg13g2_tiehi _09574__323 (.L_HI(net323));
 sg13g2_tiehi _09573__324 (.L_HI(net324));
 sg13g2_tiehi _09572__325 (.L_HI(net325));
 sg13g2_tiehi _09571__326 (.L_HI(net326));
 sg13g2_tiehi _09570__327 (.L_HI(net327));
 sg13g2_tiehi _09569__328 (.L_HI(net328));
 sg13g2_tiehi _09568__329 (.L_HI(net329));
 sg13g2_tiehi _09567__330 (.L_HI(net330));
 sg13g2_tiehi _09566__331 (.L_HI(net331));
 sg13g2_tiehi _09565__332 (.L_HI(net332));
 sg13g2_tiehi _09564__333 (.L_HI(net333));
 sg13g2_tiehi _09563__334 (.L_HI(net334));
 sg13g2_tiehi _09562__335 (.L_HI(net335));
 sg13g2_tiehi _09561__336 (.L_HI(net336));
 sg13g2_tiehi _09560__337 (.L_HI(net337));
 sg13g2_tiehi _09559__338 (.L_HI(net338));
 sg13g2_tiehi _09558__339 (.L_HI(net339));
 sg13g2_tiehi _09557__340 (.L_HI(net340));
 sg13g2_tiehi _09556__341 (.L_HI(net341));
 sg13g2_tiehi _09555__342 (.L_HI(net342));
 sg13g2_tiehi _09554__343 (.L_HI(net343));
 sg13g2_tiehi _09553__344 (.L_HI(net344));
 sg13g2_tiehi _09552__345 (.L_HI(net345));
 sg13g2_tiehi _09551__346 (.L_HI(net346));
 sg13g2_tiehi _09550__347 (.L_HI(net347));
 sg13g2_tiehi _09549__348 (.L_HI(net348));
 sg13g2_tiehi _09548__349 (.L_HI(net349));
 sg13g2_tiehi _09547__350 (.L_HI(net350));
 sg13g2_tiehi _09546__351 (.L_HI(net351));
 sg13g2_tiehi _09545__352 (.L_HI(net352));
 sg13g2_tiehi _09544__353 (.L_HI(net353));
 sg13g2_tiehi _09543__354 (.L_HI(net354));
 sg13g2_tiehi _09542__355 (.L_HI(net355));
 sg13g2_tiehi _09541__356 (.L_HI(net356));
 sg13g2_tiehi _09540__357 (.L_HI(net357));
 sg13g2_tiehi _09539__358 (.L_HI(net358));
 sg13g2_tiehi _09538__359 (.L_HI(net359));
 sg13g2_tiehi _09537__360 (.L_HI(net360));
 sg13g2_tiehi _09536__361 (.L_HI(net361));
 sg13g2_tiehi _09535__362 (.L_HI(net362));
 sg13g2_tiehi _09534__363 (.L_HI(net363));
 sg13g2_tiehi _09533__364 (.L_HI(net364));
 sg13g2_tiehi _09532__365 (.L_HI(net365));
 sg13g2_tiehi _09531__366 (.L_HI(net366));
 sg13g2_tiehi _09530__367 (.L_HI(net367));
 sg13g2_tiehi _09529__368 (.L_HI(net368));
 sg13g2_tiehi _09528__369 (.L_HI(net369));
 sg13g2_tiehi _09527__370 (.L_HI(net370));
 sg13g2_tiehi _09526__371 (.L_HI(net371));
 sg13g2_tiehi _09525__372 (.L_HI(net372));
 sg13g2_tiehi _09524__373 (.L_HI(net373));
 sg13g2_tiehi _09523__374 (.L_HI(net374));
 sg13g2_tiehi _09522__375 (.L_HI(net375));
 sg13g2_tiehi _09521__376 (.L_HI(net376));
 sg13g2_tiehi _09520__377 (.L_HI(net377));
 sg13g2_tiehi _09519__378 (.L_HI(net378));
 sg13g2_tiehi _09518__379 (.L_HI(net379));
 sg13g2_tiehi _09517__380 (.L_HI(net380));
 sg13g2_tiehi _09516__381 (.L_HI(net381));
 sg13g2_tiehi _09515__382 (.L_HI(net382));
 sg13g2_tiehi _09514__383 (.L_HI(net383));
 sg13g2_tiehi _09513__384 (.L_HI(net384));
 sg13g2_tiehi _09512__385 (.L_HI(net385));
 sg13g2_tiehi _09511__386 (.L_HI(net386));
 sg13g2_tiehi _09510__387 (.L_HI(net387));
 sg13g2_tiehi _09509__388 (.L_HI(net388));
 sg13g2_tiehi _09508__389 (.L_HI(net389));
 sg13g2_tiehi _09507__390 (.L_HI(net390));
 sg13g2_tiehi _09506__391 (.L_HI(net391));
 sg13g2_tiehi _09505__392 (.L_HI(net392));
 sg13g2_tiehi _09504__393 (.L_HI(net393));
 sg13g2_tiehi _09503__394 (.L_HI(net394));
 sg13g2_tiehi _09502__395 (.L_HI(net395));
 sg13g2_tiehi _09501__396 (.L_HI(net396));
 sg13g2_tiehi _09500__397 (.L_HI(net397));
 sg13g2_tiehi _09499__398 (.L_HI(net398));
 sg13g2_tiehi _09498__399 (.L_HI(net399));
 sg13g2_tiehi _09497__400 (.L_HI(net400));
 sg13g2_tiehi _09496__401 (.L_HI(net401));
 sg13g2_tiehi _09495__402 (.L_HI(net402));
 sg13g2_tiehi _09494__403 (.L_HI(net403));
 sg13g2_tiehi _09493__404 (.L_HI(net404));
 sg13g2_tiehi _09492__405 (.L_HI(net405));
 sg13g2_tiehi _09491__406 (.L_HI(net406));
 sg13g2_tiehi _09490__407 (.L_HI(net407));
 sg13g2_tiehi _09489__408 (.L_HI(net408));
 sg13g2_tiehi _09488__409 (.L_HI(net409));
 sg13g2_tiehi _09487__410 (.L_HI(net410));
 sg13g2_tiehi _09486__411 (.L_HI(net411));
 sg13g2_tiehi _09485__412 (.L_HI(net412));
 sg13g2_tiehi _09484__413 (.L_HI(net413));
 sg13g2_tiehi _09483__414 (.L_HI(net414));
 sg13g2_tiehi _09482__415 (.L_HI(net415));
 sg13g2_tiehi _09481__416 (.L_HI(net416));
 sg13g2_tiehi _09480__417 (.L_HI(net417));
 sg13g2_tiehi _09479__418 (.L_HI(net418));
 sg13g2_tiehi _09478__419 (.L_HI(net419));
 sg13g2_tiehi _09477__420 (.L_HI(net420));
 sg13g2_tiehi _09476__421 (.L_HI(net421));
 sg13g2_tiehi _09475__422 (.L_HI(net422));
 sg13g2_tiehi _09474__423 (.L_HI(net423));
 sg13g2_tiehi _09473__424 (.L_HI(net424));
 sg13g2_tiehi _09472__425 (.L_HI(net425));
 sg13g2_tiehi _09471__426 (.L_HI(net426));
 sg13g2_tiehi _09470__427 (.L_HI(net427));
 sg13g2_tiehi _09469__428 (.L_HI(net428));
 sg13g2_tiehi _09468__429 (.L_HI(net429));
 sg13g2_tiehi _09467__430 (.L_HI(net430));
 sg13g2_tiehi _09466__431 (.L_HI(net431));
 sg13g2_tiehi _09465__432 (.L_HI(net432));
 sg13g2_tiehi _09464__433 (.L_HI(net433));
 sg13g2_tiehi _09463__434 (.L_HI(net434));
 sg13g2_tiehi _09462__435 (.L_HI(net435));
 sg13g2_tiehi _09461__436 (.L_HI(net436));
 sg13g2_tiehi _09460__437 (.L_HI(net437));
 sg13g2_tiehi _09459__438 (.L_HI(net438));
 sg13g2_tiehi _09458__439 (.L_HI(net439));
 sg13g2_tiehi _09457__440 (.L_HI(net440));
 sg13g2_tiehi _09456__441 (.L_HI(net441));
 sg13g2_tiehi _09455__442 (.L_HI(net442));
 sg13g2_tiehi _09454__443 (.L_HI(net443));
 sg13g2_tiehi _09453__444 (.L_HI(net444));
 sg13g2_tiehi _09452__445 (.L_HI(net445));
 sg13g2_tiehi _09451__446 (.L_HI(net446));
 sg13g2_tiehi _09450__447 (.L_HI(net447));
 sg13g2_tiehi _09449__448 (.L_HI(net448));
 sg13g2_tiehi _09448__449 (.L_HI(net449));
 sg13g2_tiehi _09447__450 (.L_HI(net450));
 sg13g2_tiehi _09446__451 (.L_HI(net451));
 sg13g2_tiehi _09445__452 (.L_HI(net452));
 sg13g2_tiehi _09444__453 (.L_HI(net453));
 sg13g2_tiehi _09443__454 (.L_HI(net454));
 sg13g2_tiehi _09442__455 (.L_HI(net455));
 sg13g2_tiehi _09441__456 (.L_HI(net456));
 sg13g2_tiehi _09440__457 (.L_HI(net457));
 sg13g2_tiehi _09439__458 (.L_HI(net458));
 sg13g2_tiehi _09438__459 (.L_HI(net459));
 sg13g2_tiehi _09437__460 (.L_HI(net460));
 sg13g2_tiehi _09436__461 (.L_HI(net461));
 sg13g2_tiehi _09435__462 (.L_HI(net462));
 sg13g2_tiehi _09434__463 (.L_HI(net463));
 sg13g2_tiehi _09433__464 (.L_HI(net464));
 sg13g2_tiehi _09432__465 (.L_HI(net465));
 sg13g2_tiehi _09431__466 (.L_HI(net466));
 sg13g2_tiehi _09430__467 (.L_HI(net467));
 sg13g2_tiehi _09429__468 (.L_HI(net468));
 sg13g2_tiehi _09428__469 (.L_HI(net469));
 sg13g2_tiehi _09427__470 (.L_HI(net470));
 sg13g2_tiehi _09426__471 (.L_HI(net471));
 sg13g2_tiehi _09425__472 (.L_HI(net472));
 sg13g2_tiehi _09424__473 (.L_HI(net473));
 sg13g2_tiehi _09423__474 (.L_HI(net474));
 sg13g2_tiehi _09422__475 (.L_HI(net475));
 sg13g2_tiehi _09421__476 (.L_HI(net476));
 sg13g2_tiehi _09420__477 (.L_HI(net477));
 sg13g2_tiehi _09419__478 (.L_HI(net478));
 sg13g2_tiehi _09418__479 (.L_HI(net479));
 sg13g2_tiehi _09417__480 (.L_HI(net480));
 sg13g2_tiehi _09416__481 (.L_HI(net481));
 sg13g2_tiehi _09415__482 (.L_HI(net482));
 sg13g2_tiehi _09414__483 (.L_HI(net483));
 sg13g2_tiehi _09413__484 (.L_HI(net484));
 sg13g2_tiehi _09412__485 (.L_HI(net485));
 sg13g2_tiehi _09411__486 (.L_HI(net486));
 sg13g2_tiehi _09410__487 (.L_HI(net487));
 sg13g2_tiehi _09409__488 (.L_HI(net488));
 sg13g2_tiehi _09408__489 (.L_HI(net489));
 sg13g2_tiehi _09407__490 (.L_HI(net490));
 sg13g2_tiehi _09406__491 (.L_HI(net491));
 sg13g2_tiehi _09405__492 (.L_HI(net492));
 sg13g2_tiehi _09404__493 (.L_HI(net493));
 sg13g2_tiehi _09403__494 (.L_HI(net494));
 sg13g2_tiehi _09402__495 (.L_HI(net495));
 sg13g2_tiehi _09401__496 (.L_HI(net496));
 sg13g2_tiehi _09400__497 (.L_HI(net497));
 sg13g2_tiehi _09399__498 (.L_HI(net498));
 sg13g2_tiehi _09398__499 (.L_HI(net499));
 sg13g2_tiehi _09397__500 (.L_HI(net500));
 sg13g2_tiehi _09396__501 (.L_HI(net501));
 sg13g2_tiehi _09395__502 (.L_HI(net502));
 sg13g2_tiehi _09394__503 (.L_HI(net503));
 sg13g2_tiehi _09393__504 (.L_HI(net504));
 sg13g2_tiehi _09392__505 (.L_HI(net505));
 sg13g2_tiehi _09391__506 (.L_HI(net506));
 sg13g2_tiehi _09390__507 (.L_HI(net507));
 sg13g2_tiehi _09389__508 (.L_HI(net508));
 sg13g2_tiehi _09388__509 (.L_HI(net509));
 sg13g2_tiehi _10569__510 (.L_HI(net510));
 sg13g2_tiehi _09387__511 (.L_HI(net511));
 sg13g2_tiehi _10558__512 (.L_HI(net512));
 sg13g2_tiehi _09386__513 (.L_HI(net513));
 sg13g2_tiehi _10576__514 (.L_HI(net514));
 sg13g2_tiehi _09385__515 (.L_HI(net515));
 sg13g2_tiehi _10557__516 (.L_HI(net516));
 sg13g2_tiehi _09384__517 (.L_HI(net517));
 sg13g2_tiehi _09383__518 (.L_HI(net518));
 sg13g2_tiehi _09382__519 (.L_HI(net519));
 sg13g2_tiehi _09381__520 (.L_HI(net520));
 sg13g2_tiehi _09380__521 (.L_HI(net521));
 sg13g2_tiehi _09379__522 (.L_HI(net522));
 sg13g2_tiehi _09378__523 (.L_HI(net523));
 sg13g2_tiehi _09377__524 (.L_HI(net524));
 sg13g2_tiehi _09376__525 (.L_HI(net525));
 sg13g2_tiehi _09375__526 (.L_HI(net526));
 sg13g2_tiehi _09374__527 (.L_HI(net527));
 sg13g2_tiehi _09373__528 (.L_HI(net528));
 sg13g2_tiehi _09372__529 (.L_HI(net529));
 sg13g2_tiehi _09371__530 (.L_HI(net530));
 sg13g2_tiehi _09370__531 (.L_HI(net531));
 sg13g2_tiehi _09369__532 (.L_HI(net532));
 sg13g2_tiehi _09368__533 (.L_HI(net533));
 sg13g2_tiehi _09367__534 (.L_HI(net534));
 sg13g2_tiehi _09366__535 (.L_HI(net535));
 sg13g2_tiehi _09365__536 (.L_HI(net536));
 sg13g2_tiehi _09364__537 (.L_HI(net537));
 sg13g2_tiehi _09363__538 (.L_HI(net538));
 sg13g2_tiehi _09362__539 (.L_HI(net539));
 sg13g2_tiehi _09361__540 (.L_HI(net540));
 sg13g2_tiehi _09360__541 (.L_HI(net541));
 sg13g2_tiehi _09359__542 (.L_HI(net542));
 sg13g2_tiehi _09358__543 (.L_HI(net543));
 sg13g2_tiehi _09357__544 (.L_HI(net544));
 sg13g2_tiehi _09356__545 (.L_HI(net545));
 sg13g2_tiehi _09355__546 (.L_HI(net546));
 sg13g2_tiehi _09354__547 (.L_HI(net547));
 sg13g2_tiehi _09353__548 (.L_HI(net548));
 sg13g2_tiehi _09352__549 (.L_HI(net549));
 sg13g2_tiehi _09351__550 (.L_HI(net550));
 sg13g2_tiehi _09350__551 (.L_HI(net551));
 sg13g2_tiehi _09349__552 (.L_HI(net552));
 sg13g2_tiehi _09348__553 (.L_HI(net553));
 sg13g2_tiehi _09347__554 (.L_HI(net554));
 sg13g2_tiehi _09346__555 (.L_HI(net555));
 sg13g2_tiehi _09345__556 (.L_HI(net556));
 sg13g2_tiehi _09344__557 (.L_HI(net557));
 sg13g2_tiehi _09343__558 (.L_HI(net558));
 sg13g2_tiehi _09342__559 (.L_HI(net559));
 sg13g2_tiehi _09341__560 (.L_HI(net560));
 sg13g2_tiehi _09340__561 (.L_HI(net561));
 sg13g2_tiehi _09339__562 (.L_HI(net562));
 sg13g2_tiehi _09338__563 (.L_HI(net563));
 sg13g2_tiehi _09337__564 (.L_HI(net564));
 sg13g2_tiehi _09336__565 (.L_HI(net565));
 sg13g2_tiehi _09335__566 (.L_HI(net566));
 sg13g2_tiehi _09334__567 (.L_HI(net567));
 sg13g2_tiehi _09333__568 (.L_HI(net568));
 sg13g2_tiehi _09332__569 (.L_HI(net569));
 sg13g2_tiehi _09331__570 (.L_HI(net570));
 sg13g2_tiehi _09330__571 (.L_HI(net571));
 sg13g2_tiehi _09329__572 (.L_HI(net572));
 sg13g2_tiehi _09328__573 (.L_HI(net573));
 sg13g2_tiehi _09327__574 (.L_HI(net574));
 sg13g2_tiehi _09326__575 (.L_HI(net575));
 sg13g2_tiehi _09325__576 (.L_HI(net576));
 sg13g2_tiehi _09324__577 (.L_HI(net577));
 sg13g2_tiehi _09323__578 (.L_HI(net578));
 sg13g2_tiehi _09322__579 (.L_HI(net579));
 sg13g2_tiehi _09321__580 (.L_HI(net580));
 sg13g2_tiehi _09320__581 (.L_HI(net581));
 sg13g2_tiehi _09319__582 (.L_HI(net582));
 sg13g2_tiehi _09318__583 (.L_HI(net583));
 sg13g2_tiehi _09317__584 (.L_HI(net584));
 sg13g2_tiehi _09316__585 (.L_HI(net585));
 sg13g2_tiehi _09315__586 (.L_HI(net586));
 sg13g2_tiehi _09314__587 (.L_HI(net587));
 sg13g2_tiehi _09313__588 (.L_HI(net588));
 sg13g2_tiehi _09312__589 (.L_HI(net589));
 sg13g2_tiehi _09311__590 (.L_HI(net590));
 sg13g2_tiehi _09310__591 (.L_HI(net591));
 sg13g2_tiehi _09309__592 (.L_HI(net592));
 sg13g2_tiehi _09308__593 (.L_HI(net593));
 sg13g2_tiehi _09307__594 (.L_HI(net594));
 sg13g2_tiehi _09306__595 (.L_HI(net595));
 sg13g2_tiehi _09305__596 (.L_HI(net596));
 sg13g2_tiehi _09304__597 (.L_HI(net597));
 sg13g2_tiehi _09303__598 (.L_HI(net598));
 sg13g2_tiehi _09302__599 (.L_HI(net599));
 sg13g2_tiehi _09301__600 (.L_HI(net600));
 sg13g2_tiehi _09300__601 (.L_HI(net601));
 sg13g2_tiehi _09299__602 (.L_HI(net602));
 sg13g2_tiehi _09298__603 (.L_HI(net603));
 sg13g2_tiehi _09297__604 (.L_HI(net604));
 sg13g2_tiehi _09296__605 (.L_HI(net605));
 sg13g2_tiehi _09295__606 (.L_HI(net606));
 sg13g2_tiehi _09294__607 (.L_HI(net607));
 sg13g2_tiehi _09293__608 (.L_HI(net608));
 sg13g2_tiehi _09292__609 (.L_HI(net609));
 sg13g2_tiehi _09291__610 (.L_HI(net610));
 sg13g2_tiehi _09290__611 (.L_HI(net611));
 sg13g2_tiehi _09289__612 (.L_HI(net612));
 sg13g2_tiehi _09288__613 (.L_HI(net613));
 sg13g2_tiehi _09276__614 (.L_HI(net614));
 sg13g2_tiehi _09275__615 (.L_HI(net615));
 sg13g2_tiehi _09274__616 (.L_HI(net616));
 sg13g2_tiehi _09273__617 (.L_HI(net617));
 sg13g2_tiehi _09272__618 (.L_HI(net618));
 sg13g2_tiehi _09271__619 (.L_HI(net619));
 sg13g2_tiehi _09270__620 (.L_HI(net620));
 sg13g2_tiehi _09269__621 (.L_HI(net621));
 sg13g2_tiehi _09268__622 (.L_HI(net622));
 sg13g2_tiehi _09267__623 (.L_HI(net623));
 sg13g2_tiehi _09266__624 (.L_HI(net624));
 sg13g2_tiehi _09265__625 (.L_HI(net625));
 sg13g2_tiehi _09264__626 (.L_HI(net626));
 sg13g2_tiehi _09263__627 (.L_HI(net627));
 sg13g2_tiehi _09262__628 (.L_HI(net628));
 sg13g2_tiehi _09261__629 (.L_HI(net629));
 sg13g2_tiehi _09260__630 (.L_HI(net630));
 sg13g2_tiehi _09259__631 (.L_HI(net631));
 sg13g2_tiehi _09258__632 (.L_HI(net632));
 sg13g2_tiehi _09257__633 (.L_HI(net633));
 sg13g2_tiehi _09256__634 (.L_HI(net634));
 sg13g2_tiehi _09255__635 (.L_HI(net635));
 sg13g2_tiehi _09254__636 (.L_HI(net636));
 sg13g2_tiehi _09253__637 (.L_HI(net637));
 sg13g2_tiehi _09252__638 (.L_HI(net638));
 sg13g2_tiehi _09251__639 (.L_HI(net639));
 sg13g2_tiehi _09250__640 (.L_HI(net640));
 sg13g2_tiehi _09249__641 (.L_HI(net641));
 sg13g2_tiehi _09248__642 (.L_HI(net642));
 sg13g2_tiehi _09247__643 (.L_HI(net643));
 sg13g2_tiehi _09246__644 (.L_HI(net644));
 sg13g2_tiehi _09245__645 (.L_HI(net645));
 sg13g2_tiehi _09244__646 (.L_HI(net646));
 sg13g2_tiehi _09243__647 (.L_HI(net647));
 sg13g2_tiehi _09242__648 (.L_HI(net648));
 sg13g2_tiehi _09241__649 (.L_HI(net649));
 sg13g2_tiehi _09240__650 (.L_HI(net650));
 sg13g2_tiehi _09239__651 (.L_HI(net651));
 sg13g2_tiehi _09238__652 (.L_HI(net652));
 sg13g2_tiehi _09237__653 (.L_HI(net653));
 sg13g2_tiehi _09236__654 (.L_HI(net654));
 sg13g2_tiehi _09235__655 (.L_HI(net655));
 sg13g2_tiehi _09234__656 (.L_HI(net656));
 sg13g2_tiehi _09233__657 (.L_HI(net657));
 sg13g2_tiehi _09232__658 (.L_HI(net658));
 sg13g2_tiehi _09231__659 (.L_HI(net659));
 sg13g2_tiehi _09230__660 (.L_HI(net660));
 sg13g2_tiehi _09229__661 (.L_HI(net661));
 sg13g2_tiehi _09228__662 (.L_HI(net662));
 sg13g2_tiehi _09227__663 (.L_HI(net663));
 sg13g2_tiehi _09226__664 (.L_HI(net664));
 sg13g2_tiehi _09225__665 (.L_HI(net665));
 sg13g2_tiehi _09224__666 (.L_HI(net666));
 sg13g2_tiehi _09223__667 (.L_HI(net667));
 sg13g2_tiehi _09222__668 (.L_HI(net668));
 sg13g2_tiehi _09221__669 (.L_HI(net669));
 sg13g2_tiehi _09220__670 (.L_HI(net670));
 sg13g2_tiehi _09219__671 (.L_HI(net671));
 sg13g2_tiehi _09218__672 (.L_HI(net672));
 sg13g2_tiehi _09217__673 (.L_HI(net673));
 sg13g2_tiehi _09216__674 (.L_HI(net674));
 sg13g2_tiehi _09215__675 (.L_HI(net675));
 sg13g2_tiehi _10568__676 (.L_HI(net676));
 sg13g2_tiehi _10556__677 (.L_HI(net677));
 sg13g2_tiehi _10575__678 (.L_HI(net678));
 sg13g2_tiehi _10555__679 (.L_HI(net679));
 sg13g2_tiehi _10567__680 (.L_HI(net680));
 sg13g2_tiehi _10554__681 (.L_HI(net681));
 sg13g2_tiehi _10574__682 (.L_HI(net682));
 sg13g2_tiehi _10553__683 (.L_HI(net683));
 sg13g2_tiehi _10566__684 (.L_HI(net684));
 sg13g2_tiehi _10552__685 (.L_HI(net685));
 sg13g2_tiehi _10572__686 (.L_HI(net686));
 sg13g2_tiehi _10551__687 (.L_HI(net687));
 sg13g2_tiehi _10565__688 (.L_HI(net688));
 sg13g2_tiehi _10550__689 (.L_HI(net689));
 sg13g2_tiehi _10573__690 (.L_HI(net690));
 sg13g2_tiehi _10549__691 (.L_HI(net691));
 sg13g2_tiehi _10564__692 (.L_HI(net692));
 sg13g2_tiehi _10548__693 (.L_HI(net693));
 sg13g2_tiehi _10579__694 (.L_HI(net694));
 sg13g2_tiehi _10547__695 (.L_HI(net695));
 sg13g2_tiehi _10563__696 (.L_HI(net696));
 sg13g2_tiehi _10546__697 (.L_HI(net697));
 sg13g2_tiehi _10571__698 (.L_HI(net698));
 sg13g2_tiehi _10545__699 (.L_HI(net699));
 sg13g2_tiehi _10562__700 (.L_HI(net700));
 sg13g2_tiehi _10544__701 (.L_HI(net701));
 sg13g2_tiehi _10578__702 (.L_HI(net702));
 sg13g2_tiehi _10543__703 (.L_HI(net703));
 sg13g2_tiehi _10561__704 (.L_HI(net704));
 sg13g2_tiehi _10542__705 (.L_HI(net705));
 sg13g2_tiehi _10570__706 (.L_HI(net706));
 sg13g2_tiehi _10541__707 (.L_HI(net707));
 sg13g2_tiehi _10540__708 (.L_HI(net708));
 sg13g2_tiehi _10537__709 (.L_HI(net709));
 sg13g2_tiehi _10536__710 (.L_HI(net710));
 sg13g2_tiehi _10535__711 (.L_HI(net711));
 sg13g2_tiehi _10534__712 (.L_HI(net712));
 sg13g2_tiehi _10533__713 (.L_HI(net713));
 sg13g2_tiehi _10532__714 (.L_HI(net714));
 sg13g2_tiehi _10531__715 (.L_HI(net715));
 sg13g2_tiehi _10530__716 (.L_HI(net716));
 sg13g2_tiehi _10529__717 (.L_HI(net717));
 sg13g2_tiehi _10528__718 (.L_HI(net718));
 sg13g2_tiehi _10527__719 (.L_HI(net719));
 sg13g2_tiehi _10526__720 (.L_HI(net720));
 sg13g2_tiehi _10525__721 (.L_HI(net721));
 sg13g2_tiehi _10524__722 (.L_HI(net722));
 sg13g2_tiehi _10523__723 (.L_HI(net723));
 sg13g2_tiehi _10522__724 (.L_HI(net724));
 sg13g2_tiehi _10521__725 (.L_HI(net725));
 sg13g2_tiehi _10520__726 (.L_HI(net726));
 sg13g2_tiehi _10519__727 (.L_HI(net727));
 sg13g2_tiehi _10518__728 (.L_HI(net728));
 sg13g2_tiehi _10517__729 (.L_HI(net729));
 sg13g2_tiehi _10516__730 (.L_HI(net730));
 sg13g2_tiehi _10515__731 (.L_HI(net731));
 sg13g2_tiehi _10514__732 (.L_HI(net732));
 sg13g2_tiehi _10513__733 (.L_HI(net733));
 sg13g2_tiehi _10512__734 (.L_HI(net734));
 sg13g2_tiehi _10511__735 (.L_HI(net735));
 sg13g2_tiehi _10510__736 (.L_HI(net736));
 sg13g2_tiehi _10509__737 (.L_HI(net737));
 sg13g2_tiehi _10508__738 (.L_HI(net738));
 sg13g2_tiehi _10507__739 (.L_HI(net739));
 sg13g2_tiehi _10506__740 (.L_HI(net740));
 sg13g2_tiehi _10505__741 (.L_HI(net741));
 sg13g2_tiehi _10504__742 (.L_HI(net742));
 sg13g2_tiehi _10503__743 (.L_HI(net743));
 sg13g2_tiehi _10502__744 (.L_HI(net744));
 sg13g2_tiehi _10501__745 (.L_HI(net745));
 sg13g2_tiehi _10500__746 (.L_HI(net746));
 sg13g2_tiehi _10499__747 (.L_HI(net747));
 sg13g2_tiehi _10498__748 (.L_HI(net748));
 sg13g2_tiehi _10497__749 (.L_HI(net749));
 sg13g2_tiehi _10496__750 (.L_HI(net750));
 sg13g2_tiehi _10494__751 (.L_HI(net751));
 sg13g2_tiehi _10493__752 (.L_HI(net752));
 sg13g2_tiehi _10492__753 (.L_HI(net753));
 sg13g2_tiehi _10491__754 (.L_HI(net754));
 sg13g2_tiehi _10490__755 (.L_HI(net755));
 sg13g2_tiehi _10489__756 (.L_HI(net756));
 sg13g2_tiehi _10488__757 (.L_HI(net757));
 sg13g2_tiehi _10487__758 (.L_HI(net758));
 sg13g2_tiehi _10486__759 (.L_HI(net759));
 sg13g2_tiehi _10485__760 (.L_HI(net760));
 sg13g2_tiehi _10484__761 (.L_HI(net761));
 sg13g2_tiehi _10483__762 (.L_HI(net762));
 sg13g2_tiehi _10482__763 (.L_HI(net763));
 sg13g2_tiehi _10481__764 (.L_HI(net764));
 sg13g2_tiehi _10480__765 (.L_HI(net765));
 sg13g2_tiehi _10479__766 (.L_HI(net766));
 sg13g2_tiehi _10478__767 (.L_HI(net767));
 sg13g2_tiehi _10477__768 (.L_HI(net768));
 sg13g2_tiehi _10476__769 (.L_HI(net769));
 sg13g2_tiehi _10475__770 (.L_HI(net770));
 sg13g2_tiehi _10474__771 (.L_HI(net771));
 sg13g2_tiehi _10473__772 (.L_HI(net772));
 sg13g2_tiehi _10472__773 (.L_HI(net773));
 sg13g2_tiehi _10471__774 (.L_HI(net774));
 sg13g2_tiehi _10470__775 (.L_HI(net775));
 sg13g2_tiehi _10469__776 (.L_HI(net776));
 sg13g2_tiehi _10468__777 (.L_HI(net777));
 sg13g2_tiehi _10467__778 (.L_HI(net778));
 sg13g2_tiehi _10466__779 (.L_HI(net779));
 sg13g2_tiehi _10465__780 (.L_HI(net780));
 sg13g2_tiehi _10464__781 (.L_HI(net781));
 sg13g2_tiehi _10463__782 (.L_HI(net782));
 sg13g2_tiehi _10462__783 (.L_HI(net783));
 sg13g2_tiehi _10461__784 (.L_HI(net784));
 sg13g2_tiehi _10460__785 (.L_HI(net785));
 sg13g2_tiehi _10459__786 (.L_HI(net786));
 sg13g2_tiehi _10458__787 (.L_HI(net787));
 sg13g2_tiehi _10457__788 (.L_HI(net788));
 sg13g2_tiehi _10456__789 (.L_HI(net789));
 sg13g2_tiehi _10455__790 (.L_HI(net790));
 sg13g2_tiehi _10454__791 (.L_HI(net791));
 sg13g2_tiehi _10453__792 (.L_HI(net792));
 sg13g2_tiehi _10452__793 (.L_HI(net793));
 sg13g2_tiehi _10451__794 (.L_HI(net794));
 sg13g2_tiehi _10450__795 (.L_HI(net795));
 sg13g2_tiehi _10449__796 (.L_HI(net796));
 sg13g2_tiehi _10448__797 (.L_HI(net797));
 sg13g2_tiehi _10447__798 (.L_HI(net798));
 sg13g2_tiehi _10446__799 (.L_HI(net799));
 sg13g2_tiehi _10445__800 (.L_HI(net800));
 sg13g2_tiehi _10444__801 (.L_HI(net801));
 sg13g2_tiehi _10443__802 (.L_HI(net802));
 sg13g2_tiehi _10442__803 (.L_HI(net803));
 sg13g2_tiehi _10441__804 (.L_HI(net804));
 sg13g2_tiehi _10440__805 (.L_HI(net805));
 sg13g2_tiehi _10439__806 (.L_HI(net806));
 sg13g2_tiehi _10438__807 (.L_HI(net807));
 sg13g2_tiehi _10437__808 (.L_HI(net808));
 sg13g2_tiehi _10436__809 (.L_HI(net809));
 sg13g2_tiehi _10435__810 (.L_HI(net810));
 sg13g2_tiehi _10560__811 (.L_HI(net811));
 sg13g2_tiehi _10434__812 (.L_HI(net812));
 sg13g2_tiehi _10577__813 (.L_HI(net813));
 sg13g2_tiehi _10433__814 (.L_HI(net814));
 sg13g2_tiehi _10432__815 (.L_HI(net815));
 sg13g2_tiehi _10431__816 (.L_HI(net816));
 sg13g2_tiehi _10430__817 (.L_HI(net817));
 sg13g2_tiehi _10429__818 (.L_HI(net818));
 sg13g2_tiehi _10428__819 (.L_HI(net819));
 sg13g2_tiehi _10427__820 (.L_HI(net820));
 sg13g2_tiehi _10426__821 (.L_HI(net821));
 sg13g2_tiehi _10559__822 (.L_HI(net822));
 sg13g2_tiehi _10393__823 (.L_HI(net823));
 sg13g2_tiehi _10392__824 (.L_HI(net824));
 sg13g2_tiehi _10390__825 (.L_HI(net825));
 sg13g2_tiehi _10389__826 (.L_HI(net826));
 sg13g2_tiehi _10388__827 (.L_HI(net827));
 sg13g2_tiehi _10386__828 (.L_HI(net828));
 sg13g2_tiehi _10385__829 (.L_HI(net829));
 sg13g2_tiehi _10384__830 (.L_HI(net830));
 sg13g2_tiehi _10383__831 (.L_HI(net831));
 sg13g2_tiehi _10382__832 (.L_HI(net832));
 sg13g2_tiehi _10381__833 (.L_HI(net833));
 sg13g2_tiehi _10380__834 (.L_HI(net834));
 sg13g2_tiehi _10379__835 (.L_HI(net835));
 sg13g2_tiehi _10378__836 (.L_HI(net836));
 sg13g2_tiehi _10377__837 (.L_HI(net837));
 sg13g2_tiehi _10376__838 (.L_HI(net838));
 sg13g2_tiehi _10375__839 (.L_HI(net839));
 sg13g2_tiehi _10374__840 (.L_HI(net840));
 sg13g2_tiehi _10373__841 (.L_HI(net841));
 sg13g2_tiehi _10372__842 (.L_HI(net842));
 sg13g2_tiehi _10371__843 (.L_HI(net843));
 sg13g2_tiehi _10370__844 (.L_HI(net844));
 sg13g2_tiehi _10369__845 (.L_HI(net845));
 sg13g2_tiehi _10368__846 (.L_HI(net846));
 sg13g2_tiehi _10367__847 (.L_HI(net847));
 sg13g2_tiehi _10366__848 (.L_HI(net848));
 sg13g2_tiehi _10365__849 (.L_HI(net849));
 sg13g2_tiehi _10364__850 (.L_HI(net850));
 sg13g2_tiehi _10363__851 (.L_HI(net851));
 sg13g2_tiehi _10362__852 (.L_HI(net852));
 sg13g2_tiehi _10361__853 (.L_HI(net853));
 sg13g2_tiehi _10360__854 (.L_HI(net854));
 sg13g2_tiehi _10359__855 (.L_HI(net855));
 sg13g2_tiehi _10358__856 (.L_HI(net856));
 sg13g2_tiehi _10357__857 (.L_HI(net857));
 sg13g2_tiehi _10356__858 (.L_HI(net858));
 sg13g2_tiehi _10355__859 (.L_HI(net859));
 sg13g2_tiehi _10354__860 (.L_HI(net860));
 sg13g2_tiehi _10292__861 (.L_HI(net861));
 sg13g2_tiehi _10291__862 (.L_HI(net862));
 sg13g2_tiehi _10290__863 (.L_HI(net863));
 sg13g2_tiehi _10289__864 (.L_HI(net864));
 sg13g2_tiehi _10288__865 (.L_HI(net865));
 sg13g2_tiehi _10287__866 (.L_HI(net866));
 sg13g2_tiehi _10286__867 (.L_HI(net867));
 sg13g2_tiehi _10285__868 (.L_HI(net868));
 sg13g2_tiehi _10284__869 (.L_HI(net869));
 sg13g2_tiehi _10283__870 (.L_HI(net870));
 sg13g2_tiehi _10282__871 (.L_HI(net871));
 sg13g2_tiehi _10281__872 (.L_HI(net872));
 sg13g2_tiehi _10280__873 (.L_HI(net873));
 sg13g2_tiehi _10279__874 (.L_HI(net874));
 sg13g2_tiehi _10278__875 (.L_HI(net875));
 sg13g2_tiehi _10277__876 (.L_HI(net876));
 sg13g2_tiehi _10276__877 (.L_HI(net877));
 sg13g2_tiehi _10275__878 (.L_HI(net878));
 sg13g2_tiehi _10274__879 (.L_HI(net879));
 sg13g2_tiehi _10273__880 (.L_HI(net880));
 sg13g2_tiehi _10272__881 (.L_HI(net881));
 sg13g2_tiehi _10271__882 (.L_HI(net882));
 sg13g2_tiehi _10270__883 (.L_HI(net883));
 sg13g2_tiehi _10269__884 (.L_HI(net884));
 sg13g2_tiehi _10268__885 (.L_HI(net885));
 sg13g2_tiehi _10267__886 (.L_HI(net886));
 sg13g2_tiehi _10266__887 (.L_HI(net887));
 sg13g2_tiehi _10265__888 (.L_HI(net888));
 sg13g2_tiehi _10264__889 (.L_HI(net889));
 sg13g2_tiehi _10263__890 (.L_HI(net890));
 sg13g2_tiehi _10262__891 (.L_HI(net891));
 sg13g2_tiehi _10261__892 (.L_HI(net892));
 sg13g2_tiehi _10260__893 (.L_HI(net893));
 sg13g2_tiehi _10259__894 (.L_HI(net894));
 sg13g2_tiehi _10258__895 (.L_HI(net895));
 sg13g2_tiehi _10257__896 (.L_HI(net896));
 sg13g2_tiehi _10256__897 (.L_HI(net897));
 sg13g2_tiehi _10255__898 (.L_HI(net898));
 sg13g2_tiehi _10254__899 (.L_HI(net899));
 sg13g2_tiehi _10253__900 (.L_HI(net900));
 sg13g2_tiehi _10252__901 (.L_HI(net901));
 sg13g2_tiehi _10251__902 (.L_HI(net902));
 sg13g2_tiehi _10250__903 (.L_HI(net903));
 sg13g2_tiehi _10249__904 (.L_HI(net904));
 sg13g2_tiehi _10248__905 (.L_HI(net905));
 sg13g2_tiehi _10247__906 (.L_HI(net906));
 sg13g2_tiehi _10246__907 (.L_HI(net907));
 sg13g2_tiehi _10245__908 (.L_HI(net908));
 sg13g2_tiehi _10244__909 (.L_HI(net909));
 sg13g2_tiehi _10243__910 (.L_HI(net910));
 sg13g2_tiehi _10242__911 (.L_HI(net911));
 sg13g2_tiehi _10241__912 (.L_HI(net912));
 sg13g2_tiehi _10240__913 (.L_HI(net913));
 sg13g2_tiehi _10239__914 (.L_HI(net914));
 sg13g2_tiehi _10238__915 (.L_HI(net915));
 sg13g2_tiehi _10237__916 (.L_HI(net916));
 sg13g2_tiehi _10236__917 (.L_HI(net917));
 sg13g2_tiehi _10235__918 (.L_HI(net918));
 sg13g2_tiehi _10234__919 (.L_HI(net919));
 sg13g2_tiehi _10233__920 (.L_HI(net920));
 sg13g2_tiehi _10232__921 (.L_HI(net921));
 sg13g2_tiehi _10231__922 (.L_HI(net922));
 sg13g2_tiehi _10230__923 (.L_HI(net923));
 sg13g2_tiehi _10229__924 (.L_HI(net924));
 sg13g2_tiehi _10228__925 (.L_HI(net925));
 sg13g2_tiehi _10227__926 (.L_HI(net926));
 sg13g2_tiehi _10226__927 (.L_HI(net927));
 sg13g2_tiehi _10225__928 (.L_HI(net928));
 sg13g2_tiehi _10224__929 (.L_HI(net929));
 sg13g2_tiehi _10223__930 (.L_HI(net930));
 sg13g2_tiehi _10222__931 (.L_HI(net931));
 sg13g2_tiehi _10221__932 (.L_HI(net932));
 sg13g2_tiehi _10220__933 (.L_HI(net933));
 sg13g2_tiehi _10219__934 (.L_HI(net934));
 sg13g2_tiehi _10218__935 (.L_HI(net935));
 sg13g2_tiehi _10217__936 (.L_HI(net936));
 sg13g2_tiehi _10216__937 (.L_HI(net937));
 sg13g2_tiehi _10215__938 (.L_HI(net938));
 sg13g2_tiehi _10214__939 (.L_HI(net939));
 sg13g2_tiehi _10213__940 (.L_HI(net940));
 sg13g2_tiehi _10212__941 (.L_HI(net941));
 sg13g2_tiehi _10211__942 (.L_HI(net942));
 sg13g2_tiehi _10210__943 (.L_HI(net943));
 sg13g2_tiehi _10209__944 (.L_HI(net944));
 sg13g2_tiehi _10208__945 (.L_HI(net945));
 sg13g2_tiehi _10207__946 (.L_HI(net946));
 sg13g2_tiehi _10206__947 (.L_HI(net947));
 sg13g2_tiehi _10205__948 (.L_HI(net948));
 sg13g2_tiehi _10204__949 (.L_HI(net949));
 sg13g2_tiehi _10203__950 (.L_HI(net950));
 sg13g2_tiehi _10202__951 (.L_HI(net951));
 sg13g2_tiehi _10201__952 (.L_HI(net952));
 sg13g2_tiehi _10200__953 (.L_HI(net953));
 sg13g2_tiehi _10199__954 (.L_HI(net954));
 sg13g2_tiehi _10198__955 (.L_HI(net955));
 sg13g2_tiehi _10197__956 (.L_HI(net956));
 sg13g2_tiehi _10196__957 (.L_HI(net957));
 sg13g2_tiehi _10195__958 (.L_HI(net958));
 sg13g2_tiehi _10194__959 (.L_HI(net959));
 sg13g2_tiehi _10193__960 (.L_HI(net960));
 sg13g2_tiehi _10192__961 (.L_HI(net961));
 sg13g2_tiehi _10191__962 (.L_HI(net962));
 sg13g2_tiehi _10190__963 (.L_HI(net963));
 sg13g2_tiehi _10189__964 (.L_HI(net964));
 sg13g2_tiehi _10188__965 (.L_HI(net965));
 sg13g2_tiehi _10187__966 (.L_HI(net966));
 sg13g2_tiehi _10186__967 (.L_HI(net967));
 sg13g2_tiehi _10185__968 (.L_HI(net968));
 sg13g2_tiehi _10184__969 (.L_HI(net969));
 sg13g2_tiehi _10183__970 (.L_HI(net970));
 sg13g2_tiehi _10182__971 (.L_HI(net971));
 sg13g2_tiehi _10181__972 (.L_HI(net972));
 sg13g2_tiehi _10180__973 (.L_HI(net973));
 sg13g2_tiehi _10179__974 (.L_HI(net974));
 sg13g2_tiehi _10178__975 (.L_HI(net975));
 sg13g2_tiehi _10177__976 (.L_HI(net976));
 sg13g2_tiehi _10176__977 (.L_HI(net977));
 sg13g2_tiehi _10175__978 (.L_HI(net978));
 sg13g2_tiehi _10174__979 (.L_HI(net979));
 sg13g2_tiehi _10173__980 (.L_HI(net980));
 sg13g2_tiehi _10172__981 (.L_HI(net981));
 sg13g2_tiehi _10171__982 (.L_HI(net982));
 sg13g2_tiehi _10170__983 (.L_HI(net983));
 sg13g2_tiehi _10169__984 (.L_HI(net984));
 sg13g2_tiehi _10168__985 (.L_HI(net985));
 sg13g2_tiehi _10167__986 (.L_HI(net986));
 sg13g2_tiehi _10166__987 (.L_HI(net987));
 sg13g2_tiehi _10165__988 (.L_HI(net988));
 sg13g2_tiehi _10164__989 (.L_HI(net989));
 sg13g2_tiehi _10163__990 (.L_HI(net990));
 sg13g2_tiehi _10162__991 (.L_HI(net991));
 sg13g2_tiehi _10161__992 (.L_HI(net992));
 sg13g2_tiehi _10160__993 (.L_HI(net993));
 sg13g2_tiehi _10159__994 (.L_HI(net994));
 sg13g2_tiehi _10158__995 (.L_HI(net995));
 sg13g2_tiehi _10157__996 (.L_HI(net996));
 sg13g2_tiehi _10156__997 (.L_HI(net997));
 sg13g2_tiehi _10155__998 (.L_HI(net998));
 sg13g2_tiehi _10154__999 (.L_HI(net999));
 sg13g2_tiehi _10153__1000 (.L_HI(net1000));
 sg13g2_tiehi _10152__1001 (.L_HI(net1001));
 sg13g2_tiehi _10151__1002 (.L_HI(net1002));
 sg13g2_tiehi _10150__1003 (.L_HI(net1003));
 sg13g2_tiehi _10149__1004 (.L_HI(net1004));
 sg13g2_tiehi _10148__1005 (.L_HI(net1005));
 sg13g2_tiehi _10147__1006 (.L_HI(net1006));
 sg13g2_tiehi _10146__1007 (.L_HI(net1007));
 sg13g2_tiehi _10145__1008 (.L_HI(net1008));
 sg13g2_tiehi _10144__1009 (.L_HI(net1009));
 sg13g2_tiehi _10143__1010 (.L_HI(net1010));
 sg13g2_tiehi _10142__1011 (.L_HI(net1011));
 sg13g2_tiehi _10141__1012 (.L_HI(net1012));
 sg13g2_tiehi _10140__1013 (.L_HI(net1013));
 sg13g2_tiehi _10139__1014 (.L_HI(net1014));
 sg13g2_tiehi _10138__1015 (.L_HI(net1015));
 sg13g2_tiehi _10137__1016 (.L_HI(net1016));
 sg13g2_tiehi _10136__1017 (.L_HI(net1017));
 sg13g2_tiehi _10135__1018 (.L_HI(net1018));
 sg13g2_tiehi _10134__1019 (.L_HI(net1019));
 sg13g2_tiehi _10133__1020 (.L_HI(net1020));
 sg13g2_tiehi _10132__1021 (.L_HI(net1021));
 sg13g2_tiehi _10131__1022 (.L_HI(net1022));
 sg13g2_tiehi _10130__1023 (.L_HI(net1023));
 sg13g2_tiehi _10129__1024 (.L_HI(net1024));
 sg13g2_tiehi _10128__1025 (.L_HI(net1025));
 sg13g2_tiehi _10127__1026 (.L_HI(net1026));
 sg13g2_tiehi _10126__1027 (.L_HI(net1027));
 sg13g2_tiehi _10125__1028 (.L_HI(net1028));
 sg13g2_tiehi _10124__1029 (.L_HI(net1029));
 sg13g2_tiehi _10123__1030 (.L_HI(net1030));
 sg13g2_tiehi _10122__1031 (.L_HI(net1031));
 sg13g2_tiehi _10121__1032 (.L_HI(net1032));
 sg13g2_tiehi _10120__1033 (.L_HI(net1033));
 sg13g2_tiehi _10119__1034 (.L_HI(net1034));
 sg13g2_tiehi _10118__1035 (.L_HI(net1035));
 sg13g2_tiehi _10117__1036 (.L_HI(net1036));
 sg13g2_tiehi _10116__1037 (.L_HI(net1037));
 sg13g2_tiehi _10115__1038 (.L_HI(net1038));
 sg13g2_tiehi _10114__1039 (.L_HI(net1039));
 sg13g2_tiehi _10113__1040 (.L_HI(net1040));
 sg13g2_tiehi _10112__1041 (.L_HI(net1041));
 sg13g2_tiehi _10111__1042 (.L_HI(net1042));
 sg13g2_tiehi _10110__1043 (.L_HI(net1043));
 sg13g2_tiehi _10109__1044 (.L_HI(net1044));
 sg13g2_tiehi _10108__1045 (.L_HI(net1045));
 sg13g2_tiehi _10107__1046 (.L_HI(net1046));
 sg13g2_tiehi _10106__1047 (.L_HI(net1047));
 sg13g2_tiehi _10105__1048 (.L_HI(net1048));
 sg13g2_tiehi _10104__1049 (.L_HI(net1049));
 sg13g2_tiehi _10103__1050 (.L_HI(net1050));
 sg13g2_tiehi _10102__1051 (.L_HI(net1051));
 sg13g2_tiehi _10101__1052 (.L_HI(net1052));
 sg13g2_tiehi _10100__1053 (.L_HI(net1053));
 sg13g2_tiehi _10099__1054 (.L_HI(net1054));
 sg13g2_tiehi _10098__1055 (.L_HI(net1055));
 sg13g2_tiehi _10097__1056 (.L_HI(net1056));
 sg13g2_tiehi _10096__1057 (.L_HI(net1057));
 sg13g2_tiehi _10095__1058 (.L_HI(net1058));
 sg13g2_tiehi _10094__1059 (.L_HI(net1059));
 sg13g2_tiehi _10093__1060 (.L_HI(net1060));
 sg13g2_tiehi _10092__1061 (.L_HI(net1061));
 sg13g2_tiehi _10091__1062 (.L_HI(net1062));
 sg13g2_tiehi _10090__1063 (.L_HI(net1063));
 sg13g2_tiehi _10089__1064 (.L_HI(net1064));
 sg13g2_tiehi _10088__1065 (.L_HI(net1065));
 sg13g2_tiehi _10087__1066 (.L_HI(net1066));
 sg13g2_tiehi _10086__1067 (.L_HI(net1067));
 sg13g2_tiehi _10085__1068 (.L_HI(net1068));
 sg13g2_tiehi _10084__1069 (.L_HI(net1069));
 sg13g2_tiehi _10083__1070 (.L_HI(net1070));
 sg13g2_tiehi _10082__1071 (.L_HI(net1071));
 sg13g2_tiehi _10081__1072 (.L_HI(net1072));
 sg13g2_tiehi _10080__1073 (.L_HI(net1073));
 sg13g2_tiehi _10079__1074 (.L_HI(net1074));
 sg13g2_tiehi _10078__1075 (.L_HI(net1075));
 sg13g2_tiehi _10077__1076 (.L_HI(net1076));
 sg13g2_tiehi _10076__1077 (.L_HI(net1077));
 sg13g2_tiehi _10075__1078 (.L_HI(net1078));
 sg13g2_tiehi _10074__1079 (.L_HI(net1079));
 sg13g2_tiehi _10073__1080 (.L_HI(net1080));
 sg13g2_tiehi _10072__1081 (.L_HI(net1081));
 sg13g2_tiehi _10071__1082 (.L_HI(net1082));
 sg13g2_tiehi _10070__1083 (.L_HI(net1083));
 sg13g2_tiehi _10069__1084 (.L_HI(net1084));
 sg13g2_tiehi _10068__1085 (.L_HI(net1085));
 sg13g2_tiehi _10067__1086 (.L_HI(net1086));
 sg13g2_tiehi _10066__1087 (.L_HI(net1087));
 sg13g2_tiehi _10065__1088 (.L_HI(net1088));
 sg13g2_tiehi _10293__1089 (.L_HI(net1089));
 sg13g2_tiehi _10294__1090 (.L_HI(net1090));
 sg13g2_tiehi _10295__1091 (.L_HI(net1091));
 sg13g2_tiehi _10296__1092 (.L_HI(net1092));
 sg13g2_tiehi _10297__1093 (.L_HI(net1093));
 sg13g2_tiehi _10298__1094 (.L_HI(net1094));
 sg13g2_tiehi _10299__1095 (.L_HI(net1095));
 sg13g2_tiehi _10300__1096 (.L_HI(net1096));
 sg13g2_tiehi _10301__1097 (.L_HI(net1097));
 sg13g2_tiehi _10302__1098 (.L_HI(net1098));
 sg13g2_tiehi _10303__1099 (.L_HI(net1099));
 sg13g2_tiehi _10304__1100 (.L_HI(net1100));
 sg13g2_tiehi _10305__1101 (.L_HI(net1101));
 sg13g2_tiehi _10306__1102 (.L_HI(net1102));
 sg13g2_tiehi _10307__1103 (.L_HI(net1103));
 sg13g2_tiehi _10308__1104 (.L_HI(net1104));
 sg13g2_tiehi _10309__1105 (.L_HI(net1105));
 sg13g2_tiehi _10310__1106 (.L_HI(net1106));
 sg13g2_tiehi _10311__1107 (.L_HI(net1107));
 sg13g2_tiehi _10312__1108 (.L_HI(net1108));
 sg13g2_tiehi _10313__1109 (.L_HI(net1109));
 sg13g2_tiehi _10314__1110 (.L_HI(net1110));
 sg13g2_tiehi _10315__1111 (.L_HI(net1111));
 sg13g2_tiehi _10316__1112 (.L_HI(net1112));
 sg13g2_tiehi _10317__1113 (.L_HI(net1113));
 sg13g2_tiehi _10318__1114 (.L_HI(net1114));
 sg13g2_tiehi _10319__1115 (.L_HI(net1115));
 sg13g2_tiehi _10320__1116 (.L_HI(net1116));
 sg13g2_tiehi _10321__1117 (.L_HI(net1117));
 sg13g2_tiehi _10322__1118 (.L_HI(net1118));
 sg13g2_tiehi _10323__1119 (.L_HI(net1119));
 sg13g2_tiehi _10324__1120 (.L_HI(net1120));
 sg13g2_tiehi _10325__1121 (.L_HI(net1121));
 sg13g2_tiehi _10326__1122 (.L_HI(net1122));
 sg13g2_tiehi _10327__1123 (.L_HI(net1123));
 sg13g2_tiehi _10328__1124 (.L_HI(net1124));
 sg13g2_tiehi _10329__1125 (.L_HI(net1125));
 sg13g2_tiehi _10330__1126 (.L_HI(net1126));
 sg13g2_tiehi _10331__1127 (.L_HI(net1127));
 sg13g2_tiehi _10332__1128 (.L_HI(net1128));
 sg13g2_tiehi _10333__1129 (.L_HI(net1129));
 sg13g2_tiehi _10334__1130 (.L_HI(net1130));
 sg13g2_tiehi _10335__1131 (.L_HI(net1131));
 sg13g2_tiehi _10336__1132 (.L_HI(net1132));
 sg13g2_tiehi _10337__1133 (.L_HI(net1133));
 sg13g2_tiehi _10338__1134 (.L_HI(net1134));
 sg13g2_tiehi _10339__1135 (.L_HI(net1135));
 sg13g2_tiehi _10340__1136 (.L_HI(net1136));
 sg13g2_tiehi _10341__1137 (.L_HI(net1137));
 sg13g2_tiehi _10342__1138 (.L_HI(net1138));
 sg13g2_tiehi _10343__1139 (.L_HI(net1139));
 sg13g2_tiehi _10344__1140 (.L_HI(net1140));
 sg13g2_tiehi _10345__1141 (.L_HI(net1141));
 sg13g2_tiehi _10346__1142 (.L_HI(net1142));
 sg13g2_tiehi _10347__1143 (.L_HI(net1143));
 sg13g2_tiehi _10348__1144 (.L_HI(net1144));
 sg13g2_tiehi _10349__1145 (.L_HI(net1145));
 sg13g2_tiehi _10350__1146 (.L_HI(net1146));
 sg13g2_tiehi _10351__1147 (.L_HI(net1147));
 sg13g2_tiehi _10352__1148 (.L_HI(net1148));
 sg13g2_tiehi _10064__1149 (.L_HI(net1149));
 sg13g2_tiehi _10063__1150 (.L_HI(net1150));
 sg13g2_tiehi _10062__1151 (.L_HI(net1151));
 sg13g2_tiehi _10061__1152 (.L_HI(net1152));
 sg13g2_tiehi _10060__1153 (.L_HI(net1153));
 sg13g2_tiehi _10059__1154 (.L_HI(net1154));
 sg13g2_tiehi _10058__1155 (.L_HI(net1155));
 sg13g2_tiehi _10057__1156 (.L_HI(net1156));
 sg13g2_tiehi _10056__1157 (.L_HI(net1157));
 sg13g2_tiehi _10055__1158 (.L_HI(net1158));
 sg13g2_tiehi _10054__1159 (.L_HI(net1159));
 sg13g2_tiehi _10053__1160 (.L_HI(net1160));
 sg13g2_tiehi _10052__1161 (.L_HI(net1161));
 sg13g2_tiehi _10051__1162 (.L_HI(net1162));
 sg13g2_tiehi _10050__1163 (.L_HI(net1163));
 sg13g2_tiehi _10049__1164 (.L_HI(net1164));
 sg13g2_tiehi _10048__1165 (.L_HI(net1165));
 sg13g2_tiehi _10047__1166 (.L_HI(net1166));
 sg13g2_tiehi _10046__1167 (.L_HI(net1167));
 sg13g2_tiehi _10045__1168 (.L_HI(net1168));
 sg13g2_tiehi _10044__1169 (.L_HI(net1169));
 sg13g2_tiehi _10043__1170 (.L_HI(net1170));
 sg13g2_tiehi _10042__1171 (.L_HI(net1171));
 sg13g2_tiehi _10041__1172 (.L_HI(net1172));
 sg13g2_tiehi _10040__1173 (.L_HI(net1173));
 sg13g2_tiehi _10039__1174 (.L_HI(net1174));
 sg13g2_tiehi _10038__1175 (.L_HI(net1175));
 sg13g2_tiehi _10037__1176 (.L_HI(net1176));
 sg13g2_tiehi _10036__1177 (.L_HI(net1177));
 sg13g2_tiehi _10035__1178 (.L_HI(net1178));
 sg13g2_tiehi _10034__1179 (.L_HI(net1179));
 sg13g2_tiehi _10033__1180 (.L_HI(net1180));
 sg13g2_tiehi _10032__1181 (.L_HI(net1181));
 sg13g2_tiehi _10353__1182 (.L_HI(net1182));
 sg13g2_tiehi _10031__1183 (.L_HI(net1183));
 sg13g2_tiehi _10030__1184 (.L_HI(net1184));
 sg13g2_tiehi _10029__1185 (.L_HI(net1185));
 sg13g2_tiehi _10387__1186 (.L_HI(net1186));
 sg13g2_tiehi _10028__1187 (.L_HI(net1187));
 sg13g2_tiehi _10027__1188 (.L_HI(net1188));
 sg13g2_tiehi _10391__1189 (.L_HI(net1189));
 sg13g2_tiehi _10394__1190 (.L_HI(net1190));
 sg13g2_tiehi _10395__1191 (.L_HI(net1191));
 sg13g2_tiehi _10396__1192 (.L_HI(net1192));
 sg13g2_tiehi _10397__1193 (.L_HI(net1193));
 sg13g2_tiehi _10398__1194 (.L_HI(net1194));
 sg13g2_tiehi _10399__1195 (.L_HI(net1195));
 sg13g2_tiehi _10400__1196 (.L_HI(net1196));
 sg13g2_tiehi _10401__1197 (.L_HI(net1197));
 sg13g2_tiehi _10402__1198 (.L_HI(net1198));
 sg13g2_tiehi _10403__1199 (.L_HI(net1199));
 sg13g2_tiehi _10404__1200 (.L_HI(net1200));
 sg13g2_tiehi _10405__1201 (.L_HI(net1201));
 sg13g2_tiehi _10406__1202 (.L_HI(net1202));
 sg13g2_tiehi _10407__1203 (.L_HI(net1203));
 sg13g2_tiehi _10408__1204 (.L_HI(net1204));
 sg13g2_tiehi _10409__1205 (.L_HI(net1205));
 sg13g2_tiehi _10410__1206 (.L_HI(net1206));
 sg13g2_tiehi _10411__1207 (.L_HI(net1207));
 sg13g2_tiehi _10412__1208 (.L_HI(net1208));
 sg13g2_tiehi _10413__1209 (.L_HI(net1209));
 sg13g2_tiehi _10414__1210 (.L_HI(net1210));
 sg13g2_tiehi _10415__1211 (.L_HI(net1211));
 sg13g2_tiehi _10416__1212 (.L_HI(net1212));
 sg13g2_tiehi _10417__1213 (.L_HI(net1213));
 sg13g2_tiehi _10418__1214 (.L_HI(net1214));
 sg13g2_tiehi _10419__1215 (.L_HI(net1215));
 sg13g2_tiehi _10420__1216 (.L_HI(net1216));
 sg13g2_tiehi _10421__1217 (.L_HI(net1217));
 sg13g2_tiehi _10422__1218 (.L_HI(net1218));
 sg13g2_tiehi _10423__1219 (.L_HI(net1219));
 sg13g2_tiehi _10424__1220 (.L_HI(net1220));
 sg13g2_tiehi _10026__1221 (.L_HI(net1221));
 sg13g2_tiehi _10025__1222 (.L_HI(net1222));
 sg13g2_tiehi _10024__1223 (.L_HI(net1223));
 sg13g2_tiehi _10023__1224 (.L_HI(net1224));
 sg13g2_tiehi _10022__1225 (.L_HI(net1225));
 sg13g2_tiehi _10021__1226 (.L_HI(net1226));
 sg13g2_tiehi _10020__1227 (.L_HI(net1227));
 sg13g2_tiehi _10019__1228 (.L_HI(net1228));
 sg13g2_tiehi _10018__1229 (.L_HI(net1229));
 sg13g2_tiehi _10017__1230 (.L_HI(net1230));
 sg13g2_tiehi _10016__1231 (.L_HI(net1231));
 sg13g2_tiehi _10015__1232 (.L_HI(net1232));
 sg13g2_tiehi _10014__1233 (.L_HI(net1233));
 sg13g2_tiehi _10013__1234 (.L_HI(net1234));
 sg13g2_tiehi _10012__1235 (.L_HI(net1235));
 sg13g2_tiehi _10011__1236 (.L_HI(net1236));
 sg13g2_tiehi _10010__1237 (.L_HI(net1237));
 sg13g2_tiehi _10009__1238 (.L_HI(net1238));
 sg13g2_tiehi _10008__1239 (.L_HI(net1239));
 sg13g2_tiehi _10007__1240 (.L_HI(net1240));
 sg13g2_tiehi _10006__1241 (.L_HI(net1241));
 sg13g2_tiehi _10005__1242 (.L_HI(net1242));
 sg13g2_tiehi _10004__1243 (.L_HI(net1243));
 sg13g2_tiehi _10003__1244 (.L_HI(net1244));
 sg13g2_tiehi _10002__1245 (.L_HI(net1245));
 sg13g2_tiehi _10001__1246 (.L_HI(net1246));
 sg13g2_tiehi _10000__1247 (.L_HI(net1247));
 sg13g2_tiehi _09999__1248 (.L_HI(net1248));
 sg13g2_tiehi _09998__1249 (.L_HI(net1249));
 sg13g2_tiehi _09997__1250 (.L_HI(net1250));
 sg13g2_tiehi _09996__1251 (.L_HI(net1251));
 sg13g2_tiehi _09995__1252 (.L_HI(net1252));
 sg13g2_tiehi _09994__1253 (.L_HI(net1253));
 sg13g2_tiehi _09993__1254 (.L_HI(net1254));
 sg13g2_tiehi _09992__1255 (.L_HI(net1255));
 sg13g2_tiehi _09991__1256 (.L_HI(net1256));
 sg13g2_tiehi _09990__1257 (.L_HI(net1257));
 sg13g2_tiehi _09989__1258 (.L_HI(net1258));
 sg13g2_tiehi _09988__1259 (.L_HI(net1259));
 sg13g2_tiehi _09987__1260 (.L_HI(net1260));
 sg13g2_tiehi _09986__1261 (.L_HI(net1261));
 sg13g2_tiehi _09985__1262 (.L_HI(net1262));
 sg13g2_tiehi _09984__1263 (.L_HI(net1263));
 sg13g2_tiehi _09983__1264 (.L_HI(net1264));
 sg13g2_tiehi _09982__1265 (.L_HI(net1265));
 sg13g2_tiehi _09981__1266 (.L_HI(net1266));
 sg13g2_tiehi _09980__1267 (.L_HI(net1267));
 sg13g2_tiehi _09979__1268 (.L_HI(net1268));
 sg13g2_tiehi _09978__1269 (.L_HI(net1269));
 sg13g2_tiehi _09977__1270 (.L_HI(net1270));
 sg13g2_tiehi _09976__1271 (.L_HI(net1271));
 sg13g2_tiehi _09975__1272 (.L_HI(net1272));
 sg13g2_tiehi _09974__1273 (.L_HI(net1273));
 sg13g2_tiehi _09973__1274 (.L_HI(net1274));
 sg13g2_tiehi _09972__1275 (.L_HI(net1275));
 sg13g2_tiehi _09971__1276 (.L_HI(net1276));
 sg13g2_tiehi _09970__1277 (.L_HI(net1277));
 sg13g2_tiehi _09969__1278 (.L_HI(net1278));
 sg13g2_tiehi _09968__1279 (.L_HI(net1279));
 sg13g2_tiehi _09967__1280 (.L_HI(net1280));
 sg13g2_tiehi _09966__1281 (.L_HI(net1281));
 sg13g2_tiehi _09965__1282 (.L_HI(net1282));
 sg13g2_tiehi _09964__1283 (.L_HI(net1283));
 sg13g2_tiehi _09963__1284 (.L_HI(net1284));
 sg13g2_tiehi _09962__1285 (.L_HI(net1285));
 sg13g2_tiehi _09961__1286 (.L_HI(net1286));
 sg13g2_tiehi _09960__1287 (.L_HI(net1287));
 sg13g2_tiehi _09959__1288 (.L_HI(net1288));
 sg13g2_tiehi _09958__1289 (.L_HI(net1289));
 sg13g2_tiehi _10425__1290 (.L_HI(net1290));
 sg13g2_tiehi _09957__1291 (.L_HI(net1291));
 sg13g2_tiehi _09956__1292 (.L_HI(net1292));
 sg13g2_tiehi _09955__1293 (.L_HI(net1293));
 sg13g2_tiehi _09954__1294 (.L_HI(net1294));
 sg13g2_tiehi _09953__1295 (.L_HI(net1295));
 sg13g2_tiehi _09952__1296 (.L_HI(net1296));
 sg13g2_tiehi _09951__1297 (.L_HI(net1297));
 sg13g2_tiehi _09950__1298 (.L_HI(net1298));
 sg13g2_tiehi _09949__1299 (.L_HI(net1299));
 sg13g2_tiehi _09948__1300 (.L_HI(net1300));
 sg13g2_tiehi _09947__1301 (.L_HI(net1301));
 sg13g2_tiehi _09946__1302 (.L_HI(net1302));
 sg13g2_tiehi _09945__1303 (.L_HI(net1303));
 sg13g2_tiehi _09944__1304 (.L_HI(net1304));
 sg13g2_tiehi _09943__1305 (.L_HI(net1305));
 sg13g2_tiehi _09942__1306 (.L_HI(net1306));
 sg13g2_tiehi _09941__1307 (.L_HI(net1307));
 sg13g2_tiehi _09940__1308 (.L_HI(net1308));
 sg13g2_tiehi _09939__1309 (.L_HI(net1309));
 sg13g2_tiehi _09938__1310 (.L_HI(net1310));
 sg13g2_tiehi _09937__1311 (.L_HI(net1311));
 sg13g2_tiehi _09936__1312 (.L_HI(net1312));
 sg13g2_tiehi _09935__1313 (.L_HI(net1313));
 sg13g2_tiehi _09934__1314 (.L_HI(net1314));
 sg13g2_tiehi _09933__1315 (.L_HI(net1315));
 sg13g2_tiehi _09932__1316 (.L_HI(net1316));
 sg13g2_tiehi _09931__1317 (.L_HI(net1317));
 sg13g2_tiehi _09930__1318 (.L_HI(net1318));
 sg13g2_tiehi _09929__1319 (.L_HI(net1319));
 sg13g2_tiehi _09928__1320 (.L_HI(net1320));
 sg13g2_tiehi _09927__1321 (.L_HI(net1321));
 sg13g2_tiehi _09926__1322 (.L_HI(net1322));
 sg13g2_tiehi _09925__1323 (.L_HI(net1323));
 sg13g2_tiehi _09924__1324 (.L_HI(net1324));
 sg13g2_tiehi _09923__1325 (.L_HI(net1325));
 sg13g2_tiehi _09922__1326 (.L_HI(net1326));
 sg13g2_tiehi _09921__1327 (.L_HI(net1327));
 sg13g2_tiehi _09920__1328 (.L_HI(net1328));
 sg13g2_tiehi _09919__1329 (.L_HI(net1329));
 sg13g2_tiehi _09918__1330 (.L_HI(net1330));
 sg13g2_tiehi _09917__1331 (.L_HI(net1331));
 sg13g2_tiehi _09916__1332 (.L_HI(net1332));
 sg13g2_tiehi _10495__1333 (.L_HI(net1333));
 sg13g2_tiehi _10538__1334 (.L_HI(net1334));
 sg13g2_tiehi _09915__1335 (.L_HI(net1335));
 sg13g2_tiehi _09914__1336 (.L_HI(net1336));
 sg13g2_tiehi _09913__1337 (.L_HI(net1337));
 sg13g2_tiehi _09912__1338 (.L_HI(net1338));
 sg13g2_tiehi _09911__1339 (.L_HI(net1339));
 sg13g2_tiehi _09910__1340 (.L_HI(net1340));
 sg13g2_tiehi _09909__1341 (.L_HI(net1341));
 sg13g2_tiehi _09908__1342 (.L_HI(net1342));
 sg13g2_tiehi _09907__1343 (.L_HI(net1343));
 sg13g2_tiehi _09906__1344 (.L_HI(net1344));
 sg13g2_tiehi _09905__1345 (.L_HI(net1345));
 sg13g2_tiehi _09904__1346 (.L_HI(net1346));
 sg13g2_tiehi _09903__1347 (.L_HI(net1347));
 sg13g2_tiehi _09902__1348 (.L_HI(net1348));
 sg13g2_tiehi _09901__1349 (.L_HI(net1349));
 sg13g2_tiehi _09900__1350 (.L_HI(net1350));
 sg13g2_tiehi _09899__1351 (.L_HI(net1351));
 sg13g2_tiehi _09898__1352 (.L_HI(net1352));
 sg13g2_tiehi _09897__1353 (.L_HI(net1353));
 sg13g2_tiehi _09896__1354 (.L_HI(net1354));
 sg13g2_tiehi _09895__1355 (.L_HI(net1355));
 sg13g2_tiehi _09894__1356 (.L_HI(net1356));
 sg13g2_tiehi _09893__1357 (.L_HI(net1357));
 sg13g2_tiehi _09892__1358 (.L_HI(net1358));
 sg13g2_tiehi _09891__1359 (.L_HI(net1359));
 sg13g2_tiehi _09890__1360 (.L_HI(net1360));
 sg13g2_tiehi _09889__1361 (.L_HI(net1361));
 sg13g2_tiehi _09888__1362 (.L_HI(net1362));
 sg13g2_tiehi _09887__1363 (.L_HI(net1363));
 sg13g2_tiehi _09886__1364 (.L_HI(net1364));
 sg13g2_tiehi _09885__1365 (.L_HI(net1365));
 sg13g2_tiehi _09884__1366 (.L_HI(net1366));
 sg13g2_tiehi _10539__1367 (.L_HI(net1367));
 sg13g2_tiehi _09883__1368 (.L_HI(net1368));
 sg13g2_tiehi _09882__1369 (.L_HI(net1369));
 sg13g2_tiehi _09881__1370 (.L_HI(net1370));
 sg13g2_tiehi _09880__1371 (.L_HI(net1371));
 sg13g2_tiehi _09879__1372 (.L_HI(net1372));
 sg13g2_tiehi _09878__1373 (.L_HI(net1373));
 sg13g2_tiehi tt_um_ECM24_serv_soc_top_1374 (.L_HI(net1374));
 sg13g2_tiehi tt_um_ECM24_serv_soc_top_1375 (.L_HI(net1375));
 sg13g2_tiehi tt_um_ECM24_serv_soc_top_1376 (.L_HI(net1376));
 sg13g2_tiehi tt_um_ECM24_serv_soc_top_1377 (.L_HI(net1377));
 sg13g2_tiehi tt_um_ECM24_serv_soc_top_1378 (.L_HI(net1378));
 sg13g2_tiehi tt_um_ECM24_serv_soc_top_1379 (.L_HI(net1379));
 sg13g2_inv_1 _05321__1 (.Y(net1380),
    .A(clknet_1_1__leaf_clk));
 sg13g2_tielo tt_um_ECM24_serv_soc_top_8 (.L_LO(net8));
 sg13g2_tielo tt_um_ECM24_serv_soc_top_9 (.L_LO(net9));
 sg13g2_tielo tt_um_ECM24_serv_soc_top_10 (.L_LO(net10));
 sg13g2_tielo tt_um_ECM24_serv_soc_top_11 (.L_LO(net11));
 sg13g2_tielo tt_um_ECM24_serv_soc_top_12 (.L_LO(net12));
 sg13g2_tielo tt_um_ECM24_serv_soc_top_13 (.L_LO(net13));
 sg13g2_tielo tt_um_ECM24_serv_soc_top_14 (.L_LO(net14));
 sg13g2_tielo tt_um_ECM24_serv_soc_top_15 (.L_LO(net15));
 sg13g2_tielo tt_um_ECM24_serv_soc_top_16 (.L_LO(net16));
 sg13g2_tielo tt_um_ECM24_serv_soc_top_17 (.L_LO(net17));
 sg13g2_tiehi _09877__18 (.L_HI(net18));
 sg13g2_buf_1 _11953_ (.A(\ram_spi_if.spi_cs_n ),
    .X(uio_out[0]));
 sg13g2_buf_1 _11954_ (.A(\ram_spi_if.spi_mosi ),
    .X(uio_out[1]));
 sg13g2_buf_1 _11955_ (.A(\ram_spi_if.spi_clk ),
    .X(uio_out[3]));
 sg13g2_buf_8 fanout1749 (.A(net1753),
    .X(net1749));
 sg13g2_buf_8 fanout1750 (.A(net1753),
    .X(net1750));
 sg13g2_buf_8 fanout1751 (.A(net1753),
    .X(net1751));
 sg13g2_buf_8 fanout1752 (.A(net1753),
    .X(net1752));
 sg13g2_buf_8 fanout1753 (.A(net1759),
    .X(net1753));
 sg13g2_buf_8 fanout1754 (.A(net1759),
    .X(net1754));
 sg13g2_buf_8 fanout1755 (.A(net1759),
    .X(net1755));
 sg13g2_buf_8 fanout1756 (.A(net1757),
    .X(net1756));
 sg13g2_buf_8 fanout1757 (.A(net1758),
    .X(net1757));
 sg13g2_buf_8 fanout1758 (.A(net1759),
    .X(net1758));
 sg13g2_buf_8 fanout1759 (.A(_03851_),
    .X(net1759));
 sg13g2_buf_8 fanout1760 (.A(net1761),
    .X(net1760));
 sg13g2_buf_8 fanout1761 (.A(net1764),
    .X(net1761));
 sg13g2_buf_8 fanout1762 (.A(net1763),
    .X(net1762));
 sg13g2_buf_8 fanout1763 (.A(net1764),
    .X(net1763));
 sg13g2_buf_8 fanout1764 (.A(_02769_),
    .X(net1764));
 sg13g2_buf_8 fanout1765 (.A(net1769),
    .X(net1765));
 sg13g2_buf_8 fanout1766 (.A(net1769),
    .X(net1766));
 sg13g2_buf_8 fanout1767 (.A(net1768),
    .X(net1767));
 sg13g2_buf_8 fanout1768 (.A(net1769),
    .X(net1768));
 sg13g2_buf_8 fanout1769 (.A(_02769_),
    .X(net1769));
 sg13g2_buf_8 fanout1770 (.A(net1771),
    .X(net1770));
 sg13g2_buf_8 fanout1771 (.A(net1774),
    .X(net1771));
 sg13g2_buf_8 fanout1772 (.A(net1773),
    .X(net1772));
 sg13g2_buf_8 fanout1773 (.A(net1774),
    .X(net1773));
 sg13g2_buf_8 fanout1774 (.A(_02736_),
    .X(net1774));
 sg13g2_buf_8 fanout1775 (.A(net1779),
    .X(net1775));
 sg13g2_buf_8 fanout1776 (.A(net1779),
    .X(net1776));
 sg13g2_buf_8 fanout1777 (.A(net1778),
    .X(net1777));
 sg13g2_buf_8 fanout1778 (.A(net1779),
    .X(net1778));
 sg13g2_buf_8 fanout1779 (.A(_02736_),
    .X(net1779));
 sg13g2_buf_8 fanout1780 (.A(net1790),
    .X(net1780));
 sg13g2_buf_8 fanout1781 (.A(net1790),
    .X(net1781));
 sg13g2_buf_8 fanout1782 (.A(net1783),
    .X(net1782));
 sg13g2_buf_8 fanout1783 (.A(net1790),
    .X(net1783));
 sg13g2_buf_8 fanout1784 (.A(net1789),
    .X(net1784));
 sg13g2_buf_1 fanout1785 (.A(net1789),
    .X(net1785));
 sg13g2_buf_8 fanout1786 (.A(net1789),
    .X(net1786));
 sg13g2_buf_8 fanout1787 (.A(net1789),
    .X(net1787));
 sg13g2_buf_8 fanout1788 (.A(net1789),
    .X(net1788));
 sg13g2_buf_8 fanout1789 (.A(net1790),
    .X(net1789));
 sg13g2_buf_8 fanout1790 (.A(_02642_),
    .X(net1790));
 sg13g2_buf_8 fanout1791 (.A(net1800),
    .X(net1791));
 sg13g2_buf_8 fanout1792 (.A(net1800),
    .X(net1792));
 sg13g2_buf_8 fanout1793 (.A(net1794),
    .X(net1793));
 sg13g2_buf_8 fanout1794 (.A(net1800),
    .X(net1794));
 sg13g2_buf_8 fanout1795 (.A(net1797),
    .X(net1795));
 sg13g2_buf_1 fanout1796 (.A(net1797),
    .X(net1796));
 sg13g2_buf_8 fanout1797 (.A(net1800),
    .X(net1797));
 sg13g2_buf_8 fanout1798 (.A(net1799),
    .X(net1798));
 sg13g2_buf_8 fanout1799 (.A(net1800),
    .X(net1799));
 sg13g2_buf_8 fanout1800 (.A(_02609_),
    .X(net1800));
 sg13g2_buf_8 fanout1801 (.A(net1810),
    .X(net1801));
 sg13g2_buf_8 fanout1802 (.A(net1810),
    .X(net1802));
 sg13g2_buf_8 fanout1803 (.A(net1804),
    .X(net1803));
 sg13g2_buf_8 fanout1804 (.A(net1810),
    .X(net1804));
 sg13g2_buf_8 fanout1805 (.A(net1807),
    .X(net1805));
 sg13g2_buf_1 fanout1806 (.A(net1807),
    .X(net1806));
 sg13g2_buf_8 fanout1807 (.A(net1810),
    .X(net1807));
 sg13g2_buf_8 fanout1808 (.A(net1810),
    .X(net1808));
 sg13g2_buf_8 fanout1809 (.A(net1810),
    .X(net1809));
 sg13g2_buf_8 fanout1810 (.A(_02576_),
    .X(net1810));
 sg13g2_buf_8 fanout1811 (.A(net1820),
    .X(net1811));
 sg13g2_buf_8 fanout1812 (.A(net1820),
    .X(net1812));
 sg13g2_buf_8 fanout1813 (.A(net1814),
    .X(net1813));
 sg13g2_buf_8 fanout1814 (.A(net1820),
    .X(net1814));
 sg13g2_buf_8 fanout1815 (.A(net1817),
    .X(net1815));
 sg13g2_buf_1 fanout1816 (.A(net1817),
    .X(net1816));
 sg13g2_buf_8 fanout1817 (.A(net1820),
    .X(net1817));
 sg13g2_buf_8 fanout1818 (.A(net1820),
    .X(net1818));
 sg13g2_buf_8 fanout1819 (.A(net1820),
    .X(net1819));
 sg13g2_buf_8 fanout1820 (.A(_02543_),
    .X(net1820));
 sg13g2_buf_8 fanout1821 (.A(net1825),
    .X(net1821));
 sg13g2_buf_8 fanout1822 (.A(net1825),
    .X(net1822));
 sg13g2_buf_8 fanout1823 (.A(net1825),
    .X(net1823));
 sg13g2_buf_2 fanout1824 (.A(net1825),
    .X(net1824));
 sg13g2_buf_8 fanout1825 (.A(_02508_),
    .X(net1825));
 sg13g2_buf_8 fanout1826 (.A(net1828),
    .X(net1826));
 sg13g2_buf_1 fanout1827 (.A(net1828),
    .X(net1827));
 sg13g2_buf_8 fanout1828 (.A(_02508_),
    .X(net1828));
 sg13g2_buf_8 fanout1829 (.A(net1831),
    .X(net1829));
 sg13g2_buf_1 fanout1830 (.A(net1831),
    .X(net1830));
 sg13g2_buf_8 fanout1831 (.A(_02508_),
    .X(net1831));
 sg13g2_buf_8 fanout1832 (.A(net1836),
    .X(net1832));
 sg13g2_buf_8 fanout1833 (.A(net1835),
    .X(net1833));
 sg13g2_buf_8 fanout1834 (.A(net1835),
    .X(net1834));
 sg13g2_buf_8 fanout1835 (.A(net1836),
    .X(net1835));
 sg13g2_buf_8 fanout1836 (.A(net1842),
    .X(net1836));
 sg13g2_buf_8 fanout1837 (.A(net1842),
    .X(net1837));
 sg13g2_buf_8 fanout1838 (.A(net1842),
    .X(net1838));
 sg13g2_buf_8 fanout1839 (.A(net1841),
    .X(net1839));
 sg13g2_buf_1 fanout1840 (.A(net1841),
    .X(net1840));
 sg13g2_buf_8 fanout1841 (.A(net1842),
    .X(net1841));
 sg13g2_buf_8 fanout1842 (.A(_02475_),
    .X(net1842));
 sg13g2_buf_8 fanout1843 (.A(net1847),
    .X(net1843));
 sg13g2_buf_8 fanout1844 (.A(net1846),
    .X(net1844));
 sg13g2_buf_8 fanout1845 (.A(net1846),
    .X(net1845));
 sg13g2_buf_8 fanout1846 (.A(net1847),
    .X(net1846));
 sg13g2_buf_8 fanout1847 (.A(net1853),
    .X(net1847));
 sg13g2_buf_8 fanout1848 (.A(net1853),
    .X(net1848));
 sg13g2_buf_8 fanout1849 (.A(net1853),
    .X(net1849));
 sg13g2_buf_8 fanout1850 (.A(net1852),
    .X(net1850));
 sg13g2_buf_1 fanout1851 (.A(net1852),
    .X(net1851));
 sg13g2_buf_8 fanout1852 (.A(net1853),
    .X(net1852));
 sg13g2_buf_8 fanout1853 (.A(_02442_),
    .X(net1853));
 sg13g2_buf_8 fanout1854 (.A(net1855),
    .X(net1854));
 sg13g2_buf_8 fanout1855 (.A(_02409_),
    .X(net1855));
 sg13g2_buf_8 fanout1856 (.A(net1858),
    .X(net1856));
 sg13g2_buf_1 fanout1857 (.A(net1858),
    .X(net1857));
 sg13g2_buf_8 fanout1858 (.A(_02409_),
    .X(net1858));
 sg13g2_buf_8 fanout1859 (.A(net1863),
    .X(net1859));
 sg13g2_buf_8 fanout1860 (.A(net1863),
    .X(net1860));
 sg13g2_buf_8 fanout1861 (.A(net1862),
    .X(net1861));
 sg13g2_buf_8 fanout1862 (.A(net1863),
    .X(net1862));
 sg13g2_buf_8 fanout1863 (.A(_02409_),
    .X(net1863));
 sg13g2_buf_8 fanout1864 (.A(net1865),
    .X(net1864));
 sg13g2_buf_8 fanout1865 (.A(net1868),
    .X(net1865));
 sg13g2_buf_8 fanout1866 (.A(net1868),
    .X(net1866));
 sg13g2_buf_1 fanout1867 (.A(net1868),
    .X(net1867));
 sg13g2_buf_8 fanout1868 (.A(net1874),
    .X(net1868));
 sg13g2_buf_8 fanout1869 (.A(net1870),
    .X(net1869));
 sg13g2_buf_8 fanout1870 (.A(net1874),
    .X(net1870));
 sg13g2_buf_8 fanout1871 (.A(net1873),
    .X(net1871));
 sg13g2_buf_8 fanout1872 (.A(net1873),
    .X(net1872));
 sg13g2_buf_8 fanout1873 (.A(net1874),
    .X(net1873));
 sg13g2_buf_8 fanout1874 (.A(_02376_),
    .X(net1874));
 sg13g2_buf_8 fanout1875 (.A(net1876),
    .X(net1875));
 sg13g2_buf_8 fanout1876 (.A(_02343_),
    .X(net1876));
 sg13g2_buf_8 fanout1877 (.A(net1879),
    .X(net1877));
 sg13g2_buf_1 fanout1878 (.A(net1879),
    .X(net1878));
 sg13g2_buf_8 fanout1879 (.A(_02343_),
    .X(net1879));
 sg13g2_buf_8 fanout1880 (.A(net1884),
    .X(net1880));
 sg13g2_buf_8 fanout1881 (.A(net1884),
    .X(net1881));
 sg13g2_buf_8 fanout1882 (.A(net1883),
    .X(net1882));
 sg13g2_buf_8 fanout1883 (.A(net1884),
    .X(net1883));
 sg13g2_buf_8 fanout1884 (.A(_02343_),
    .X(net1884));
 sg13g2_buf_8 fanout1885 (.A(net1888),
    .X(net1885));
 sg13g2_buf_8 fanout1886 (.A(net1888),
    .X(net1886));
 sg13g2_buf_8 fanout1887 (.A(net1888),
    .X(net1887));
 sg13g2_buf_8 fanout1888 (.A(_02307_),
    .X(net1888));
 sg13g2_buf_8 fanout1889 (.A(net1891),
    .X(net1889));
 sg13g2_buf_1 fanout1890 (.A(net1891),
    .X(net1890));
 sg13g2_buf_8 fanout1891 (.A(_02307_),
    .X(net1891));
 sg13g2_buf_8 fanout1892 (.A(net1894),
    .X(net1892));
 sg13g2_buf_8 fanout1893 (.A(net1894),
    .X(net1893));
 sg13g2_buf_8 fanout1894 (.A(_02307_),
    .X(net1894));
 sg13g2_buf_8 fanout1895 (.A(net1896),
    .X(net1895));
 sg13g2_buf_8 fanout1896 (.A(net1904),
    .X(net1896));
 sg13g2_buf_8 fanout1897 (.A(net1904),
    .X(net1897));
 sg13g2_buf_2 fanout1898 (.A(net1904),
    .X(net1898));
 sg13g2_buf_8 fanout1899 (.A(net1900),
    .X(net1899));
 sg13g2_buf_8 fanout1900 (.A(net1904),
    .X(net1900));
 sg13g2_buf_8 fanout1901 (.A(net1903),
    .X(net1901));
 sg13g2_buf_8 fanout1902 (.A(net1903),
    .X(net1902));
 sg13g2_buf_8 fanout1903 (.A(net1904),
    .X(net1903));
 sg13g2_buf_8 fanout1904 (.A(_02274_),
    .X(net1904));
 sg13g2_buf_8 fanout1905 (.A(net1906),
    .X(net1905));
 sg13g2_buf_8 fanout1906 (.A(net1909),
    .X(net1906));
 sg13g2_buf_8 fanout1907 (.A(net1909),
    .X(net1907));
 sg13g2_buf_1 fanout1908 (.A(net1909),
    .X(net1908));
 sg13g2_buf_8 fanout1909 (.A(net1915),
    .X(net1909));
 sg13g2_buf_8 fanout1910 (.A(net1912),
    .X(net1910));
 sg13g2_buf_1 fanout1911 (.A(net1912),
    .X(net1911));
 sg13g2_buf_8 fanout1912 (.A(net1915),
    .X(net1912));
 sg13g2_buf_8 fanout1913 (.A(net1914),
    .X(net1913));
 sg13g2_buf_8 fanout1914 (.A(net1915),
    .X(net1914));
 sg13g2_buf_8 fanout1915 (.A(_02241_),
    .X(net1915));
 sg13g2_buf_8 fanout1916 (.A(net1917),
    .X(net1916));
 sg13g2_buf_8 fanout1917 (.A(net1920),
    .X(net1917));
 sg13g2_buf_8 fanout1918 (.A(net1919),
    .X(net1918));
 sg13g2_buf_8 fanout1919 (.A(net1920),
    .X(net1919));
 sg13g2_buf_8 fanout1920 (.A(_02208_),
    .X(net1920));
 sg13g2_buf_8 fanout1921 (.A(net1925),
    .X(net1921));
 sg13g2_buf_8 fanout1922 (.A(net1925),
    .X(net1922));
 sg13g2_buf_8 fanout1923 (.A(net1924),
    .X(net1923));
 sg13g2_buf_8 fanout1924 (.A(net1925),
    .X(net1924));
 sg13g2_buf_8 fanout1925 (.A(_02208_),
    .X(net1925));
 sg13g2_buf_8 fanout1926 (.A(net1928),
    .X(net1926));
 sg13g2_buf_1 fanout1927 (.A(net1928),
    .X(net1927));
 sg13g2_buf_8 fanout1928 (.A(net1931),
    .X(net1928));
 sg13g2_buf_8 fanout1929 (.A(net1931),
    .X(net1929));
 sg13g2_buf_1 fanout1930 (.A(net1931),
    .X(net1930));
 sg13g2_buf_8 fanout1931 (.A(_02175_),
    .X(net1931));
 sg13g2_buf_8 fanout1932 (.A(net1936),
    .X(net1932));
 sg13g2_buf_8 fanout1933 (.A(net1936),
    .X(net1933));
 sg13g2_buf_8 fanout1934 (.A(net1935),
    .X(net1934));
 sg13g2_buf_8 fanout1935 (.A(net1936),
    .X(net1935));
 sg13g2_buf_8 fanout1936 (.A(_02175_),
    .X(net1936));
 sg13g2_buf_8 fanout1937 (.A(net1938),
    .X(net1937));
 sg13g2_buf_8 fanout1938 (.A(net1941),
    .X(net1938));
 sg13g2_buf_8 fanout1939 (.A(net1940),
    .X(net1939));
 sg13g2_buf_8 fanout1940 (.A(net1941),
    .X(net1940));
 sg13g2_buf_8 fanout1941 (.A(_02142_),
    .X(net1941));
 sg13g2_buf_8 fanout1942 (.A(net1946),
    .X(net1942));
 sg13g2_buf_8 fanout1943 (.A(net1946),
    .X(net1943));
 sg13g2_buf_8 fanout1944 (.A(net1945),
    .X(net1944));
 sg13g2_buf_8 fanout1945 (.A(net1946),
    .X(net1945));
 sg13g2_buf_8 fanout1946 (.A(_02142_),
    .X(net1946));
 sg13g2_buf_8 fanout1947 (.A(net1951),
    .X(net1947));
 sg13g2_buf_8 fanout1948 (.A(net1951),
    .X(net1948));
 sg13g2_buf_8 fanout1949 (.A(net1951),
    .X(net1949));
 sg13g2_buf_1 fanout1950 (.A(net1951),
    .X(net1950));
 sg13g2_buf_8 fanout1951 (.A(_02109_),
    .X(net1951));
 sg13g2_buf_8 fanout1952 (.A(net1954),
    .X(net1952));
 sg13g2_buf_1 fanout1953 (.A(net1954),
    .X(net1953));
 sg13g2_buf_8 fanout1954 (.A(_02109_),
    .X(net1954));
 sg13g2_buf_8 fanout1955 (.A(net1957),
    .X(net1955));
 sg13g2_buf_1 fanout1956 (.A(net1957),
    .X(net1956));
 sg13g2_buf_8 fanout1957 (.A(_02109_),
    .X(net1957));
 sg13g2_buf_8 fanout1958 (.A(net1959),
    .X(net1958));
 sg13g2_buf_8 fanout1959 (.A(net1962),
    .X(net1959));
 sg13g2_buf_8 fanout1960 (.A(net1961),
    .X(net1960));
 sg13g2_buf_8 fanout1961 (.A(net1962),
    .X(net1961));
 sg13g2_buf_8 fanout1962 (.A(_01994_),
    .X(net1962));
 sg13g2_buf_8 fanout1963 (.A(net1967),
    .X(net1963));
 sg13g2_buf_8 fanout1964 (.A(net1967),
    .X(net1964));
 sg13g2_buf_8 fanout1965 (.A(net1966),
    .X(net1965));
 sg13g2_buf_8 fanout1966 (.A(net1967),
    .X(net1966));
 sg13g2_buf_8 fanout1967 (.A(_01994_),
    .X(net1967));
 sg13g2_buf_8 fanout1968 (.A(net1969),
    .X(net1968));
 sg13g2_buf_8 fanout1969 (.A(net1972),
    .X(net1969));
 sg13g2_buf_8 fanout1970 (.A(net1972),
    .X(net1970));
 sg13g2_buf_1 fanout1971 (.A(net1972),
    .X(net1971));
 sg13g2_buf_8 fanout1972 (.A(net1978),
    .X(net1972));
 sg13g2_buf_8 fanout1973 (.A(net1975),
    .X(net1973));
 sg13g2_buf_1 fanout1974 (.A(net1975),
    .X(net1974));
 sg13g2_buf_8 fanout1975 (.A(net1978),
    .X(net1975));
 sg13g2_buf_8 fanout1976 (.A(net1977),
    .X(net1976));
 sg13g2_buf_8 fanout1977 (.A(net1978),
    .X(net1977));
 sg13g2_buf_8 fanout1978 (.A(_01959_),
    .X(net1978));
 sg13g2_buf_8 fanout1979 (.A(net1981),
    .X(net1979));
 sg13g2_buf_1 fanout1980 (.A(net1981),
    .X(net1980));
 sg13g2_buf_8 fanout1981 (.A(net1989),
    .X(net1981));
 sg13g2_buf_8 fanout1982 (.A(net1989),
    .X(net1982));
 sg13g2_buf_1 fanout1983 (.A(net1989),
    .X(net1983));
 sg13g2_buf_8 fanout1984 (.A(net1988),
    .X(net1984));
 sg13g2_buf_8 fanout1985 (.A(net1988),
    .X(net1985));
 sg13g2_buf_8 fanout1986 (.A(net1988),
    .X(net1986));
 sg13g2_buf_8 fanout1987 (.A(net1988),
    .X(net1987));
 sg13g2_buf_8 fanout1988 (.A(net1989),
    .X(net1988));
 sg13g2_buf_8 fanout1989 (.A(_01926_),
    .X(net1989));
 sg13g2_buf_8 fanout1990 (.A(net1991),
    .X(net1990));
 sg13g2_buf_8 fanout1991 (.A(net1994),
    .X(net1991));
 sg13g2_buf_8 fanout1992 (.A(net1994),
    .X(net1992));
 sg13g2_buf_1 fanout1993 (.A(net1994),
    .X(net1993));
 sg13g2_buf_8 fanout1994 (.A(net2000),
    .X(net1994));
 sg13g2_buf_8 fanout1995 (.A(net1997),
    .X(net1995));
 sg13g2_buf_8 fanout1996 (.A(net1997),
    .X(net1996));
 sg13g2_buf_8 fanout1997 (.A(net2000),
    .X(net1997));
 sg13g2_buf_8 fanout1998 (.A(net2000),
    .X(net1998));
 sg13g2_buf_8 fanout1999 (.A(net2000),
    .X(net1999));
 sg13g2_buf_8 fanout2000 (.A(_01893_),
    .X(net2000));
 sg13g2_buf_8 fanout2001 (.A(net2003),
    .X(net2001));
 sg13g2_buf_1 fanout2002 (.A(net2003),
    .X(net2002));
 sg13g2_buf_8 fanout2003 (.A(net2011),
    .X(net2003));
 sg13g2_buf_8 fanout2004 (.A(net2011),
    .X(net2004));
 sg13g2_buf_1 fanout2005 (.A(net2011),
    .X(net2005));
 sg13g2_buf_8 fanout2006 (.A(net2010),
    .X(net2006));
 sg13g2_buf_8 fanout2007 (.A(net2010),
    .X(net2007));
 sg13g2_buf_8 fanout2008 (.A(net2010),
    .X(net2008));
 sg13g2_buf_8 fanout2009 (.A(net2010),
    .X(net2009));
 sg13g2_buf_8 fanout2010 (.A(net2011),
    .X(net2010));
 sg13g2_buf_8 fanout2011 (.A(_01860_),
    .X(net2011));
 sg13g2_buf_8 fanout2012 (.A(net2016),
    .X(net2012));
 sg13g2_buf_8 fanout2013 (.A(net2016),
    .X(net2013));
 sg13g2_buf_8 fanout2014 (.A(net2016),
    .X(net2014));
 sg13g2_buf_8 fanout2015 (.A(net2016),
    .X(net2015));
 sg13g2_buf_8 fanout2016 (.A(net2022),
    .X(net2016));
 sg13g2_buf_8 fanout2017 (.A(net2019),
    .X(net2017));
 sg13g2_buf_8 fanout2018 (.A(net2019),
    .X(net2018));
 sg13g2_buf_8 fanout2019 (.A(net2022),
    .X(net2019));
 sg13g2_buf_8 fanout2020 (.A(net2022),
    .X(net2020));
 sg13g2_buf_8 fanout2021 (.A(net2022),
    .X(net2021));
 sg13g2_buf_8 fanout2022 (.A(_01827_),
    .X(net2022));
 sg13g2_buf_8 fanout2023 (.A(net2025),
    .X(net2023));
 sg13g2_buf_1 fanout2024 (.A(net2025),
    .X(net2024));
 sg13g2_buf_8 fanout2025 (.A(net2028),
    .X(net2025));
 sg13g2_buf_8 fanout2026 (.A(net2028),
    .X(net2026));
 sg13g2_buf_1 fanout2027 (.A(net2028),
    .X(net2027));
 sg13g2_buf_8 fanout2028 (.A(_01752_),
    .X(net2028));
 sg13g2_buf_8 fanout2029 (.A(net2033),
    .X(net2029));
 sg13g2_buf_8 fanout2030 (.A(net2033),
    .X(net2030));
 sg13g2_buf_8 fanout2031 (.A(net2032),
    .X(net2031));
 sg13g2_buf_8 fanout2032 (.A(net2033),
    .X(net2032));
 sg13g2_buf_8 fanout2033 (.A(_01752_),
    .X(net2033));
 sg13g2_buf_8 fanout2034 (.A(net2038),
    .X(net2034));
 sg13g2_buf_8 fanout2035 (.A(net2038),
    .X(net2035));
 sg13g2_buf_8 fanout2036 (.A(net2038),
    .X(net2036));
 sg13g2_buf_8 fanout2037 (.A(net2038),
    .X(net2037));
 sg13g2_buf_8 fanout2038 (.A(net2044),
    .X(net2038));
 sg13g2_buf_8 fanout2039 (.A(net2044),
    .X(net2039));
 sg13g2_buf_8 fanout2040 (.A(net2044),
    .X(net2040));
 sg13g2_buf_8 fanout2041 (.A(net2042),
    .X(net2041));
 sg13g2_buf_8 fanout2042 (.A(net2043),
    .X(net2042));
 sg13g2_buf_8 fanout2043 (.A(net2044),
    .X(net2043));
 sg13g2_buf_8 fanout2044 (.A(_01717_),
    .X(net2044));
 sg13g2_buf_8 fanout2045 (.A(net2046),
    .X(net2045));
 sg13g2_buf_8 fanout2046 (.A(net2049),
    .X(net2046));
 sg13g2_buf_8 fanout2047 (.A(net2048),
    .X(net2047));
 sg13g2_buf_8 fanout2048 (.A(net2049),
    .X(net2048));
 sg13g2_buf_8 fanout2049 (.A(_01680_),
    .X(net2049));
 sg13g2_buf_8 fanout2050 (.A(net2054),
    .X(net2050));
 sg13g2_buf_8 fanout2051 (.A(net2054),
    .X(net2051));
 sg13g2_buf_8 fanout2052 (.A(net2053),
    .X(net2052));
 sg13g2_buf_8 fanout2053 (.A(net2054),
    .X(net2053));
 sg13g2_buf_8 fanout2054 (.A(_01680_),
    .X(net2054));
 sg13g2_buf_8 fanout2055 (.A(net2056),
    .X(net2055));
 sg13g2_buf_8 fanout2056 (.A(net2064),
    .X(net2056));
 sg13g2_buf_8 fanout2057 (.A(net2058),
    .X(net2057));
 sg13g2_buf_8 fanout2058 (.A(net2064),
    .X(net2058));
 sg13g2_buf_8 fanout2059 (.A(net2063),
    .X(net2059));
 sg13g2_buf_8 fanout2060 (.A(net2063),
    .X(net2060));
 sg13g2_buf_8 fanout2061 (.A(net2063),
    .X(net2061));
 sg13g2_buf_8 fanout2062 (.A(net2063),
    .X(net2062));
 sg13g2_buf_8 fanout2063 (.A(net2064),
    .X(net2063));
 sg13g2_buf_8 fanout2064 (.A(_01617_),
    .X(net2064));
 sg13g2_buf_8 fanout2065 (.A(net2066),
    .X(net2065));
 sg13g2_buf_8 fanout2066 (.A(_03817_),
    .X(net2066));
 sg13g2_buf_8 fanout2067 (.A(net2071),
    .X(net2067));
 sg13g2_buf_8 fanout2068 (.A(net2071),
    .X(net2068));
 sg13g2_buf_8 fanout2069 (.A(net2071),
    .X(net2069));
 sg13g2_buf_8 fanout2070 (.A(net2071),
    .X(net2070));
 sg13g2_buf_8 fanout2071 (.A(_02542_),
    .X(net2071));
 sg13g2_buf_8 fanout2072 (.A(net2076),
    .X(net2072));
 sg13g2_buf_8 fanout2073 (.A(net2076),
    .X(net2073));
 sg13g2_buf_8 fanout2074 (.A(net2076),
    .X(net2074));
 sg13g2_buf_8 fanout2075 (.A(net2076),
    .X(net2075));
 sg13g2_buf_8 fanout2076 (.A(_02342_),
    .X(net2076));
 sg13g2_buf_8 fanout2077 (.A(net2081),
    .X(net2077));
 sg13g2_buf_8 fanout2078 (.A(net2081),
    .X(net2078));
 sg13g2_buf_8 fanout2079 (.A(net2081),
    .X(net2079));
 sg13g2_buf_8 fanout2080 (.A(net2081),
    .X(net2080));
 sg13g2_buf_8 fanout2081 (.A(_01993_),
    .X(net2081));
 sg13g2_buf_8 fanout2082 (.A(net2086),
    .X(net2082));
 sg13g2_buf_8 fanout2083 (.A(net2086),
    .X(net2083));
 sg13g2_buf_8 fanout2084 (.A(net2085),
    .X(net2084));
 sg13g2_buf_8 fanout2085 (.A(net2086),
    .X(net2085));
 sg13g2_buf_8 fanout2086 (.A(_01826_),
    .X(net2086));
 sg13g2_buf_8 fanout2087 (.A(net2088),
    .X(net2087));
 sg13g2_buf_8 fanout2088 (.A(net2096),
    .X(net2088));
 sg13g2_buf_8 fanout2089 (.A(net2090),
    .X(net2089));
 sg13g2_buf_8 fanout2090 (.A(net2096),
    .X(net2090));
 sg13g2_buf_8 fanout2091 (.A(net2095),
    .X(net2091));
 sg13g2_buf_8 fanout2092 (.A(net2095),
    .X(net2092));
 sg13g2_buf_8 fanout2093 (.A(net2095),
    .X(net2093));
 sg13g2_buf_8 fanout2094 (.A(net2095),
    .X(net2094));
 sg13g2_buf_8 fanout2095 (.A(net2096),
    .X(net2095));
 sg13g2_buf_8 fanout2096 (.A(_01791_),
    .X(net2096));
 sg13g2_buf_8 fanout2097 (.A(net2101),
    .X(net2097));
 sg13g2_buf_8 fanout2098 (.A(net2101),
    .X(net2098));
 sg13g2_buf_8 fanout2099 (.A(net2101),
    .X(net2099));
 sg13g2_buf_8 fanout2100 (.A(net2101),
    .X(net2100));
 sg13g2_buf_8 fanout2101 (.A(_01714_),
    .X(net2101));
 sg13g2_buf_8 fanout2102 (.A(net2103),
    .X(net2102));
 sg13g2_buf_8 fanout2103 (.A(net2106),
    .X(net2103));
 sg13g2_buf_8 fanout2104 (.A(net2105),
    .X(net2104));
 sg13g2_buf_8 fanout2105 (.A(net2106),
    .X(net2105));
 sg13g2_buf_8 fanout2106 (.A(_01679_),
    .X(net2106));
 sg13g2_buf_8 fanout2107 (.A(net2110),
    .X(net2107));
 sg13g2_buf_8 fanout2108 (.A(net2110),
    .X(net2108));
 sg13g2_buf_8 fanout2109 (.A(net2110),
    .X(net2109));
 sg13g2_buf_8 fanout2110 (.A(_01548_),
    .X(net2110));
 sg13g2_buf_8 fanout2111 (.A(net2113),
    .X(net2111));
 sg13g2_buf_1 fanout2112 (.A(net2113),
    .X(net2112));
 sg13g2_buf_8 fanout2113 (.A(_01548_),
    .X(net2113));
 sg13g2_buf_8 fanout2114 (.A(net2116),
    .X(net2114));
 sg13g2_buf_2 fanout2115 (.A(net2116),
    .X(net2115));
 sg13g2_buf_8 fanout2116 (.A(_01548_),
    .X(net2116));
 sg13g2_buf_8 fanout2117 (.A(_03795_),
    .X(net2117));
 sg13g2_buf_2 fanout2118 (.A(net2122),
    .X(net2118));
 sg13g2_buf_8 fanout2119 (.A(net2121),
    .X(net2119));
 sg13g2_buf_1 fanout2120 (.A(net2121),
    .X(net2120));
 sg13g2_buf_1 fanout2121 (.A(net2122),
    .X(net2121));
 sg13g2_buf_8 fanout2122 (.A(net2126),
    .X(net2122));
 sg13g2_buf_2 fanout2123 (.A(net2125),
    .X(net2123));
 sg13g2_buf_2 fanout2124 (.A(net2125),
    .X(net2124));
 sg13g2_buf_2 fanout2125 (.A(net2126),
    .X(net2125));
 sg13g2_buf_1 fanout2126 (.A(_03677_),
    .X(net2126));
 sg13g2_buf_8 fanout2127 (.A(net2128),
    .X(net2127));
 sg13g2_buf_8 fanout2128 (.A(net2129),
    .X(net2128));
 sg13g2_buf_8 fanout2129 (.A(_02692_),
    .X(net2129));
 sg13g2_buf_8 fanout2130 (.A(net2132),
    .X(net2130));
 sg13g2_buf_2 fanout2131 (.A(net2132),
    .X(net2131));
 sg13g2_buf_8 fanout2132 (.A(net2135),
    .X(net2132));
 sg13g2_buf_8 fanout2133 (.A(net2135),
    .X(net2133));
 sg13g2_buf_1 fanout2134 (.A(net2135),
    .X(net2134));
 sg13g2_buf_8 fanout2135 (.A(net2151),
    .X(net2135));
 sg13g2_buf_8 fanout2136 (.A(net2138),
    .X(net2136));
 sg13g2_buf_8 fanout2137 (.A(net2138),
    .X(net2137));
 sg13g2_buf_8 fanout2138 (.A(net2141),
    .X(net2138));
 sg13g2_buf_8 fanout2139 (.A(net2141),
    .X(net2139));
 sg13g2_buf_8 fanout2140 (.A(net2141),
    .X(net2140));
 sg13g2_buf_8 fanout2141 (.A(net2151),
    .X(net2141));
 sg13g2_buf_8 fanout2142 (.A(net2146),
    .X(net2142));
 sg13g2_buf_1 fanout2143 (.A(net2146),
    .X(net2143));
 sg13g2_buf_8 fanout2144 (.A(net2146),
    .X(net2144));
 sg13g2_buf_8 fanout2145 (.A(net2146),
    .X(net2145));
 sg13g2_buf_8 fanout2146 (.A(net2151),
    .X(net2146));
 sg13g2_buf_8 fanout2147 (.A(net2150),
    .X(net2147));
 sg13g2_buf_8 fanout2148 (.A(net2149),
    .X(net2148));
 sg13g2_buf_8 fanout2149 (.A(net2150),
    .X(net2149));
 sg13g2_buf_8 fanout2150 (.A(net2151),
    .X(net2150));
 sg13g2_buf_8 fanout2151 (.A(net2173),
    .X(net2151));
 sg13g2_buf_8 fanout2152 (.A(net2155),
    .X(net2152));
 sg13g2_buf_8 fanout2153 (.A(net2155),
    .X(net2153));
 sg13g2_buf_8 fanout2154 (.A(net2155),
    .X(net2154));
 sg13g2_buf_8 fanout2155 (.A(net2161),
    .X(net2155));
 sg13g2_buf_8 fanout2156 (.A(net2158),
    .X(net2156));
 sg13g2_buf_8 fanout2157 (.A(net2161),
    .X(net2157));
 sg13g2_buf_1 fanout2158 (.A(net2161),
    .X(net2158));
 sg13g2_buf_8 fanout2159 (.A(net2160),
    .X(net2159));
 sg13g2_buf_8 fanout2160 (.A(net2161),
    .X(net2160));
 sg13g2_buf_8 fanout2161 (.A(net2173),
    .X(net2161));
 sg13g2_buf_8 fanout2162 (.A(net2163),
    .X(net2162));
 sg13g2_buf_8 fanout2163 (.A(net2166),
    .X(net2163));
 sg13g2_buf_8 fanout2164 (.A(net2165),
    .X(net2164));
 sg13g2_buf_8 fanout2165 (.A(net2166),
    .X(net2165));
 sg13g2_buf_8 fanout2166 (.A(net2173),
    .X(net2166));
 sg13g2_buf_8 fanout2167 (.A(net2168),
    .X(net2167));
 sg13g2_buf_8 fanout2168 (.A(net2172),
    .X(net2168));
 sg13g2_buf_8 fanout2169 (.A(net2171),
    .X(net2169));
 sg13g2_buf_8 fanout2170 (.A(net2171),
    .X(net2170));
 sg13g2_buf_8 fanout2171 (.A(net2172),
    .X(net2171));
 sg13g2_buf_8 fanout2172 (.A(net2173),
    .X(net2172));
 sg13g2_buf_8 fanout2173 (.A(_01750_),
    .X(net2173));
 sg13g2_buf_8 fanout2174 (.A(net2176),
    .X(net2174));
 sg13g2_buf_2 fanout2175 (.A(net2176),
    .X(net2175));
 sg13g2_buf_8 fanout2176 (.A(net2179),
    .X(net2176));
 sg13g2_buf_8 fanout2177 (.A(net2179),
    .X(net2177));
 sg13g2_buf_1 fanout2178 (.A(net2179),
    .X(net2178));
 sg13g2_buf_8 fanout2179 (.A(net2195),
    .X(net2179));
 sg13g2_buf_8 fanout2180 (.A(net2182),
    .X(net2180));
 sg13g2_buf_8 fanout2181 (.A(net2182),
    .X(net2181));
 sg13g2_buf_8 fanout2182 (.A(net2185),
    .X(net2182));
 sg13g2_buf_8 fanout2183 (.A(net2185),
    .X(net2183));
 sg13g2_buf_8 fanout2184 (.A(net2185),
    .X(net2184));
 sg13g2_buf_8 fanout2185 (.A(net2195),
    .X(net2185));
 sg13g2_buf_8 fanout2186 (.A(net2190),
    .X(net2186));
 sg13g2_buf_1 fanout2187 (.A(net2190),
    .X(net2187));
 sg13g2_buf_8 fanout2188 (.A(net2190),
    .X(net2188));
 sg13g2_buf_8 fanout2189 (.A(net2190),
    .X(net2189));
 sg13g2_buf_8 fanout2190 (.A(net2195),
    .X(net2190));
 sg13g2_buf_8 fanout2191 (.A(net2194),
    .X(net2191));
 sg13g2_buf_8 fanout2192 (.A(net2193),
    .X(net2192));
 sg13g2_buf_8 fanout2193 (.A(net2194),
    .X(net2193));
 sg13g2_buf_8 fanout2194 (.A(net2195),
    .X(net2194));
 sg13g2_buf_8 fanout2195 (.A(net2217),
    .X(net2195));
 sg13g2_buf_8 fanout2196 (.A(net2197),
    .X(net2196));
 sg13g2_buf_8 fanout2197 (.A(net2199),
    .X(net2197));
 sg13g2_buf_8 fanout2198 (.A(net2199),
    .X(net2198));
 sg13g2_buf_8 fanout2199 (.A(net2205),
    .X(net2199));
 sg13g2_buf_8 fanout2200 (.A(net2202),
    .X(net2200));
 sg13g2_buf_8 fanout2201 (.A(net2205),
    .X(net2201));
 sg13g2_buf_1 fanout2202 (.A(net2205),
    .X(net2202));
 sg13g2_buf_8 fanout2203 (.A(net2204),
    .X(net2203));
 sg13g2_buf_8 fanout2204 (.A(net2205),
    .X(net2204));
 sg13g2_buf_8 fanout2205 (.A(net2217),
    .X(net2205));
 sg13g2_buf_8 fanout2206 (.A(net2207),
    .X(net2206));
 sg13g2_buf_8 fanout2207 (.A(net2210),
    .X(net2207));
 sg13g2_buf_8 fanout2208 (.A(net2209),
    .X(net2208));
 sg13g2_buf_8 fanout2209 (.A(net2210),
    .X(net2209));
 sg13g2_buf_8 fanout2210 (.A(net2217),
    .X(net2210));
 sg13g2_buf_8 fanout2211 (.A(net2212),
    .X(net2211));
 sg13g2_buf_8 fanout2212 (.A(net2216),
    .X(net2212));
 sg13g2_buf_8 fanout2213 (.A(net2215),
    .X(net2213));
 sg13g2_buf_8 fanout2214 (.A(net2215),
    .X(net2214));
 sg13g2_buf_8 fanout2215 (.A(net2216),
    .X(net2215));
 sg13g2_buf_8 fanout2216 (.A(net2217),
    .X(net2216));
 sg13g2_buf_8 fanout2217 (.A(_01715_),
    .X(net2217));
 sg13g2_buf_8 fanout2218 (.A(net2220),
    .X(net2218));
 sg13g2_buf_2 fanout2219 (.A(net2220),
    .X(net2219));
 sg13g2_buf_8 fanout2220 (.A(net2223),
    .X(net2220));
 sg13g2_buf_8 fanout2221 (.A(net2223),
    .X(net2221));
 sg13g2_buf_8 fanout2222 (.A(net2223),
    .X(net2222));
 sg13g2_buf_8 fanout2223 (.A(net2238),
    .X(net2223));
 sg13g2_buf_8 fanout2224 (.A(net2225),
    .X(net2224));
 sg13g2_buf_8 fanout2225 (.A(net2228),
    .X(net2225));
 sg13g2_buf_8 fanout2226 (.A(net2228),
    .X(net2226));
 sg13g2_buf_8 fanout2227 (.A(net2228),
    .X(net2227));
 sg13g2_buf_8 fanout2228 (.A(net2238),
    .X(net2228));
 sg13g2_buf_8 fanout2229 (.A(net2232),
    .X(net2229));
 sg13g2_buf_8 fanout2230 (.A(net2232),
    .X(net2230));
 sg13g2_buf_8 fanout2231 (.A(net2232),
    .X(net2231));
 sg13g2_buf_8 fanout2232 (.A(net2238),
    .X(net2232));
 sg13g2_buf_8 fanout2233 (.A(net2237),
    .X(net2233));
 sg13g2_buf_8 fanout2234 (.A(net2236),
    .X(net2234));
 sg13g2_buf_8 fanout2235 (.A(net2236),
    .X(net2235));
 sg13g2_buf_8 fanout2236 (.A(net2237),
    .X(net2236));
 sg13g2_buf_8 fanout2237 (.A(net2238),
    .X(net2237));
 sg13g2_buf_8 fanout2238 (.A(_01615_),
    .X(net2238));
 sg13g2_buf_8 fanout2239 (.A(net2242),
    .X(net2239));
 sg13g2_buf_8 fanout2240 (.A(net2242),
    .X(net2240));
 sg13g2_buf_8 fanout2241 (.A(net2242),
    .X(net2241));
 sg13g2_buf_8 fanout2242 (.A(net2259),
    .X(net2242));
 sg13g2_buf_8 fanout2243 (.A(net2247),
    .X(net2243));
 sg13g2_buf_8 fanout2244 (.A(net2247),
    .X(net2244));
 sg13g2_buf_8 fanout2245 (.A(net2246),
    .X(net2245));
 sg13g2_buf_8 fanout2246 (.A(net2247),
    .X(net2246));
 sg13g2_buf_8 fanout2247 (.A(net2259),
    .X(net2247));
 sg13g2_buf_8 fanout2248 (.A(net2249),
    .X(net2248));
 sg13g2_buf_8 fanout2249 (.A(net2252),
    .X(net2249));
 sg13g2_buf_8 fanout2250 (.A(net2252),
    .X(net2250));
 sg13g2_buf_8 fanout2251 (.A(net2252),
    .X(net2251));
 sg13g2_buf_8 fanout2252 (.A(net2259),
    .X(net2252));
 sg13g2_buf_8 fanout2253 (.A(net2258),
    .X(net2253));
 sg13g2_buf_8 fanout2254 (.A(net2258),
    .X(net2254));
 sg13g2_buf_8 fanout2255 (.A(net2257),
    .X(net2255));
 sg13g2_buf_8 fanout2256 (.A(net2257),
    .X(net2256));
 sg13g2_buf_8 fanout2257 (.A(net2258),
    .X(net2257));
 sg13g2_buf_8 fanout2258 (.A(net2259),
    .X(net2258));
 sg13g2_buf_8 fanout2259 (.A(_01615_),
    .X(net2259));
 sg13g2_buf_8 fanout2260 (.A(net2261),
    .X(net2260));
 sg13g2_buf_8 fanout2261 (.A(net2264),
    .X(net2261));
 sg13g2_buf_8 fanout2262 (.A(net2264),
    .X(net2262));
 sg13g2_buf_8 fanout2263 (.A(net2264),
    .X(net2263));
 sg13g2_buf_8 fanout2264 (.A(_01614_),
    .X(net2264));
 sg13g2_buf_8 fanout2265 (.A(net2267),
    .X(net2265));
 sg13g2_buf_2 fanout2266 (.A(net2267),
    .X(net2266));
 sg13g2_buf_8 fanout2267 (.A(net2270),
    .X(net2267));
 sg13g2_buf_8 fanout2268 (.A(net2270),
    .X(net2268));
 sg13g2_buf_8 fanout2269 (.A(net2270),
    .X(net2269));
 sg13g2_buf_8 fanout2270 (.A(net2284),
    .X(net2270));
 sg13g2_buf_8 fanout2271 (.A(net2272),
    .X(net2271));
 sg13g2_buf_8 fanout2272 (.A(net2275),
    .X(net2272));
 sg13g2_buf_8 fanout2273 (.A(net2275),
    .X(net2273));
 sg13g2_buf_8 fanout2274 (.A(net2275),
    .X(net2274));
 sg13g2_buf_8 fanout2275 (.A(net2284),
    .X(net2275));
 sg13g2_buf_8 fanout2276 (.A(net2279),
    .X(net2276));
 sg13g2_buf_8 fanout2277 (.A(net2279),
    .X(net2277));
 sg13g2_buf_8 fanout2278 (.A(net2279),
    .X(net2278));
 sg13g2_buf_8 fanout2279 (.A(net2284),
    .X(net2279));
 sg13g2_buf_8 fanout2280 (.A(net2283),
    .X(net2280));
 sg13g2_buf_8 fanout2281 (.A(net2282),
    .X(net2281));
 sg13g2_buf_8 fanout2282 (.A(net2283),
    .X(net2282));
 sg13g2_buf_8 fanout2283 (.A(net2284),
    .X(net2283));
 sg13g2_buf_8 fanout2284 (.A(net2306),
    .X(net2284));
 sg13g2_buf_8 fanout2285 (.A(net2288),
    .X(net2285));
 sg13g2_buf_8 fanout2286 (.A(net2288),
    .X(net2286));
 sg13g2_buf_8 fanout2287 (.A(net2288),
    .X(net2287));
 sg13g2_buf_8 fanout2288 (.A(net2306),
    .X(net2288));
 sg13g2_buf_8 fanout2289 (.A(net2293),
    .X(net2289));
 sg13g2_buf_8 fanout2290 (.A(net2293),
    .X(net2290));
 sg13g2_buf_8 fanout2291 (.A(net2292),
    .X(net2291));
 sg13g2_buf_8 fanout2292 (.A(net2293),
    .X(net2292));
 sg13g2_buf_8 fanout2293 (.A(net2306),
    .X(net2293));
 sg13g2_buf_8 fanout2294 (.A(net2295),
    .X(net2294));
 sg13g2_buf_8 fanout2295 (.A(net2305),
    .X(net2295));
 sg13g2_buf_8 fanout2296 (.A(net2298),
    .X(net2296));
 sg13g2_buf_8 fanout2297 (.A(net2298),
    .X(net2297));
 sg13g2_buf_8 fanout2298 (.A(net2305),
    .X(net2298));
 sg13g2_buf_8 fanout2299 (.A(net2304),
    .X(net2299));
 sg13g2_buf_8 fanout2300 (.A(net2304),
    .X(net2300));
 sg13g2_buf_8 fanout2301 (.A(net2303),
    .X(net2301));
 sg13g2_buf_8 fanout2302 (.A(net2303),
    .X(net2302));
 sg13g2_buf_8 fanout2303 (.A(net2304),
    .X(net2303));
 sg13g2_buf_8 fanout2304 (.A(net2305),
    .X(net2304));
 sg13g2_buf_8 fanout2305 (.A(net2306),
    .X(net2305));
 sg13g2_buf_8 fanout2306 (.A(_01546_),
    .X(net2306));
 sg13g2_buf_8 fanout2307 (.A(net2312),
    .X(net2307));
 sg13g2_buf_8 fanout2308 (.A(net2312),
    .X(net2308));
 sg13g2_buf_8 fanout2309 (.A(net2311),
    .X(net2309));
 sg13g2_buf_8 fanout2310 (.A(net2311),
    .X(net2310));
 sg13g2_buf_8 fanout2311 (.A(net2312),
    .X(net2311));
 sg13g2_buf_8 fanout2312 (.A(_01539_),
    .X(net2312));
 sg13g2_buf_8 fanout2313 (.A(_03794_),
    .X(net2313));
 sg13g2_buf_8 fanout2314 (.A(net2315),
    .X(net2314));
 sg13g2_buf_8 fanout2315 (.A(_03766_),
    .X(net2315));
 sg13g2_buf_8 fanout2316 (.A(net2317),
    .X(net2316));
 sg13g2_buf_8 fanout2317 (.A(net2318),
    .X(net2317));
 sg13g2_buf_2 fanout2318 (.A(_02691_),
    .X(net2318));
 sg13g2_buf_8 fanout2319 (.A(net2320),
    .X(net2319));
 sg13g2_buf_2 fanout2320 (.A(net2321),
    .X(net2320));
 sg13g2_buf_1 fanout2321 (.A(net2324),
    .X(net2321));
 sg13g2_buf_8 fanout2322 (.A(net2324),
    .X(net2322));
 sg13g2_buf_1 fanout2323 (.A(net2324),
    .X(net2323));
 sg13g2_buf_8 fanout2324 (.A(_02030_),
    .X(net2324));
 sg13g2_buf_8 fanout2325 (.A(_01533_),
    .X(net2325));
 sg13g2_buf_8 fanout2326 (.A(net2328),
    .X(net2326));
 sg13g2_buf_8 fanout2327 (.A(net2328),
    .X(net2327));
 sg13g2_buf_8 fanout2328 (.A(net2329),
    .X(net2328));
 sg13g2_buf_8 fanout2329 (.A(_01470_),
    .X(net2329));
 sg13g2_buf_8 fanout2330 (.A(_01470_),
    .X(net2330));
 sg13g2_buf_8 fanout2331 (.A(_01470_),
    .X(net2331));
 sg13g2_buf_8 fanout2332 (.A(net2333),
    .X(net2332));
 sg13g2_buf_8 fanout2333 (.A(net2334),
    .X(net2333));
 sg13g2_buf_2 fanout2334 (.A(net2335),
    .X(net2334));
 sg13g2_buf_1 fanout2335 (.A(net2337),
    .X(net2335));
 sg13g2_buf_8 fanout2336 (.A(net2337),
    .X(net2336));
 sg13g2_buf_8 fanout2337 (.A(_03884_),
    .X(net2337));
 sg13g2_buf_8 fanout2338 (.A(net2340),
    .X(net2338));
 sg13g2_buf_1 fanout2339 (.A(net2340),
    .X(net2339));
 sg13g2_buf_8 fanout2340 (.A(net2341),
    .X(net2340));
 sg13g2_buf_8 fanout2341 (.A(net2343),
    .X(net2341));
 sg13g2_buf_8 fanout2342 (.A(net2343),
    .X(net2342));
 sg13g2_buf_8 fanout2343 (.A(_03641_),
    .X(net2343));
 sg13g2_buf_8 fanout2344 (.A(net2347),
    .X(net2344));
 sg13g2_buf_1 fanout2345 (.A(net2347),
    .X(net2345));
 sg13g2_buf_8 fanout2346 (.A(net2347),
    .X(net2346));
 sg13g2_buf_8 fanout2347 (.A(_00471_),
    .X(net2347));
 sg13g2_buf_8 fanout2348 (.A(net2349),
    .X(net2348));
 sg13g2_buf_8 fanout2349 (.A(net2350),
    .X(net2349));
 sg13g2_buf_8 fanout2350 (.A(_00471_),
    .X(net2350));
 sg13g2_buf_8 fanout2351 (.A(net2352),
    .X(net2351));
 sg13g2_buf_8 fanout2352 (.A(net2353),
    .X(net2352));
 sg13g2_buf_8 fanout2353 (.A(_02680_),
    .X(net2353));
 sg13g2_buf_8 fanout2354 (.A(net2355),
    .X(net2354));
 sg13g2_buf_2 fanout2355 (.A(net2356),
    .X(net2355));
 sg13g2_buf_1 fanout2356 (.A(net2357),
    .X(net2356));
 sg13g2_buf_2 fanout2357 (.A(_02680_),
    .X(net2357));
 sg13g2_buf_8 fanout2358 (.A(net2359),
    .X(net2358));
 sg13g2_buf_8 fanout2359 (.A(net2360),
    .X(net2359));
 sg13g2_buf_8 fanout2360 (.A(_01415_),
    .X(net2360));
 sg13g2_buf_8 fanout2361 (.A(net2362),
    .X(net2361));
 sg13g2_buf_2 fanout2362 (.A(_01415_),
    .X(net2362));
 sg13g2_buf_8 fanout2363 (.A(net2364),
    .X(net2363));
 sg13g2_buf_8 fanout2364 (.A(net2366),
    .X(net2364));
 sg13g2_buf_8 fanout2365 (.A(net2366),
    .X(net2365));
 sg13g2_buf_8 fanout2366 (.A(_02683_),
    .X(net2366));
 sg13g2_buf_8 fanout2367 (.A(net2368),
    .X(net2367));
 sg13g2_buf_2 fanout2368 (.A(_01460_),
    .X(net2368));
 sg13g2_buf_8 fanout2369 (.A(net2370),
    .X(net2369));
 sg13g2_buf_8 fanout2370 (.A(net2371),
    .X(net2370));
 sg13g2_buf_8 fanout2371 (.A(_03718_),
    .X(net2371));
 sg13g2_buf_8 fanout2372 (.A(net2373),
    .X(net2372));
 sg13g2_buf_8 fanout2373 (.A(_01673_),
    .X(net2373));
 sg13g2_buf_8 fanout2374 (.A(net2375),
    .X(net2374));
 sg13g2_buf_8 fanout2375 (.A(_01670_),
    .X(net2375));
 sg13g2_buf_8 fanout2376 (.A(_01455_),
    .X(net2376));
 sg13g2_buf_8 fanout2377 (.A(net2378),
    .X(net2377));
 sg13g2_buf_8 fanout2378 (.A(net2379),
    .X(net2378));
 sg13g2_buf_8 fanout2379 (.A(_01404_),
    .X(net2379));
 sg13g2_buf_8 fanout2380 (.A(net2383),
    .X(net2380));
 sg13g2_buf_8 fanout2381 (.A(net2383),
    .X(net2381));
 sg13g2_buf_8 fanout2382 (.A(net2383),
    .X(net2382));
 sg13g2_buf_8 fanout2383 (.A(_01404_),
    .X(net2383));
 sg13g2_buf_8 fanout2384 (.A(net2388),
    .X(net2384));
 sg13g2_buf_8 fanout2385 (.A(net2388),
    .X(net2385));
 sg13g2_buf_8 fanout2386 (.A(net2387),
    .X(net2386));
 sg13g2_buf_8 fanout2387 (.A(net2388),
    .X(net2387));
 sg13g2_buf_8 fanout2388 (.A(net3769),
    .X(net2388));
 sg13g2_buf_8 fanout2389 (.A(net2390),
    .X(net2389));
 sg13g2_buf_8 fanout2390 (.A(_01669_),
    .X(net2390));
 sg13g2_buf_8 fanout2391 (.A(_01656_),
    .X(net2391));
 sg13g2_buf_8 fanout2392 (.A(_01656_),
    .X(net2392));
 sg13g2_buf_8 fanout2393 (.A(net2394),
    .X(net2393));
 sg13g2_buf_8 fanout2394 (.A(_01655_),
    .X(net2394));
 sg13g2_buf_8 fanout2395 (.A(_01654_),
    .X(net2395));
 sg13g2_buf_8 fanout2396 (.A(_01653_),
    .X(net2396));
 sg13g2_buf_8 fanout2397 (.A(net2398),
    .X(net2397));
 sg13g2_buf_8 fanout2398 (.A(net2401),
    .X(net2398));
 sg13g2_buf_8 fanout2399 (.A(net2400),
    .X(net2399));
 sg13g2_buf_8 fanout2400 (.A(net2401),
    .X(net2400));
 sg13g2_buf_8 fanout2401 (.A(_01611_),
    .X(net2401));
 sg13g2_buf_8 fanout2402 (.A(net2404),
    .X(net2402));
 sg13g2_buf_8 fanout2403 (.A(net2407),
    .X(net2403));
 sg13g2_buf_1 fanout2404 (.A(net2407),
    .X(net2404));
 sg13g2_buf_8 fanout2405 (.A(net2407),
    .X(net2405));
 sg13g2_buf_1 fanout2406 (.A(net2407),
    .X(net2406));
 sg13g2_buf_2 fanout2407 (.A(_01609_),
    .X(net2407));
 sg13g2_buf_8 fanout2408 (.A(net2410),
    .X(net2408));
 sg13g2_buf_1 fanout2409 (.A(net2410),
    .X(net2409));
 sg13g2_buf_8 fanout2410 (.A(_01607_),
    .X(net2410));
 sg13g2_buf_8 fanout2411 (.A(net2412),
    .X(net2411));
 sg13g2_buf_8 fanout2412 (.A(_01607_),
    .X(net2412));
 sg13g2_buf_8 fanout2413 (.A(net2417),
    .X(net2413));
 sg13g2_buf_2 fanout2414 (.A(net2417),
    .X(net2414));
 sg13g2_buf_8 fanout2415 (.A(net2416),
    .X(net2415));
 sg13g2_buf_8 fanout2416 (.A(net2417),
    .X(net2416));
 sg13g2_buf_8 fanout2417 (.A(_01605_),
    .X(net2417));
 sg13g2_buf_8 fanout2418 (.A(net2422),
    .X(net2418));
 sg13g2_buf_2 fanout2419 (.A(net2422),
    .X(net2419));
 sg13g2_buf_8 fanout2420 (.A(net2422),
    .X(net2420));
 sg13g2_buf_8 fanout2421 (.A(net2422),
    .X(net2421));
 sg13g2_buf_8 fanout2422 (.A(_01603_),
    .X(net2422));
 sg13g2_buf_8 fanout2423 (.A(net2425),
    .X(net2423));
 sg13g2_buf_1 fanout2424 (.A(net2425),
    .X(net2424));
 sg13g2_buf_8 fanout2425 (.A(_01601_),
    .X(net2425));
 sg13g2_buf_8 fanout2426 (.A(net2427),
    .X(net2426));
 sg13g2_buf_8 fanout2427 (.A(_01601_),
    .X(net2427));
 sg13g2_buf_8 fanout2428 (.A(net2433),
    .X(net2428));
 sg13g2_buf_8 fanout2429 (.A(net2430),
    .X(net2429));
 sg13g2_buf_1 fanout2430 (.A(net2433),
    .X(net2430));
 sg13g2_buf_8 fanout2431 (.A(net2433),
    .X(net2431));
 sg13g2_buf_1 fanout2432 (.A(net2433),
    .X(net2432));
 sg13g2_buf_8 fanout2433 (.A(_01599_),
    .X(net2433));
 sg13g2_buf_8 fanout2434 (.A(net2435),
    .X(net2434));
 sg13g2_buf_8 fanout2435 (.A(_01597_),
    .X(net2435));
 sg13g2_buf_8 fanout2436 (.A(net2438),
    .X(net2436));
 sg13g2_buf_1 fanout2437 (.A(net2438),
    .X(net2437));
 sg13g2_buf_8 fanout2438 (.A(_01597_),
    .X(net2438));
 sg13g2_buf_8 fanout2439 (.A(net2440),
    .X(net2439));
 sg13g2_buf_8 fanout2440 (.A(_01595_),
    .X(net2440));
 sg13g2_buf_8 fanout2441 (.A(net2442),
    .X(net2441));
 sg13g2_buf_8 fanout2442 (.A(_01595_),
    .X(net2442));
 sg13g2_buf_1 fanout2443 (.A(_01595_),
    .X(net2443));
 sg13g2_buf_8 fanout2444 (.A(net2449),
    .X(net2444));
 sg13g2_buf_1 fanout2445 (.A(net2449),
    .X(net2445));
 sg13g2_buf_8 fanout2446 (.A(net2449),
    .X(net2446));
 sg13g2_buf_8 fanout2447 (.A(net2449),
    .X(net2447));
 sg13g2_buf_1 fanout2448 (.A(net2449),
    .X(net2448));
 sg13g2_buf_8 fanout2449 (.A(_01593_),
    .X(net2449));
 sg13g2_buf_8 fanout2450 (.A(net2452),
    .X(net2450));
 sg13g2_buf_8 fanout2451 (.A(net2452),
    .X(net2451));
 sg13g2_buf_2 fanout2452 (.A(_01591_),
    .X(net2452));
 sg13g2_buf_8 fanout2453 (.A(_01591_),
    .X(net2453));
 sg13g2_buf_2 fanout2454 (.A(_01591_),
    .X(net2454));
 sg13g2_buf_8 fanout2455 (.A(net2457),
    .X(net2455));
 sg13g2_buf_8 fanout2456 (.A(net2457),
    .X(net2456));
 sg13g2_buf_8 fanout2457 (.A(_01589_),
    .X(net2457));
 sg13g2_buf_8 fanout2458 (.A(net2459),
    .X(net2458));
 sg13g2_buf_8 fanout2459 (.A(_01589_),
    .X(net2459));
 sg13g2_buf_8 fanout2460 (.A(net2464),
    .X(net2460));
 sg13g2_buf_8 fanout2461 (.A(net2464),
    .X(net2461));
 sg13g2_buf_8 fanout2462 (.A(net2464),
    .X(net2462));
 sg13g2_buf_8 fanout2463 (.A(net2464),
    .X(net2463));
 sg13g2_buf_8 fanout2464 (.A(_01587_),
    .X(net2464));
 sg13g2_buf_8 fanout2465 (.A(net2469),
    .X(net2465));
 sg13g2_buf_8 fanout2466 (.A(net2469),
    .X(net2466));
 sg13g2_buf_8 fanout2467 (.A(net2468),
    .X(net2467));
 sg13g2_buf_8 fanout2468 (.A(net2469),
    .X(net2468));
 sg13g2_buf_8 fanout2469 (.A(_01585_),
    .X(net2469));
 sg13g2_buf_8 fanout2470 (.A(net2472),
    .X(net2470));
 sg13g2_buf_8 fanout2471 (.A(net2472),
    .X(net2471));
 sg13g2_buf_2 fanout2472 (.A(_01583_),
    .X(net2472));
 sg13g2_buf_8 fanout2473 (.A(_01583_),
    .X(net2473));
 sg13g2_buf_2 fanout2474 (.A(_01583_),
    .X(net2474));
 sg13g2_buf_8 fanout2475 (.A(net2477),
    .X(net2475));
 sg13g2_buf_1 fanout2476 (.A(net2477),
    .X(net2476));
 sg13g2_buf_2 fanout2477 (.A(_01581_),
    .X(net2477));
 sg13g2_buf_8 fanout2478 (.A(net2480),
    .X(net2478));
 sg13g2_buf_1 fanout2479 (.A(net2480),
    .X(net2479));
 sg13g2_buf_8 fanout2480 (.A(_01581_),
    .X(net2480));
 sg13g2_buf_8 fanout2481 (.A(net2482),
    .X(net2481));
 sg13g2_buf_8 fanout2482 (.A(net2485),
    .X(net2482));
 sg13g2_buf_8 fanout2483 (.A(net2484),
    .X(net2483));
 sg13g2_buf_8 fanout2484 (.A(net2485),
    .X(net2484));
 sg13g2_buf_8 fanout2485 (.A(_01579_),
    .X(net2485));
 sg13g2_buf_8 fanout2486 (.A(net2487),
    .X(net2486));
 sg13g2_buf_8 fanout2487 (.A(net2490),
    .X(net2487));
 sg13g2_buf_8 fanout2488 (.A(net2490),
    .X(net2488));
 sg13g2_buf_2 fanout2489 (.A(net2490),
    .X(net2489));
 sg13g2_buf_8 fanout2490 (.A(_01577_),
    .X(net2490));
 sg13g2_buf_8 fanout2491 (.A(net2495),
    .X(net2491));
 sg13g2_buf_8 fanout2492 (.A(net2495),
    .X(net2492));
 sg13g2_buf_8 fanout2493 (.A(net2494),
    .X(net2493));
 sg13g2_buf_8 fanout2494 (.A(net2495),
    .X(net2494));
 sg13g2_buf_8 fanout2495 (.A(_01575_),
    .X(net2495));
 sg13g2_buf_8 fanout2496 (.A(net2498),
    .X(net2496));
 sg13g2_buf_1 fanout2497 (.A(net2498),
    .X(net2497));
 sg13g2_buf_1 fanout2498 (.A(_01573_),
    .X(net2498));
 sg13g2_buf_8 fanout2499 (.A(net2501),
    .X(net2499));
 sg13g2_buf_1 fanout2500 (.A(net2501),
    .X(net2500));
 sg13g2_buf_8 fanout2501 (.A(_01573_),
    .X(net2501));
 sg13g2_buf_8 fanout2502 (.A(net2503),
    .X(net2502));
 sg13g2_buf_8 fanout2503 (.A(net2506),
    .X(net2503));
 sg13g2_buf_8 fanout2504 (.A(net2506),
    .X(net2504));
 sg13g2_buf_8 fanout2505 (.A(net2506),
    .X(net2505));
 sg13g2_buf_8 fanout2506 (.A(_01571_),
    .X(net2506));
 sg13g2_buf_8 fanout2507 (.A(_01569_),
    .X(net2507));
 sg13g2_buf_8 fanout2508 (.A(_01569_),
    .X(net2508));
 sg13g2_buf_8 fanout2509 (.A(net2511),
    .X(net2509));
 sg13g2_buf_1 fanout2510 (.A(net2511),
    .X(net2510));
 sg13g2_buf_8 fanout2511 (.A(_01569_),
    .X(net2511));
 sg13g2_buf_8 fanout2512 (.A(net2513),
    .X(net2512));
 sg13g2_buf_8 fanout2513 (.A(net2517),
    .X(net2513));
 sg13g2_buf_8 fanout2514 (.A(net2516),
    .X(net2514));
 sg13g2_buf_1 fanout2515 (.A(net2516),
    .X(net2515));
 sg13g2_buf_8 fanout2516 (.A(net2517),
    .X(net2516));
 sg13g2_buf_8 fanout2517 (.A(_01567_),
    .X(net2517));
 sg13g2_buf_8 fanout2518 (.A(_01565_),
    .X(net2518));
 sg13g2_buf_1 fanout2519 (.A(_01565_),
    .X(net2519));
 sg13g2_buf_8 fanout2520 (.A(net2522),
    .X(net2520));
 sg13g2_buf_8 fanout2521 (.A(net2522),
    .X(net2521));
 sg13g2_buf_8 fanout2522 (.A(_01565_),
    .X(net2522));
 sg13g2_buf_8 fanout2523 (.A(_01563_),
    .X(net2523));
 sg13g2_buf_1 fanout2524 (.A(_01563_),
    .X(net2524));
 sg13g2_buf_8 fanout2525 (.A(net2527),
    .X(net2525));
 sg13g2_buf_8 fanout2526 (.A(net2527),
    .X(net2526));
 sg13g2_buf_8 fanout2527 (.A(_01563_),
    .X(net2527));
 sg13g2_buf_8 fanout2528 (.A(net2529),
    .X(net2528));
 sg13g2_buf_8 fanout2529 (.A(net2532),
    .X(net2529));
 sg13g2_buf_8 fanout2530 (.A(net2531),
    .X(net2530));
 sg13g2_buf_8 fanout2531 (.A(net2532),
    .X(net2531));
 sg13g2_buf_8 fanout2532 (.A(_01561_),
    .X(net2532));
 sg13g2_buf_8 fanout2533 (.A(_01559_),
    .X(net2533));
 sg13g2_buf_8 fanout2534 (.A(_01559_),
    .X(net2534));
 sg13g2_buf_8 fanout2535 (.A(net2537),
    .X(net2535));
 sg13g2_buf_1 fanout2536 (.A(net2537),
    .X(net2536));
 sg13g2_buf_8 fanout2537 (.A(_01559_),
    .X(net2537));
 sg13g2_buf_8 fanout2538 (.A(net2540),
    .X(net2538));
 sg13g2_buf_1 fanout2539 (.A(net2540),
    .X(net2539));
 sg13g2_buf_8 fanout2540 (.A(_01557_),
    .X(net2540));
 sg13g2_buf_8 fanout2541 (.A(net2543),
    .X(net2541));
 sg13g2_buf_1 fanout2542 (.A(net2543),
    .X(net2542));
 sg13g2_buf_8 fanout2543 (.A(_01557_),
    .X(net2543));
 sg13g2_buf_8 fanout2544 (.A(net2549),
    .X(net2544));
 sg13g2_buf_1 fanout2545 (.A(net2549),
    .X(net2545));
 sg13g2_buf_8 fanout2546 (.A(net2547),
    .X(net2546));
 sg13g2_buf_8 fanout2547 (.A(net2549),
    .X(net2547));
 sg13g2_buf_8 fanout2548 (.A(net2549),
    .X(net2548));
 sg13g2_buf_8 fanout2549 (.A(_01555_),
    .X(net2549));
 sg13g2_buf_8 fanout2550 (.A(_01553_),
    .X(net2550));
 sg13g2_buf_8 fanout2551 (.A(_01553_),
    .X(net2551));
 sg13g2_buf_8 fanout2552 (.A(net2554),
    .X(net2552));
 sg13g2_buf_1 fanout2553 (.A(net2554),
    .X(net2553));
 sg13g2_buf_8 fanout2554 (.A(_01553_),
    .X(net2554));
 sg13g2_buf_8 fanout2555 (.A(net2556),
    .X(net2555));
 sg13g2_buf_8 fanout2556 (.A(net2559),
    .X(net2556));
 sg13g2_buf_8 fanout2557 (.A(net2558),
    .X(net2557));
 sg13g2_buf_8 fanout2558 (.A(net2559),
    .X(net2558));
 sg13g2_buf_8 fanout2559 (.A(_01551_),
    .X(net2559));
 sg13g2_buf_8 fanout2560 (.A(net2565),
    .X(net2560));
 sg13g2_buf_1 fanout2561 (.A(net2565),
    .X(net2561));
 sg13g2_buf_8 fanout2562 (.A(net2565),
    .X(net2562));
 sg13g2_buf_1 fanout2563 (.A(net2564),
    .X(net2563));
 sg13g2_buf_8 fanout2564 (.A(net2565),
    .X(net2564));
 sg13g2_buf_8 fanout2565 (.A(_01549_),
    .X(net2565));
 sg13g2_buf_8 fanout2566 (.A(net2567),
    .X(net2566));
 sg13g2_buf_2 fanout2567 (.A(_01417_),
    .X(net2567));
 sg13g2_buf_8 fanout2568 (.A(net3746),
    .X(net2568));
 sg13g2_buf_2 fanout2569 (.A(net2570),
    .X(net2569));
 sg13g2_buf_1 fanout2570 (.A(net2571),
    .X(net2570));
 sg13g2_buf_2 fanout2571 (.A(\cpu.cpu.decode.co_mem_word ),
    .X(net2571));
 sg13g2_buf_8 fanout2572 (.A(net2573),
    .X(net2572));
 sg13g2_buf_8 fanout2573 (.A(net2574),
    .X(net2573));
 sg13g2_buf_8 fanout2574 (.A(net3737),
    .X(net2574));
 sg13g2_buf_8 fanout2575 (.A(net2576),
    .X(net2575));
 sg13g2_buf_8 fanout2576 (.A(net3590),
    .X(net2576));
 sg13g2_buf_8 fanout2577 (.A(net3736),
    .X(net2577));
 sg13g2_buf_2 fanout2578 (.A(\cpu.cpu.decode.opcode[2] ),
    .X(net2578));
 sg13g2_buf_2 fanout2579 (.A(net2580),
    .X(net2579));
 sg13g2_buf_8 fanout2580 (.A(\cpu.cpu.decode.opcode[0] ),
    .X(net2580));
 sg13g2_buf_8 fanout2581 (.A(net2583),
    .X(net2581));
 sg13g2_buf_1 fanout2582 (.A(net2583),
    .X(net2582));
 sg13g2_buf_8 fanout2583 (.A(net1416),
    .X(net2583));
 sg13g2_buf_8 fanout2584 (.A(net2587),
    .X(net2584));
 sg13g2_buf_8 fanout2585 (.A(net2587),
    .X(net2585));
 sg13g2_buf_8 fanout2586 (.A(net2587),
    .X(net2586));
 sg13g2_buf_8 fanout2587 (.A(net1416),
    .X(net2587));
 sg13g2_buf_8 fanout2588 (.A(net2593),
    .X(net2588));
 sg13g2_buf_8 fanout2589 (.A(net2592),
    .X(net2589));
 sg13g2_buf_8 fanout2590 (.A(net2592),
    .X(net2590));
 sg13g2_buf_2 fanout2591 (.A(net2592),
    .X(net2591));
 sg13g2_buf_8 fanout2592 (.A(net2593),
    .X(net2592));
 sg13g2_buf_8 fanout2593 (.A(\cpu.rf_ram_if.gen_wtrig_ratio_neq_2.wtrig0_r ),
    .X(net2593));
 sg13g2_buf_8 fanout2594 (.A(net3726),
    .X(net2594));
 sg13g2_buf_8 fanout2595 (.A(net2596),
    .X(net2595));
 sg13g2_buf_8 fanout2596 (.A(net3731),
    .X(net2596));
 sg13g2_buf_8 fanout2597 (.A(net2598),
    .X(net2597));
 sg13g2_buf_1 fanout2598 (.A(net2601),
    .X(net2598));
 sg13g2_buf_8 fanout2599 (.A(net2601),
    .X(net2599));
 sg13g2_buf_1 fanout2600 (.A(net2601),
    .X(net2600));
 sg13g2_buf_8 fanout2601 (.A(net1),
    .X(net2601));
 sg13g2_buf_8 fanout2602 (.A(net1),
    .X(net2602));
 sg13g2_buf_2 input1 (.A(rst_n),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[4]),
    .X(net2));
 sg13g2_buf_1 input3 (.A(ui_in[5]),
    .X(net3));
 sg13g2_buf_1 input4 (.A(ui_in[6]),
    .X(net4));
 sg13g2_buf_1 input5 (.A(ui_in[7]),
    .X(net5));
 sg13g2_buf_1 input6 (.A(uio_in[2]),
    .X(net6));
 sg13g2_tielo tt_um_ECM24_serv_soc_top_7 (.L_LO(net7));
 sg13g2_buf_8 clkbuf_0_clk (.A(clk),
    .X(delaynet_0_clk));
 sg13g2_buf_8 clkbuf_1_0__f_clk (.A(clknet_0_clk),
    .X(clknet_1_0__leaf_clk));
 sg13g2_buf_8 clkbuf_1_1__f_clk (.A(clknet_0_clk),
    .X(clknet_1_1__leaf_clk));
 sg13g2_buf_1 clkload0 (.A(clknet_1_0__leaf_clk));
 sg13g2_buf_8 clkbuf_leaf_0_clk_regs (.A(clknet_5_0__leaf_clk_regs),
    .X(clknet_leaf_0_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_1_clk_regs (.A(clknet_5_0__leaf_clk_regs),
    .X(clknet_leaf_1_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_2_clk_regs (.A(clknet_5_0__leaf_clk_regs),
    .X(clknet_leaf_2_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_3_clk_regs (.A(clknet_5_0__leaf_clk_regs),
    .X(clknet_leaf_3_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_4_clk_regs (.A(clknet_5_1__leaf_clk_regs),
    .X(clknet_leaf_4_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_5_clk_regs (.A(clknet_5_3__leaf_clk_regs),
    .X(clknet_leaf_5_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_6_clk_regs (.A(clknet_5_2__leaf_clk_regs),
    .X(clknet_leaf_6_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_7_clk_regs (.A(clknet_5_2__leaf_clk_regs),
    .X(clknet_leaf_7_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_8_clk_regs (.A(clknet_5_2__leaf_clk_regs),
    .X(clknet_leaf_8_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_9_clk_regs (.A(clknet_5_2__leaf_clk_regs),
    .X(clknet_leaf_9_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_10_clk_regs (.A(clknet_5_2__leaf_clk_regs),
    .X(clknet_leaf_10_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_11_clk_regs (.A(clknet_5_2__leaf_clk_regs),
    .X(clknet_leaf_11_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_12_clk_regs (.A(clknet_5_3__leaf_clk_regs),
    .X(clknet_leaf_12_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_13_clk_regs (.A(clknet_5_3__leaf_clk_regs),
    .X(clknet_leaf_13_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_14_clk_regs (.A(clknet_5_3__leaf_clk_regs),
    .X(clknet_leaf_14_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_15_clk_regs (.A(clknet_5_3__leaf_clk_regs),
    .X(clknet_leaf_15_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_16_clk_regs (.A(clknet_5_6__leaf_clk_regs),
    .X(clknet_leaf_16_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_17_clk_regs (.A(clknet_5_6__leaf_clk_regs),
    .X(clknet_leaf_17_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_18_clk_regs (.A(clknet_5_12__leaf_clk_regs),
    .X(clknet_leaf_18_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_19_clk_regs (.A(clknet_5_6__leaf_clk_regs),
    .X(clknet_leaf_19_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_20_clk_regs (.A(clknet_5_6__leaf_clk_regs),
    .X(clknet_leaf_20_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_21_clk_regs (.A(clknet_5_13__leaf_clk_regs),
    .X(clknet_leaf_21_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_22_clk_regs (.A(clknet_5_12__leaf_clk_regs),
    .X(clknet_leaf_22_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_23_clk_regs (.A(clknet_5_12__leaf_clk_regs),
    .X(clknet_leaf_23_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_24_clk_regs (.A(clknet_5_12__leaf_clk_regs),
    .X(clknet_leaf_24_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_25_clk_regs (.A(clknet_5_12__leaf_clk_regs),
    .X(clknet_leaf_25_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_26_clk_regs (.A(clknet_5_9__leaf_clk_regs),
    .X(clknet_leaf_26_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_27_clk_regs (.A(clknet_5_9__leaf_clk_regs),
    .X(clknet_leaf_27_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_28_clk_regs (.A(clknet_5_9__leaf_clk_regs),
    .X(clknet_leaf_28_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_29_clk_regs (.A(clknet_5_9__leaf_clk_regs),
    .X(clknet_leaf_29_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_30_clk_regs (.A(clknet_5_8__leaf_clk_regs),
    .X(clknet_leaf_30_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_31_clk_regs (.A(clknet_5_8__leaf_clk_regs),
    .X(clknet_leaf_31_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_32_clk_regs (.A(clknet_5_8__leaf_clk_regs),
    .X(clknet_leaf_32_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_33_clk_regs (.A(clknet_5_8__leaf_clk_regs),
    .X(clknet_leaf_33_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_34_clk_regs (.A(clknet_5_8__leaf_clk_regs),
    .X(clknet_leaf_34_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_35_clk_regs (.A(clknet_5_9__leaf_clk_regs),
    .X(clknet_leaf_35_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_36_clk_regs (.A(clknet_5_10__leaf_clk_regs),
    .X(clknet_leaf_36_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_37_clk_regs (.A(clknet_5_8__leaf_clk_regs),
    .X(clknet_leaf_37_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_38_clk_regs (.A(clknet_5_10__leaf_clk_regs),
    .X(clknet_leaf_38_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_39_clk_regs (.A(clknet_5_10__leaf_clk_regs),
    .X(clknet_leaf_39_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_40_clk_regs (.A(clknet_5_10__leaf_clk_regs),
    .X(clknet_leaf_40_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_41_clk_regs (.A(clknet_5_10__leaf_clk_regs),
    .X(clknet_leaf_41_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_42_clk_regs (.A(clknet_5_10__leaf_clk_regs),
    .X(clknet_leaf_42_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_43_clk_regs (.A(clknet_5_11__leaf_clk_regs),
    .X(clknet_leaf_43_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_44_clk_regs (.A(clknet_5_11__leaf_clk_regs),
    .X(clknet_leaf_44_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_45_clk_regs (.A(clknet_5_11__leaf_clk_regs),
    .X(clknet_leaf_45_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_46_clk_regs (.A(clknet_5_11__leaf_clk_regs),
    .X(clknet_leaf_46_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_47_clk_regs (.A(clknet_5_14__leaf_clk_regs),
    .X(clknet_leaf_47_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_48_clk_regs (.A(clknet_5_11__leaf_clk_regs),
    .X(clknet_leaf_48_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_49_clk_regs (.A(clknet_5_14__leaf_clk_regs),
    .X(clknet_leaf_49_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_50_clk_regs (.A(clknet_5_14__leaf_clk_regs),
    .X(clknet_leaf_50_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_51_clk_regs (.A(clknet_5_15__leaf_clk_regs),
    .X(clknet_leaf_51_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_52_clk_regs (.A(clknet_5_15__leaf_clk_regs),
    .X(clknet_leaf_52_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_53_clk_regs (.A(clknet_5_15__leaf_clk_regs),
    .X(clknet_leaf_53_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_54_clk_regs (.A(clknet_5_15__leaf_clk_regs),
    .X(clknet_leaf_54_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_55_clk_regs (.A(clknet_5_15__leaf_clk_regs),
    .X(clknet_leaf_55_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_56_clk_regs (.A(clknet_5_14__leaf_clk_regs),
    .X(clknet_leaf_56_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_57_clk_regs (.A(clknet_5_14__leaf_clk_regs),
    .X(clknet_leaf_57_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_58_clk_regs (.A(clknet_5_12__leaf_clk_regs),
    .X(clknet_leaf_58_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_59_clk_regs (.A(clknet_5_13__leaf_clk_regs),
    .X(clknet_leaf_59_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_60_clk_regs (.A(clknet_5_13__leaf_clk_regs),
    .X(clknet_leaf_60_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_61_clk_regs (.A(clknet_5_13__leaf_clk_regs),
    .X(clknet_leaf_61_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_62_clk_regs (.A(clknet_5_13__leaf_clk_regs),
    .X(clknet_leaf_62_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_63_clk_regs (.A(clknet_5_24__leaf_clk_regs),
    .X(clknet_leaf_63_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_64_clk_regs (.A(clknet_5_24__leaf_clk_regs),
    .X(clknet_leaf_64_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_65_clk_regs (.A(clknet_5_24__leaf_clk_regs),
    .X(clknet_leaf_65_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_66_clk_regs (.A(clknet_5_24__leaf_clk_regs),
    .X(clknet_leaf_66_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_67_clk_regs (.A(clknet_5_24__leaf_clk_regs),
    .X(clknet_leaf_67_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_68_clk_regs (.A(clknet_5_25__leaf_clk_regs),
    .X(clknet_leaf_68_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_69_clk_regs (.A(clknet_5_26__leaf_clk_regs),
    .X(clknet_leaf_69_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_70_clk_regs (.A(clknet_5_26__leaf_clk_regs),
    .X(clknet_leaf_70_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_71_clk_regs (.A(clknet_5_26__leaf_clk_regs),
    .X(clknet_leaf_71_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_72_clk_regs (.A(clknet_5_26__leaf_clk_regs),
    .X(clknet_leaf_72_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_73_clk_regs (.A(clknet_5_26__leaf_clk_regs),
    .X(clknet_leaf_73_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_74_clk_regs (.A(clknet_5_26__leaf_clk_regs),
    .X(clknet_leaf_74_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_75_clk_regs (.A(clknet_5_27__leaf_clk_regs),
    .X(clknet_leaf_75_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_76_clk_regs (.A(clknet_5_27__leaf_clk_regs),
    .X(clknet_leaf_76_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_77_clk_regs (.A(clknet_5_27__leaf_clk_regs),
    .X(clknet_leaf_77_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_78_clk_regs (.A(clknet_5_27__leaf_clk_regs),
    .X(clknet_leaf_78_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_79_clk_regs (.A(clknet_5_27__leaf_clk_regs),
    .X(clknet_leaf_79_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_80_clk_regs (.A(clknet_5_30__leaf_clk_regs),
    .X(clknet_leaf_80_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_81_clk_regs (.A(clknet_5_30__leaf_clk_regs),
    .X(clknet_leaf_81_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_82_clk_regs (.A(clknet_5_30__leaf_clk_regs),
    .X(clknet_leaf_82_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_83_clk_regs (.A(clknet_5_30__leaf_clk_regs),
    .X(clknet_leaf_83_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_84_clk_regs (.A(clknet_5_31__leaf_clk_regs),
    .X(clknet_leaf_84_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_85_clk_regs (.A(clknet_5_31__leaf_clk_regs),
    .X(clknet_leaf_85_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_86_clk_regs (.A(clknet_5_31__leaf_clk_regs),
    .X(clknet_leaf_86_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_87_clk_regs (.A(clknet_5_31__leaf_clk_regs),
    .X(clknet_leaf_87_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_88_clk_regs (.A(clknet_5_31__leaf_clk_regs),
    .X(clknet_leaf_88_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_89_clk_regs (.A(clknet_5_30__leaf_clk_regs),
    .X(clknet_leaf_89_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_90_clk_regs (.A(clknet_5_28__leaf_clk_regs),
    .X(clknet_leaf_90_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_91_clk_regs (.A(clknet_5_28__leaf_clk_regs),
    .X(clknet_leaf_91_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_92_clk_regs (.A(clknet_5_29__leaf_clk_regs),
    .X(clknet_leaf_92_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_93_clk_regs (.A(clknet_5_29__leaf_clk_regs),
    .X(clknet_leaf_93_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_94_clk_regs (.A(clknet_5_29__leaf_clk_regs),
    .X(clknet_leaf_94_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_95_clk_regs (.A(clknet_5_29__leaf_clk_regs),
    .X(clknet_leaf_95_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_96_clk_regs (.A(clknet_5_29__leaf_clk_regs),
    .X(clknet_leaf_96_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_97_clk_regs (.A(clknet_5_28__leaf_clk_regs),
    .X(clknet_leaf_97_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_98_clk_regs (.A(clknet_5_28__leaf_clk_regs),
    .X(clknet_leaf_98_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_99_clk_regs (.A(clknet_5_28__leaf_clk_regs),
    .X(clknet_leaf_99_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_100_clk_regs (.A(clknet_5_28__leaf_clk_regs),
    .X(clknet_leaf_100_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_101_clk_regs (.A(clknet_5_25__leaf_clk_regs),
    .X(clknet_leaf_101_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_102_clk_regs (.A(clknet_5_25__leaf_clk_regs),
    .X(clknet_leaf_102_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_103_clk_regs (.A(clknet_5_25__leaf_clk_regs),
    .X(clknet_leaf_103_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_104_clk_regs (.A(clknet_5_25__leaf_clk_regs),
    .X(clknet_leaf_104_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_105_clk_regs (.A(clknet_5_24__leaf_clk_regs),
    .X(clknet_leaf_105_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_107_clk_regs (.A(clknet_5_19__leaf_clk_regs),
    .X(clknet_leaf_107_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_108_clk_regs (.A(clknet_5_19__leaf_clk_regs),
    .X(clknet_leaf_108_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_109_clk_regs (.A(clknet_5_19__leaf_clk_regs),
    .X(clknet_leaf_109_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_110_clk_regs (.A(clknet_5_19__leaf_clk_regs),
    .X(clknet_leaf_110_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_111_clk_regs (.A(clknet_5_22__leaf_clk_regs),
    .X(clknet_leaf_111_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_112_clk_regs (.A(clknet_5_22__leaf_clk_regs),
    .X(clknet_leaf_112_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_113_clk_regs (.A(clknet_5_22__leaf_clk_regs),
    .X(clknet_leaf_113_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_114_clk_regs (.A(clknet_5_22__leaf_clk_regs),
    .X(clknet_leaf_114_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_115_clk_regs (.A(clknet_5_23__leaf_clk_regs),
    .X(clknet_leaf_115_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_116_clk_regs (.A(clknet_5_23__leaf_clk_regs),
    .X(clknet_leaf_116_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_117_clk_regs (.A(clknet_5_23__leaf_clk_regs),
    .X(clknet_leaf_117_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_118_clk_regs (.A(clknet_5_23__leaf_clk_regs),
    .X(clknet_leaf_118_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_119_clk_regs (.A(clknet_5_23__leaf_clk_regs),
    .X(clknet_leaf_119_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_120_clk_regs (.A(clknet_5_22__leaf_clk_regs),
    .X(clknet_leaf_120_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_121_clk_regs (.A(clknet_5_20__leaf_clk_regs),
    .X(clknet_leaf_121_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_122_clk_regs (.A(clknet_5_20__leaf_clk_regs),
    .X(clknet_leaf_122_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_123_clk_regs (.A(clknet_5_21__leaf_clk_regs),
    .X(clknet_leaf_123_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_124_clk_regs (.A(clknet_5_21__leaf_clk_regs),
    .X(clknet_leaf_124_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_125_clk_regs (.A(clknet_5_21__leaf_clk_regs),
    .X(clknet_leaf_125_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_126_clk_regs (.A(clknet_5_21__leaf_clk_regs),
    .X(clknet_leaf_126_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_127_clk_regs (.A(clknet_5_21__leaf_clk_regs),
    .X(clknet_leaf_127_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_128_clk_regs (.A(clknet_5_20__leaf_clk_regs),
    .X(clknet_leaf_128_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_129_clk_regs (.A(clknet_5_20__leaf_clk_regs),
    .X(clknet_leaf_129_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_130_clk_regs (.A(clknet_5_20__leaf_clk_regs),
    .X(clknet_leaf_130_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_131_clk_regs (.A(clknet_5_20__leaf_clk_regs),
    .X(clknet_leaf_131_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_132_clk_regs (.A(clknet_5_17__leaf_clk_regs),
    .X(clknet_leaf_132_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_133_clk_regs (.A(clknet_5_17__leaf_clk_regs),
    .X(clknet_leaf_133_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_134_clk_regs (.A(clknet_5_17__leaf_clk_regs),
    .X(clknet_leaf_134_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_135_clk_regs (.A(clknet_5_17__leaf_clk_regs),
    .X(clknet_leaf_135_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_136_clk_regs (.A(clknet_5_16__leaf_clk_regs),
    .X(clknet_leaf_136_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_137_clk_regs (.A(clknet_5_16__leaf_clk_regs),
    .X(clknet_leaf_137_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_138_clk_regs (.A(clknet_5_16__leaf_clk_regs),
    .X(clknet_leaf_138_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_139_clk_regs (.A(clknet_5_16__leaf_clk_regs),
    .X(clknet_leaf_139_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_140_clk_regs (.A(clknet_5_16__leaf_clk_regs),
    .X(clknet_leaf_140_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_141_clk_regs (.A(clknet_5_16__leaf_clk_regs),
    .X(clknet_leaf_141_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_142_clk_regs (.A(clknet_5_18__leaf_clk_regs),
    .X(clknet_leaf_142_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_143_clk_regs (.A(clknet_5_17__leaf_clk_regs),
    .X(clknet_leaf_143_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_144_clk_regs (.A(clknet_5_19__leaf_clk_regs),
    .X(clknet_leaf_144_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_145_clk_regs (.A(clknet_5_18__leaf_clk_regs),
    .X(clknet_leaf_145_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_146_clk_regs (.A(clknet_5_18__leaf_clk_regs),
    .X(clknet_leaf_146_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_147_clk_regs (.A(clknet_5_18__leaf_clk_regs),
    .X(clknet_leaf_147_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_148_clk_regs (.A(clknet_5_18__leaf_clk_regs),
    .X(clknet_leaf_148_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_149_clk_regs (.A(clknet_5_7__leaf_clk_regs),
    .X(clknet_leaf_149_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_150_clk_regs (.A(clknet_5_7__leaf_clk_regs),
    .X(clknet_leaf_150_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_151_clk_regs (.A(clknet_5_7__leaf_clk_regs),
    .X(clknet_leaf_151_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_152_clk_regs (.A(clknet_5_7__leaf_clk_regs),
    .X(clknet_leaf_152_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_153_clk_regs (.A(clknet_5_6__leaf_clk_regs),
    .X(clknet_leaf_153_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_154_clk_regs (.A(clknet_5_6__leaf_clk_regs),
    .X(clknet_leaf_154_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_155_clk_regs (.A(clknet_5_4__leaf_clk_regs),
    .X(clknet_leaf_155_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_156_clk_regs (.A(clknet_5_7__leaf_clk_regs),
    .X(clknet_leaf_156_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_157_clk_regs (.A(clknet_5_5__leaf_clk_regs),
    .X(clknet_leaf_157_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_158_clk_regs (.A(clknet_5_5__leaf_clk_regs),
    .X(clknet_leaf_158_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_159_clk_regs (.A(clknet_5_5__leaf_clk_regs),
    .X(clknet_leaf_159_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_160_clk_regs (.A(clknet_5_5__leaf_clk_regs),
    .X(clknet_leaf_160_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_161_clk_regs (.A(clknet_5_5__leaf_clk_regs),
    .X(clknet_leaf_161_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_162_clk_regs (.A(clknet_5_4__leaf_clk_regs),
    .X(clknet_leaf_162_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_163_clk_regs (.A(clknet_5_4__leaf_clk_regs),
    .X(clknet_leaf_163_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_164_clk_regs (.A(clknet_5_4__leaf_clk_regs),
    .X(clknet_leaf_164_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_165_clk_regs (.A(clknet_5_4__leaf_clk_regs),
    .X(clknet_leaf_165_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_166_clk_regs (.A(clknet_5_1__leaf_clk_regs),
    .X(clknet_leaf_166_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_167_clk_regs (.A(clknet_5_1__leaf_clk_regs),
    .X(clknet_leaf_167_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_168_clk_regs (.A(clknet_5_4__leaf_clk_regs),
    .X(clknet_leaf_168_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_169_clk_regs (.A(clknet_5_1__leaf_clk_regs),
    .X(clknet_leaf_169_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_170_clk_regs (.A(clknet_5_1__leaf_clk_regs),
    .X(clknet_leaf_170_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_171_clk_regs (.A(clknet_5_0__leaf_clk_regs),
    .X(clknet_leaf_171_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_172_clk_regs (.A(clknet_5_0__leaf_clk_regs),
    .X(clknet_leaf_172_clk_regs));
 sg13g2_buf_8 clkbuf_0_clk_regs (.A(clk_regs),
    .X(clknet_0_clk_regs));
 sg13g2_buf_8 clkbuf_4_0_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_0_0_clk_regs));
 sg13g2_buf_8 clkbuf_4_1_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_1_0_clk_regs));
 sg13g2_buf_8 clkbuf_4_2_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_2_0_clk_regs));
 sg13g2_buf_8 clkbuf_4_3_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_3_0_clk_regs));
 sg13g2_buf_8 clkbuf_4_4_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_4_0_clk_regs));
 sg13g2_buf_8 clkbuf_4_5_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_5_0_clk_regs));
 sg13g2_buf_8 clkbuf_4_6_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_6_0_clk_regs));
 sg13g2_buf_8 clkbuf_4_7_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_7_0_clk_regs));
 sg13g2_buf_8 clkbuf_4_8_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_8_0_clk_regs));
 sg13g2_buf_8 clkbuf_4_9_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_9_0_clk_regs));
 sg13g2_buf_8 clkbuf_4_10_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_10_0_clk_regs));
 sg13g2_buf_8 clkbuf_4_11_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_11_0_clk_regs));
 sg13g2_buf_8 clkbuf_4_12_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_12_0_clk_regs));
 sg13g2_buf_8 clkbuf_4_13_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_13_0_clk_regs));
 sg13g2_buf_8 clkbuf_4_14_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_14_0_clk_regs));
 sg13g2_buf_8 clkbuf_4_15_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_15_0_clk_regs));
 sg13g2_buf_8 clkbuf_5_0__f_clk_regs (.A(clknet_4_0_0_clk_regs),
    .X(clknet_5_0__leaf_clk_regs));
 sg13g2_buf_8 clkbuf_5_1__f_clk_regs (.A(clknet_4_0_0_clk_regs),
    .X(clknet_5_1__leaf_clk_regs));
 sg13g2_buf_8 clkbuf_5_2__f_clk_regs (.A(clknet_4_1_0_clk_regs),
    .X(clknet_5_2__leaf_clk_regs));
 sg13g2_buf_8 clkbuf_5_3__f_clk_regs (.A(clknet_4_1_0_clk_regs),
    .X(clknet_5_3__leaf_clk_regs));
 sg13g2_buf_8 clkbuf_5_4__f_clk_regs (.A(clknet_4_2_0_clk_regs),
    .X(clknet_5_4__leaf_clk_regs));
 sg13g2_buf_8 clkbuf_5_5__f_clk_regs (.A(clknet_4_2_0_clk_regs),
    .X(clknet_5_5__leaf_clk_regs));
 sg13g2_buf_8 clkbuf_5_6__f_clk_regs (.A(clknet_4_3_0_clk_regs),
    .X(clknet_5_6__leaf_clk_regs));
 sg13g2_buf_8 clkbuf_5_7__f_clk_regs (.A(clknet_4_3_0_clk_regs),
    .X(clknet_5_7__leaf_clk_regs));
 sg13g2_buf_8 clkbuf_5_8__f_clk_regs (.A(clknet_4_4_0_clk_regs),
    .X(clknet_5_8__leaf_clk_regs));
 sg13g2_buf_8 clkbuf_5_9__f_clk_regs (.A(clknet_4_4_0_clk_regs),
    .X(clknet_5_9__leaf_clk_regs));
 sg13g2_buf_8 clkbuf_5_10__f_clk_regs (.A(clknet_4_5_0_clk_regs),
    .X(clknet_5_10__leaf_clk_regs));
 sg13g2_buf_8 clkbuf_5_11__f_clk_regs (.A(clknet_4_5_0_clk_regs),
    .X(clknet_5_11__leaf_clk_regs));
 sg13g2_buf_8 clkbuf_5_12__f_clk_regs (.A(clknet_4_6_0_clk_regs),
    .X(clknet_5_12__leaf_clk_regs));
 sg13g2_buf_8 clkbuf_5_13__f_clk_regs (.A(clknet_4_6_0_clk_regs),
    .X(clknet_5_13__leaf_clk_regs));
 sg13g2_buf_8 clkbuf_5_14__f_clk_regs (.A(clknet_4_7_0_clk_regs),
    .X(clknet_5_14__leaf_clk_regs));
 sg13g2_buf_8 clkbuf_5_15__f_clk_regs (.A(clknet_4_7_0_clk_regs),
    .X(clknet_5_15__leaf_clk_regs));
 sg13g2_buf_8 clkbuf_5_16__f_clk_regs (.A(clknet_4_8_0_clk_regs),
    .X(clknet_5_16__leaf_clk_regs));
 sg13g2_buf_8 clkbuf_5_17__f_clk_regs (.A(clknet_4_8_0_clk_regs),
    .X(clknet_5_17__leaf_clk_regs));
 sg13g2_buf_8 clkbuf_5_18__f_clk_regs (.A(clknet_4_9_0_clk_regs),
    .X(clknet_5_18__leaf_clk_regs));
 sg13g2_buf_8 clkbuf_5_19__f_clk_regs (.A(clknet_4_9_0_clk_regs),
    .X(clknet_5_19__leaf_clk_regs));
 sg13g2_buf_8 clkbuf_5_20__f_clk_regs (.A(clknet_4_10_0_clk_regs),
    .X(clknet_5_20__leaf_clk_regs));
 sg13g2_buf_8 clkbuf_5_21__f_clk_regs (.A(clknet_4_10_0_clk_regs),
    .X(clknet_5_21__leaf_clk_regs));
 sg13g2_buf_8 clkbuf_5_22__f_clk_regs (.A(clknet_4_11_0_clk_regs),
    .X(clknet_5_22__leaf_clk_regs));
 sg13g2_buf_8 clkbuf_5_23__f_clk_regs (.A(clknet_4_11_0_clk_regs),
    .X(clknet_5_23__leaf_clk_regs));
 sg13g2_buf_8 clkbuf_5_24__f_clk_regs (.A(clknet_4_12_0_clk_regs),
    .X(clknet_5_24__leaf_clk_regs));
 sg13g2_buf_8 clkbuf_5_25__f_clk_regs (.A(clknet_4_12_0_clk_regs),
    .X(clknet_5_25__leaf_clk_regs));
 sg13g2_buf_8 clkbuf_5_26__f_clk_regs (.A(clknet_4_13_0_clk_regs),
    .X(clknet_5_26__leaf_clk_regs));
 sg13g2_buf_8 clkbuf_5_27__f_clk_regs (.A(clknet_4_13_0_clk_regs),
    .X(clknet_5_27__leaf_clk_regs));
 sg13g2_buf_8 clkbuf_5_28__f_clk_regs (.A(clknet_4_14_0_clk_regs),
    .X(clknet_5_28__leaf_clk_regs));
 sg13g2_buf_8 clkbuf_5_29__f_clk_regs (.A(clknet_4_14_0_clk_regs),
    .X(clknet_5_29__leaf_clk_regs));
 sg13g2_buf_8 clkbuf_5_30__f_clk_regs (.A(clknet_4_15_0_clk_regs),
    .X(clknet_5_30__leaf_clk_regs));
 sg13g2_buf_8 clkbuf_5_31__f_clk_regs (.A(clknet_4_15_0_clk_regs),
    .X(clknet_5_31__leaf_clk_regs));
 sg13g2_buf_8 clkload1 (.A(clknet_5_1__leaf_clk_regs));
 sg13g2_buf_8 clkload2 (.A(clknet_5_3__leaf_clk_regs));
 sg13g2_buf_8 clkload3 (.A(clknet_5_5__leaf_clk_regs));
 sg13g2_buf_8 clkload4 (.A(clknet_5_7__leaf_clk_regs));
 sg13g2_buf_8 clkload5 (.A(clknet_5_9__leaf_clk_regs));
 sg13g2_buf_8 clkload6 (.A(clknet_5_11__leaf_clk_regs));
 sg13g2_buf_8 clkload7 (.A(clknet_5_13__leaf_clk_regs));
 sg13g2_buf_8 clkload8 (.A(clknet_5_17__leaf_clk_regs));
 sg13g2_inv_1 clkload9 (.A(clknet_5_19__leaf_clk_regs));
 sg13g2_buf_8 clkload10 (.A(clknet_5_21__leaf_clk_regs));
 sg13g2_buf_8 clkload11 (.A(clknet_5_25__leaf_clk_regs));
 sg13g2_buf_8 clkload12 (.A(clknet_5_27__leaf_clk_regs));
 sg13g2_buf_8 clkload13 (.A(clknet_5_29__leaf_clk_regs));
 sg13g2_inv_1 clkload14 (.A(clknet_leaf_172_clk_regs));
 sg13g2_inv_1 clkload15 (.A(clknet_leaf_11_clk_regs));
 sg13g2_inv_1 clkload16 (.A(clknet_leaf_33_clk_regs));
 sg13g2_inv_1 clkload17 (.A(clknet_leaf_62_clk_regs));
 sg13g2_buf_8 clkload18 (.A(clknet_leaf_105_clk_regs));
 sg13g2_inv_4 clkload19 (.A(clknet_leaf_85_clk_regs));
 sg13g2_buf_8 delaybuf_0_clk (.A(delaynet_0_clk),
    .X(clknet_0_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(\cpu.rf_ram_if.wdata0_r[11] ),
    .X(net1381));
 sg13g2_dlygate4sd3_1 hold2 (.A(\cpu.rf_ram_if.wdata0_r[27] ),
    .X(net1382));
 sg13g2_dlygate4sd3_1 hold3 (.A(\cpu.rf_ram_if.wdata0_r[22] ),
    .X(net1383));
 sg13g2_dlygate4sd3_1 hold4 (.A(\cpu.rf_ram_if.wdata0_r[31] ),
    .X(net1384));
 sg13g2_dlygate4sd3_1 hold5 (.A(\cpu.rf_ram_if.wdata0_r[15] ),
    .X(net1385));
 sg13g2_dlygate4sd3_1 hold6 (.A(\cpu.rf_ram_if.wdata0_r[30] ),
    .X(net1386));
 sg13g2_dlygate4sd3_1 hold7 (.A(\cpu.rf_ram_if.wdata0_r[3] ),
    .X(net1387));
 sg13g2_dlygate4sd3_1 hold8 (.A(\cpu.rf_ram_if.wdata0_r[18] ),
    .X(net1388));
 sg13g2_dlygate4sd3_1 hold9 (.A(\cpu.rf_ram_if.wdata0_r[14] ),
    .X(net1389));
 sg13g2_dlygate4sd3_1 hold10 (.A(\cpu.rf_ram_if.wdata0_r[19] ),
    .X(net1390));
 sg13g2_dlygate4sd3_1 hold11 (.A(\cpu.rf_ram_if.wdata0_r[24] ),
    .X(net1391));
 sg13g2_dlygate4sd3_1 hold12 (.A(\cpu.rf_ram_if.wdata0_r[10] ),
    .X(net1392));
 sg13g2_dlygate4sd3_1 hold13 (.A(\cpu.rf_ram_if.wdata0_r[5] ),
    .X(net1393));
 sg13g2_dlygate4sd3_1 hold14 (.A(\cpu.rf_ram_if.wdata0_r[16] ),
    .X(net1394));
 sg13g2_dlygate4sd3_1 hold15 (.A(\cpu.rf_ram_if.wdata0_r[29] ),
    .X(net1395));
 sg13g2_dlygate4sd3_1 hold16 (.A(\cpu.rf_ram_if.wdata0_r[13] ),
    .X(net1396));
 sg13g2_dlygate4sd3_1 hold17 (.A(\cpu.rf_ram_if.wdata0_r[7] ),
    .X(net1397));
 sg13g2_dlygate4sd3_1 hold18 (.A(\cpu.rf_ram_if.wdata0_r[17] ),
    .X(net1398));
 sg13g2_dlygate4sd3_1 hold19 (.A(\cpu.rf_ram_if.wdata0_r[23] ),
    .X(net1399));
 sg13g2_dlygate4sd3_1 hold20 (.A(\cpu.rf_ram_if.wdata0_r[4] ),
    .X(net1400));
 sg13g2_dlygate4sd3_1 hold21 (.A(\cpu.rf_ram_if.wdata0_r[12] ),
    .X(net1401));
 sg13g2_dlygate4sd3_1 hold22 (.A(\cpu.rf_ram_if.wdata0_r[8] ),
    .X(net1402));
 sg13g2_dlygate4sd3_1 hold23 (.A(\cpu.rf_ram_if.wdata0_r[21] ),
    .X(net1403));
 sg13g2_dlygate4sd3_1 hold24 (.A(\cpu.rf_ram_if.rdata0[21] ),
    .X(net1404));
 sg13g2_dlygate4sd3_1 hold25 (.A(_00012_),
    .X(net1405));
 sg13g2_dlygate4sd3_1 hold26 (.A(\cpu.rf_ram_if.wdata0_r[28] ),
    .X(net1406));
 sg13g2_dlygate4sd3_1 hold27 (.A(\cpu.rf_ram_if.wdata0_r[25] ),
    .X(net1407));
 sg13g2_dlygate4sd3_1 hold28 (.A(\cpu.rf_ram_if.wdata0_r[6] ),
    .X(net1408));
 sg13g2_dlygate4sd3_1 hold29 (.A(\cpu.rf_ram_if.wdata0_r[9] ),
    .X(net1409));
 sg13g2_dlygate4sd3_1 hold30 (.A(\cpu.rf_ram_if.wdata0_r[1] ),
    .X(net1410));
 sg13g2_dlygate4sd3_1 hold31 (.A(\cpu.rf_ram_if.wdata0_r[26] ),
    .X(net1411));
 sg13g2_dlygate4sd3_1 hold32 (.A(\cpu.rf_ram_if.wdata0_r[2] ),
    .X(net1412));
 sg13g2_dlygate4sd3_1 hold33 (.A(\cpu.rf_ram_if.wdata0_r[20] ),
    .X(net1413));
 sg13g2_dlygate4sd3_1 hold34 (.A(\cpu.rf_ram_if.rreq_r ),
    .X(net1414));
 sg13g2_dlygate4sd3_1 hold35 (.A(\cpu.i_rf_rdata[31] ),
    .X(net1415));
 sg13g2_dlygate4sd3_1 hold36 (.A(\cpu.rf_ram_if.rtrig1 ),
    .X(net1416));
 sg13g2_dlygate4sd3_1 hold37 (.A(\ram_spi_if.cycle_counter[0] ),
    .X(net1417));
 sg13g2_dlygate4sd3_1 hold38 (.A(\rf_ram.RAM[10][1] ),
    .X(net1418));
 sg13g2_dlygate4sd3_1 hold39 (.A(\rf_ram.RAM[2][14] ),
    .X(net1419));
 sg13g2_dlygate4sd3_1 hold40 (.A(\rf_ram.RAM[8][12] ),
    .X(net1420));
 sg13g2_dlygate4sd3_1 hold41 (.A(\rf_ram.RAM[0][30] ),
    .X(net1421));
 sg13g2_dlygate4sd3_1 hold42 (.A(\rf_ram.RAM[14][9] ),
    .X(net1422));
 sg13g2_dlygate4sd3_1 hold43 (.A(\rf_ram.RAM[6][14] ),
    .X(net1423));
 sg13g2_dlygate4sd3_1 hold44 (.A(\rf_ram.RAM[28][7] ),
    .X(net1424));
 sg13g2_dlygate4sd3_1 hold45 (.A(\rf_ram.RAM[8][25] ),
    .X(net1425));
 sg13g2_dlygate4sd3_1 hold46 (.A(\rf_ram.RAM[26][14] ),
    .X(net1426));
 sg13g2_dlygate4sd3_1 hold47 (.A(\rf_ram.RAM[20][12] ),
    .X(net1427));
 sg13g2_dlygate4sd3_1 hold48 (.A(\rf_ram.RAM[4][4] ),
    .X(net1428));
 sg13g2_dlygate4sd3_1 hold49 (.A(\rf_ram.RAM[4][16] ),
    .X(net1429));
 sg13g2_dlygate4sd3_1 hold50 (.A(\rf_ram.RAM[22][6] ),
    .X(net1430));
 sg13g2_dlygate4sd3_1 hold51 (.A(\rf_ram.RAM[20][15] ),
    .X(net1431));
 sg13g2_dlygate4sd3_1 hold52 (.A(\rf_ram.RAM[28][19] ),
    .X(net1432));
 sg13g2_dlygate4sd3_1 hold53 (.A(\rf_ram.RAM[18][8] ),
    .X(net1433));
 sg13g2_dlygate4sd3_1 hold54 (.A(\rf_ram.RAM[2][19] ),
    .X(net1434));
 sg13g2_dlygate4sd3_1 hold55 (.A(\rf_ram.RAM[22][18] ),
    .X(net1435));
 sg13g2_dlygate4sd3_1 hold56 (.A(\rf_ram.RAM[18][14] ),
    .X(net1436));
 sg13g2_dlygate4sd3_1 hold57 (.A(\rf_ram.RAM[20][18] ),
    .X(net1437));
 sg13g2_dlygate4sd3_1 hold58 (.A(\rf_ram.RAM[12][29] ),
    .X(net1438));
 sg13g2_dlygate4sd3_1 hold59 (.A(\rf_ram.RAM[20][30] ),
    .X(net1439));
 sg13g2_dlygate4sd3_1 hold60 (.A(\rf_ram.RAM[31][19] ),
    .X(net1440));
 sg13g2_dlygate4sd3_1 hold61 (.A(\rf_ram.RAM[10][10] ),
    .X(net1441));
 sg13g2_dlygate4sd3_1 hold62 (.A(\rf_ram.RAM[25][26] ),
    .X(net1442));
 sg13g2_dlygate4sd3_1 hold63 (.A(\rf_ram.RAM[0][21] ),
    .X(net1443));
 sg13g2_dlygate4sd3_1 hold64 (.A(\rf_ram.RAM[0][17] ),
    .X(net1444));
 sg13g2_dlygate4sd3_1 hold65 (.A(\rf_ram.RAM[7][15] ),
    .X(net1445));
 sg13g2_dlygate4sd3_1 hold66 (.A(\rf_ram.RAM[4][0] ),
    .X(net1446));
 sg13g2_dlygate4sd3_1 hold67 (.A(_00652_),
    .X(net1447));
 sg13g2_dlygate4sd3_1 hold68 (.A(\rf_ram.RAM[27][29] ),
    .X(net1448));
 sg13g2_dlygate4sd3_1 hold69 (.A(\rf_ram.RAM[30][15] ),
    .X(net1449));
 sg13g2_dlygate4sd3_1 hold70 (.A(\rf_ram.RAM[4][19] ),
    .X(net1450));
 sg13g2_dlygate4sd3_1 hold71 (.A(\rf_ram.RAM[23][15] ),
    .X(net1451));
 sg13g2_dlygate4sd3_1 hold72 (.A(\rf_ram.RAM[13][17] ),
    .X(net1452));
 sg13g2_dlygate4sd3_1 hold73 (.A(\rf_ram.RAM[25][8] ),
    .X(net1453));
 sg13g2_dlygate4sd3_1 hold74 (.A(\rf_ram.RAM[18][11] ),
    .X(net1454));
 sg13g2_dlygate4sd3_1 hold75 (.A(\rf_ram.RAM[8][29] ),
    .X(net1455));
 sg13g2_dlygate4sd3_1 hold76 (.A(\rf_ram.RAM[8][14] ),
    .X(net1456));
 sg13g2_dlygate4sd3_1 hold77 (.A(\rf_ram.RAM[22][29] ),
    .X(net1457));
 sg13g2_dlygate4sd3_1 hold78 (.A(\rf_ram.RAM[24][23] ),
    .X(net1458));
 sg13g2_dlygate4sd3_1 hold79 (.A(\rf_ram.RAM[8][26] ),
    .X(net1459));
 sg13g2_dlygate4sd3_1 hold80 (.A(\rf_ram.RAM[15][17] ),
    .X(net1460));
 sg13g2_dlygate4sd3_1 hold81 (.A(\rf_ram.RAM[14][1] ),
    .X(net1461));
 sg13g2_dlygate4sd3_1 hold82 (.A(\rf_ram.RAM[18][10] ),
    .X(net1462));
 sg13g2_dlygate4sd3_1 hold83 (.A(\rf_ram.RAM[0][6] ),
    .X(net1463));
 sg13g2_dlygate4sd3_1 hold84 (.A(\rf_ram.RAM[2][25] ),
    .X(net1464));
 sg13g2_dlygate4sd3_1 hold85 (.A(\rf_ram.RAM[4][25] ),
    .X(net1465));
 sg13g2_dlygate4sd3_1 hold86 (.A(\rf_ram.RAM[28][29] ),
    .X(net1466));
 sg13g2_dlygate4sd3_1 hold87 (.A(\rf_ram.RAM[18][12] ),
    .X(net1467));
 sg13g2_dlygate4sd3_1 hold88 (.A(\rf_ram.RAM[3][10] ),
    .X(net1468));
 sg13g2_dlygate4sd3_1 hold89 (.A(\rf_ram.RAM[30][26] ),
    .X(net1469));
 sg13g2_dlygate4sd3_1 hold90 (.A(\rf_ram.RAM[20][31] ),
    .X(net1470));
 sg13g2_dlygate4sd3_1 hold91 (.A(\rf_ram.RAM[14][19] ),
    .X(net1471));
 sg13g2_dlygate4sd3_1 hold92 (.A(\rf_ram.RAM[20][9] ),
    .X(net1472));
 sg13g2_dlygate4sd3_1 hold93 (.A(\rf_ram.RAM[8][31] ),
    .X(net1473));
 sg13g2_dlygate4sd3_1 hold94 (.A(\rf_ram.RAM[27][12] ),
    .X(net1474));
 sg13g2_dlygate4sd3_1 hold95 (.A(\rf_ram.RAM[15][12] ),
    .X(net1475));
 sg13g2_dlygate4sd3_1 hold96 (.A(\rf_ram.RAM[14][22] ),
    .X(net1476));
 sg13g2_dlygate4sd3_1 hold97 (.A(\rf_ram.RAM[0][9] ),
    .X(net1477));
 sg13g2_dlygate4sd3_1 hold98 (.A(\rf_ram.RAM[0][31] ),
    .X(net1478));
 sg13g2_dlygate4sd3_1 hold99 (.A(\rf_ram.RAM[29][4] ),
    .X(net1479));
 sg13g2_dlygate4sd3_1 hold100 (.A(\rf_ram.RAM[5][4] ),
    .X(net1480));
 sg13g2_dlygate4sd3_1 hold101 (.A(\rf_ram.RAM[16][13] ),
    .X(net1481));
 sg13g2_dlygate4sd3_1 hold102 (.A(\rf_ram.RAM[0][4] ),
    .X(net1482));
 sg13g2_dlygate4sd3_1 hold103 (.A(\rf_ram.RAM[12][11] ),
    .X(net1483));
 sg13g2_dlygate4sd3_1 hold104 (.A(\rf_ram.RAM[30][8] ),
    .X(net1484));
 sg13g2_dlygate4sd3_1 hold105 (.A(\rf_ram.RAM[20][11] ),
    .X(net1485));
 sg13g2_dlygate4sd3_1 hold106 (.A(\rf_ram.RAM[8][11] ),
    .X(net1486));
 sg13g2_dlygate4sd3_1 hold107 (.A(\rf_ram.RAM[30][23] ),
    .X(net1487));
 sg13g2_dlygate4sd3_1 hold108 (.A(\rf_ram.RAM[20][8] ),
    .X(net1488));
 sg13g2_dlygate4sd3_1 hold109 (.A(\rf_ram.RAM[9][18] ),
    .X(net1489));
 sg13g2_dlygate4sd3_1 hold110 (.A(\rf_ram.RAM[10][9] ),
    .X(net1490));
 sg13g2_dlygate4sd3_1 hold111 (.A(\rf_ram.RAM[2][17] ),
    .X(net1491));
 sg13g2_dlygate4sd3_1 hold112 (.A(\rf_ram.RAM[29][11] ),
    .X(net1492));
 sg13g2_dlygate4sd3_1 hold113 (.A(\rf_ram.RAM[18][16] ),
    .X(net1493));
 sg13g2_dlygate4sd3_1 hold114 (.A(\rf_ram.RAM[26][4] ),
    .X(net1494));
 sg13g2_dlygate4sd3_1 hold115 (.A(\rf_ram.RAM[12][8] ),
    .X(net1495));
 sg13g2_dlygate4sd3_1 hold116 (.A(\rf_ram.RAM[2][27] ),
    .X(net1496));
 sg13g2_dlygate4sd3_1 hold117 (.A(\rf_ram.RAM[10][17] ),
    .X(net1497));
 sg13g2_dlygate4sd3_1 hold118 (.A(\rf_ram.RAM[9][9] ),
    .X(net1498));
 sg13g2_dlygate4sd3_1 hold119 (.A(\rf_ram.RAM[28][23] ),
    .X(net1499));
 sg13g2_dlygate4sd3_1 hold120 (.A(\rf_ram.RAM[26][18] ),
    .X(net1500));
 sg13g2_dlygate4sd3_1 hold121 (.A(\rf_ram.RAM[2][10] ),
    .X(net1501));
 sg13g2_dlygate4sd3_1 hold122 (.A(\rf_ram.RAM[3][7] ),
    .X(net1502));
 sg13g2_dlygate4sd3_1 hold123 (.A(\rf_ram.RAM[21][15] ),
    .X(net1503));
 sg13g2_dlygate4sd3_1 hold124 (.A(\rf_ram.RAM[30][6] ),
    .X(net1504));
 sg13g2_dlygate4sd3_1 hold125 (.A(\rf_ram.RAM[20][28] ),
    .X(net1505));
 sg13g2_dlygate4sd3_1 hold126 (.A(\rf_ram.RAM[11][6] ),
    .X(net1506));
 sg13g2_dlygate4sd3_1 hold127 (.A(\rf_ram.RAM[26][30] ),
    .X(net1507));
 sg13g2_dlygate4sd3_1 hold128 (.A(\rf_ram.RAM[22][19] ),
    .X(net1508));
 sg13g2_dlygate4sd3_1 hold129 (.A(\rf_ram.RAM[9][31] ),
    .X(net1509));
 sg13g2_dlygate4sd3_1 hold130 (.A(\rf_ram.RAM[30][17] ),
    .X(net1510));
 sg13g2_dlygate4sd3_1 hold131 (.A(\rf_ram.RAM[27][19] ),
    .X(net1511));
 sg13g2_dlygate4sd3_1 hold132 (.A(\rf_ram.RAM[6][18] ),
    .X(net1512));
 sg13g2_dlygate4sd3_1 hold133 (.A(\rf_ram.RAM[7][6] ),
    .X(net1513));
 sg13g2_dlygate4sd3_1 hold134 (.A(\rf_ram.RAM[16][18] ),
    .X(net1514));
 sg13g2_dlygate4sd3_1 hold135 (.A(\rf_ram.RAM[5][5] ),
    .X(net1515));
 sg13g2_dlygate4sd3_1 hold136 (.A(\rf_ram.RAM[2][13] ),
    .X(net1516));
 sg13g2_dlygate4sd3_1 hold137 (.A(\rf_ram.RAM[18][26] ),
    .X(net1517));
 sg13g2_dlygate4sd3_1 hold138 (.A(\rf_ram.RAM[13][9] ),
    .X(net1518));
 sg13g2_dlygate4sd3_1 hold139 (.A(\rf_ram.RAM[10][6] ),
    .X(net1519));
 sg13g2_dlygate4sd3_1 hold140 (.A(\rf_ram.RAM[16][26] ),
    .X(net1520));
 sg13g2_dlygate4sd3_1 hold141 (.A(\rf_ram.RAM[14][28] ),
    .X(net1521));
 sg13g2_dlygate4sd3_1 hold142 (.A(\rf_ram.RAM[20][4] ),
    .X(net1522));
 sg13g2_dlygate4sd3_1 hold143 (.A(\rf_ram.RAM[9][28] ),
    .X(net1523));
 sg13g2_dlygate4sd3_1 hold144 (.A(\rf_ram.RAM[17][19] ),
    .X(net1524));
 sg13g2_dlygate4sd3_1 hold145 (.A(\rf_ram.RAM[11][7] ),
    .X(net1525));
 sg13g2_dlygate4sd3_1 hold146 (.A(\rf_ram.RAM[20][19] ),
    .X(net1526));
 sg13g2_dlygate4sd3_1 hold147 (.A(\rf_ram.RAM[24][18] ),
    .X(net1527));
 sg13g2_dlygate4sd3_1 hold148 (.A(\rf_ram.RAM[26][12] ),
    .X(net1528));
 sg13g2_dlygate4sd3_1 hold149 (.A(\rf_ram.RAM[9][6] ),
    .X(net1529));
 sg13g2_dlygate4sd3_1 hold150 (.A(\rf_ram.RAM[16][15] ),
    .X(net1530));
 sg13g2_dlygate4sd3_1 hold151 (.A(\rf_ram.RAM[11][30] ),
    .X(net1531));
 sg13g2_dlygate4sd3_1 hold152 (.A(\rf_ram.RAM[1][30] ),
    .X(net1532));
 sg13g2_dlygate4sd3_1 hold153 (.A(\rf_ram.RAM[29][28] ),
    .X(net1533));
 sg13g2_dlygate4sd3_1 hold154 (.A(\rf_ram.RAM[12][14] ),
    .X(net1534));
 sg13g2_dlygate4sd3_1 hold155 (.A(\rf_ram.RAM[10][21] ),
    .X(net1535));
 sg13g2_dlygate4sd3_1 hold156 (.A(\rf_ram.RAM[10][25] ),
    .X(net1536));
 sg13g2_dlygate4sd3_1 hold157 (.A(\rf_ram.RAM[18][1] ),
    .X(net1537));
 sg13g2_dlygate4sd3_1 hold158 (.A(\rf_ram.RAM[10][28] ),
    .X(net1538));
 sg13g2_dlygate4sd3_1 hold159 (.A(\rf_ram.RAM[13][14] ),
    .X(net1539));
 sg13g2_dlygate4sd3_1 hold160 (.A(\rf_ram.RAM[16][9] ),
    .X(net1540));
 sg13g2_dlygate4sd3_1 hold161 (.A(\rf_ram.RAM[20][21] ),
    .X(net1541));
 sg13g2_dlygate4sd3_1 hold162 (.A(\rf_ram.RAM[26][1] ),
    .X(net1542));
 sg13g2_dlygate4sd3_1 hold163 (.A(\rf_ram.RAM[31][22] ),
    .X(net1543));
 sg13g2_dlygate4sd3_1 hold164 (.A(\rf_ram.RAM[22][25] ),
    .X(net1544));
 sg13g2_dlygate4sd3_1 hold165 (.A(\rf_ram.RAM[24][30] ),
    .X(net1545));
 sg13g2_dlygate4sd3_1 hold166 (.A(\rf_ram.RAM[9][5] ),
    .X(net1546));
 sg13g2_dlygate4sd3_1 hold167 (.A(\rf_ram.RAM[9][1] ),
    .X(net1547));
 sg13g2_dlygate4sd3_1 hold168 (.A(\rf_ram.RAM[9][24] ),
    .X(net1548));
 sg13g2_dlygate4sd3_1 hold169 (.A(\rf_ram.RAM[13][18] ),
    .X(net1549));
 sg13g2_dlygate4sd3_1 hold170 (.A(\rf_ram.RAM[0][10] ),
    .X(net1550));
 sg13g2_dlygate4sd3_1 hold171 (.A(\rf_ram.RAM[19][4] ),
    .X(net1551));
 sg13g2_dlygate4sd3_1 hold172 (.A(\rf_ram.RAM[25][9] ),
    .X(net1552));
 sg13g2_dlygate4sd3_1 hold173 (.A(\rf_ram.RAM[16][30] ),
    .X(net1553));
 sg13g2_dlygate4sd3_1 hold174 (.A(\rf_ram.RAM[14][20] ),
    .X(net1554));
 sg13g2_dlygate4sd3_1 hold175 (.A(\rf_ram.RAM[30][2] ),
    .X(net1555));
 sg13g2_dlygate4sd3_1 hold176 (.A(\rf_ram.RAM[0][24] ),
    .X(net1556));
 sg13g2_dlygate4sd3_1 hold177 (.A(\rf_ram.RAM[31][9] ),
    .X(net1557));
 sg13g2_dlygate4sd3_1 hold178 (.A(\rf_ram.RAM[19][23] ),
    .X(net1558));
 sg13g2_dlygate4sd3_1 hold179 (.A(\rf_ram.RAM[10][12] ),
    .X(net1559));
 sg13g2_dlygate4sd3_1 hold180 (.A(\rf_ram.RAM[5][10] ),
    .X(net1560));
 sg13g2_dlygate4sd3_1 hold181 (.A(\rf_ram.RAM[8][3] ),
    .X(net1561));
 sg13g2_dlygate4sd3_1 hold182 (.A(\rf_ram.RAM[17][7] ),
    .X(net1562));
 sg13g2_dlygate4sd3_1 hold183 (.A(\rf_ram.RAM[12][27] ),
    .X(net1563));
 sg13g2_dlygate4sd3_1 hold184 (.A(\rf_ram.RAM[3][13] ),
    .X(net1564));
 sg13g2_dlygate4sd3_1 hold185 (.A(\rf_ram.RAM[3][16] ),
    .X(net1565));
 sg13g2_dlygate4sd3_1 hold186 (.A(\rf_ram.RAM[0][19] ),
    .X(net1566));
 sg13g2_dlygate4sd3_1 hold187 (.A(\rf_ram.RAM[13][20] ),
    .X(net1567));
 sg13g2_dlygate4sd3_1 hold188 (.A(\rf_ram.RAM[26][21] ),
    .X(net1568));
 sg13g2_dlygate4sd3_1 hold189 (.A(\rf_ram.RAM[30][31] ),
    .X(net1569));
 sg13g2_dlygate4sd3_1 hold190 (.A(\rf_ram.RAM[11][1] ),
    .X(net1570));
 sg13g2_dlygate4sd3_1 hold191 (.A(\rf_ram.RAM[27][9] ),
    .X(net1571));
 sg13g2_dlygate4sd3_1 hold192 (.A(\rf_ram.RAM[2][0] ),
    .X(net1572));
 sg13g2_dlygate4sd3_1 hold193 (.A(_01028_),
    .X(net1573));
 sg13g2_dlygate4sd3_1 hold194 (.A(\rf_ram.RAM[19][27] ),
    .X(net1574));
 sg13g2_dlygate4sd3_1 hold195 (.A(\rf_ram.RAM[20][0] ),
    .X(net1575));
 sg13g2_dlygate4sd3_1 hold196 (.A(_00183_),
    .X(net1576));
 sg13g2_dlygate4sd3_1 hold197 (.A(\rf_ram.RAM[23][23] ),
    .X(net1577));
 sg13g2_dlygate4sd3_1 hold198 (.A(\rf_ram.RAM[7][14] ),
    .X(net1578));
 sg13g2_dlygate4sd3_1 hold199 (.A(\rf_ram.RAM[10][27] ),
    .X(net1579));
 sg13g2_dlygate4sd3_1 hold200 (.A(\rf_ram.RAM[11][19] ),
    .X(net1580));
 sg13g2_dlygate4sd3_1 hold201 (.A(\rf_ram.RAM[14][29] ),
    .X(net1581));
 sg13g2_dlygate4sd3_1 hold202 (.A(\rf_ram.RAM[13][30] ),
    .X(net1582));
 sg13g2_dlygate4sd3_1 hold203 (.A(\rf_ram.RAM[18][21] ),
    .X(net1583));
 sg13g2_dlygate4sd3_1 hold204 (.A(\rf_ram.RAM[17][26] ),
    .X(net1584));
 sg13g2_dlygate4sd3_1 hold205 (.A(\rf_ram.RAM[28][2] ),
    .X(net1585));
 sg13g2_dlygate4sd3_1 hold206 (.A(\rf_ram.RAM[13][29] ),
    .X(net1586));
 sg13g2_dlygate4sd3_1 hold207 (.A(\rf_ram.RAM[21][26] ),
    .X(net1587));
 sg13g2_dlygate4sd3_1 hold208 (.A(\rf_ram.RAM[14][15] ),
    .X(net1588));
 sg13g2_dlygate4sd3_1 hold209 (.A(\rf_ram.RAM[13][1] ),
    .X(net1589));
 sg13g2_dlygate4sd3_1 hold210 (.A(\rf_ram.RAM[25][30] ),
    .X(net1590));
 sg13g2_dlygate4sd3_1 hold211 (.A(\rf_ram.RAM[11][5] ),
    .X(net1591));
 sg13g2_dlygate4sd3_1 hold212 (.A(\rf_ram.RAM[9][20] ),
    .X(net1592));
 sg13g2_dlygate4sd3_1 hold213 (.A(\rf_ram.RAM[28][1] ),
    .X(net1593));
 sg13g2_dlygate4sd3_1 hold214 (.A(\rf_ram.RAM[25][31] ),
    .X(net1594));
 sg13g2_dlygate4sd3_1 hold215 (.A(\rf_ram.RAM[1][29] ),
    .X(net1595));
 sg13g2_dlygate4sd3_1 hold216 (.A(\rf_ram.RAM[26][26] ),
    .X(net1596));
 sg13g2_dlygate4sd3_1 hold217 (.A(\rf_ram.RAM[15][5] ),
    .X(net1597));
 sg13g2_dlygate4sd3_1 hold218 (.A(\rf_ram.RAM[19][22] ),
    .X(net1598));
 sg13g2_dlygate4sd3_1 hold219 (.A(\rf_ram.RAM[9][26] ),
    .X(net1599));
 sg13g2_dlygate4sd3_1 hold220 (.A(\rf_ram.RAM[10][4] ),
    .X(net1600));
 sg13g2_dlygate4sd3_1 hold221 (.A(\rf_ram.RAM[29][6] ),
    .X(net1601));
 sg13g2_dlygate4sd3_1 hold222 (.A(\rf_ram.RAM[8][20] ),
    .X(net1602));
 sg13g2_dlygate4sd3_1 hold223 (.A(\rf_ram.RAM[21][24] ),
    .X(net1603));
 sg13g2_dlygate4sd3_1 hold224 (.A(\rf_ram.RAM[6][22] ),
    .X(net1604));
 sg13g2_dlygate4sd3_1 hold225 (.A(\rf_ram.RAM[7][17] ),
    .X(net1605));
 sg13g2_dlygate4sd3_1 hold226 (.A(\rf_ram.RAM[0][23] ),
    .X(net1606));
 sg13g2_dlygate4sd3_1 hold227 (.A(\rf_ram.RAM[31][28] ),
    .X(net1607));
 sg13g2_dlygate4sd3_1 hold228 (.A(\rf_ram.RAM[29][23] ),
    .X(net1608));
 sg13g2_dlygate4sd3_1 hold229 (.A(\rf_ram.RAM[17][28] ),
    .X(net1609));
 sg13g2_dlygate4sd3_1 hold230 (.A(\rf_ram.RAM[29][18] ),
    .X(net1610));
 sg13g2_dlygate4sd3_1 hold231 (.A(\rf_ram.RAM[30][19] ),
    .X(net1611));
 sg13g2_dlygate4sd3_1 hold232 (.A(\rf_ram.RAM[2][8] ),
    .X(net1612));
 sg13g2_dlygate4sd3_1 hold233 (.A(\rf_ram.RAM[18][28] ),
    .X(net1613));
 sg13g2_dlygate4sd3_1 hold234 (.A(\rf_ram.RAM[3][21] ),
    .X(net1614));
 sg13g2_dlygate4sd3_1 hold235 (.A(\rf_ram.RAM[23][16] ),
    .X(net1615));
 sg13g2_dlygate4sd3_1 hold236 (.A(\rf_ram.RAM[5][20] ),
    .X(net1616));
 sg13g2_dlygate4sd3_1 hold237 (.A(\rf_ram.RAM[16][31] ),
    .X(net1617));
 sg13g2_dlygate4sd3_1 hold238 (.A(\rf_ram.RAM[6][15] ),
    .X(net1618));
 sg13g2_dlygate4sd3_1 hold239 (.A(\rf_ram.RAM[10][2] ),
    .X(net1619));
 sg13g2_dlygate4sd3_1 hold240 (.A(\rf_ram.RAM[29][15] ),
    .X(net1620));
 sg13g2_dlygate4sd3_1 hold241 (.A(\rf_ram.RAM[26][7] ),
    .X(net1621));
 sg13g2_dlygate4sd3_1 hold242 (.A(\rf_ram.RAM[10][30] ),
    .X(net1622));
 sg13g2_dlygate4sd3_1 hold243 (.A(\rf_ram.RAM[4][26] ),
    .X(net1623));
 sg13g2_dlygate4sd3_1 hold244 (.A(\rf_ram.RAM[13][15] ),
    .X(net1624));
 sg13g2_dlygate4sd3_1 hold245 (.A(\rf_ram.RAM[27][21] ),
    .X(net1625));
 sg13g2_dlygate4sd3_1 hold246 (.A(\rf_ram.RAM[1][25] ),
    .X(net1626));
 sg13g2_dlygate4sd3_1 hold247 (.A(\rf_ram.RAM[3][25] ),
    .X(net1627));
 sg13g2_dlygate4sd3_1 hold248 (.A(\rf_ram.RAM[26][28] ),
    .X(net1628));
 sg13g2_dlygate4sd3_1 hold249 (.A(\rf_ram.RAM[7][22] ),
    .X(net1629));
 sg13g2_dlygate4sd3_1 hold250 (.A(\rf_ram.RAM[12][0] ),
    .X(net1630));
 sg13g2_dlygate4sd3_1 hold251 (.A(_01124_),
    .X(net1631));
 sg13g2_dlygate4sd3_1 hold252 (.A(\rf_ram.RAM[26][29] ),
    .X(net1632));
 sg13g2_dlygate4sd3_1 hold253 (.A(\rf_ram.RAM[15][10] ),
    .X(net1633));
 sg13g2_dlygate4sd3_1 hold254 (.A(\rf_ram.RAM[4][3] ),
    .X(net1634));
 sg13g2_dlygate4sd3_1 hold255 (.A(\rf_ram.RAM[28][11] ),
    .X(net1635));
 sg13g2_dlygate4sd3_1 hold256 (.A(\rf_ram.RAM[18][0] ),
    .X(net1636));
 sg13g2_dlygate4sd3_1 hold257 (.A(\rf_ram.RAM[25][6] ),
    .X(net1637));
 sg13g2_dlygate4sd3_1 hold258 (.A(\rf_ram.RAM[5][9] ),
    .X(net1638));
 sg13g2_dlygate4sd3_1 hold259 (.A(\rf_ram.RAM[12][4] ),
    .X(net1639));
 sg13g2_dlygate4sd3_1 hold260 (.A(\rf_ram.RAM[22][15] ),
    .X(net1640));
 sg13g2_dlygate4sd3_1 hold261 (.A(\rf_ram.RAM[9][13] ),
    .X(net1641));
 sg13g2_dlygate4sd3_1 hold262 (.A(\rf_ram.RAM[6][13] ),
    .X(net1642));
 sg13g2_dlygate4sd3_1 hold263 (.A(\rf_ram.RAM[26][22] ),
    .X(net1643));
 sg13g2_dlygate4sd3_1 hold264 (.A(\rf_ram.RAM[14][3] ),
    .X(net1644));
 sg13g2_dlygate4sd3_1 hold265 (.A(\rf_ram.RAM[14][11] ),
    .X(net1645));
 sg13g2_dlygate4sd3_1 hold266 (.A(\rf_ram.RAM[25][7] ),
    .X(net1646));
 sg13g2_dlygate4sd3_1 hold267 (.A(\rf_ram.RAM[19][10] ),
    .X(net1647));
 sg13g2_dlygate4sd3_1 hold268 (.A(\rf_ram.RAM[4][18] ),
    .X(net1648));
 sg13g2_dlygate4sd3_1 hold269 (.A(\rf_ram.RAM[8][5] ),
    .X(net1649));
 sg13g2_dlygate4sd3_1 hold270 (.A(\rf_ram.RAM[14][13] ),
    .X(net1650));
 sg13g2_dlygate4sd3_1 hold271 (.A(\rf_ram.RAM[4][5] ),
    .X(net1651));
 sg13g2_dlygate4sd3_1 hold272 (.A(\rf_ram.RAM[23][25] ),
    .X(net1652));
 sg13g2_dlygate4sd3_1 hold273 (.A(\rf_ram.RAM[30][25] ),
    .X(net1653));
 sg13g2_dlygate4sd3_1 hold274 (.A(\rf_ram.RAM[18][2] ),
    .X(net1654));
 sg13g2_dlygate4sd3_1 hold275 (.A(\rf_ram.RAM[3][18] ),
    .X(net1655));
 sg13g2_dlygate4sd3_1 hold276 (.A(\rf_ram.RAM[0][8] ),
    .X(net1656));
 sg13g2_dlygate4sd3_1 hold277 (.A(\rf_ram.RAM[17][8] ),
    .X(net1657));
 sg13g2_dlygate4sd3_1 hold278 (.A(\rf_ram.RAM[14][5] ),
    .X(net1658));
 sg13g2_dlygate4sd3_1 hold279 (.A(\rf_ram.RAM[19][20] ),
    .X(net1659));
 sg13g2_dlygate4sd3_1 hold280 (.A(\rf_ram.RAM[24][11] ),
    .X(net1660));
 sg13g2_dlygate4sd3_1 hold281 (.A(\rf_ram.RAM[2][6] ),
    .X(net1661));
 sg13g2_dlygate4sd3_1 hold282 (.A(\rf_ram.RAM[18][24] ),
    .X(net1662));
 sg13g2_dlygate4sd3_1 hold283 (.A(\rf_ram.RAM[26][20] ),
    .X(net1663));
 sg13g2_dlygate4sd3_1 hold284 (.A(\rf_ram.RAM[28][22] ),
    .X(net1664));
 sg13g2_dlygate4sd3_1 hold285 (.A(\rf_ram.RAM[12][16] ),
    .X(net1665));
 sg13g2_dlygate4sd3_1 hold286 (.A(\rf_ram.RAM[23][0] ),
    .X(net1666));
 sg13g2_dlygate4sd3_1 hold287 (.A(\rf_ram.RAM[31][24] ),
    .X(net1667));
 sg13g2_dlygate4sd3_1 hold288 (.A(\rf_ram.RAM[12][31] ),
    .X(net1668));
 sg13g2_dlygate4sd3_1 hold289 (.A(\rf_ram.RAM[7][23] ),
    .X(net1669));
 sg13g2_dlygate4sd3_1 hold290 (.A(\rf_ram.RAM[11][12] ),
    .X(net1670));
 sg13g2_dlygate4sd3_1 hold291 (.A(\rf_ram.RAM[2][28] ),
    .X(net1671));
 sg13g2_dlygate4sd3_1 hold292 (.A(\rf_ram.RAM[12][15] ),
    .X(net1672));
 sg13g2_dlygate4sd3_1 hold293 (.A(\rf_ram.RAM[6][28] ),
    .X(net1673));
 sg13g2_dlygate4sd3_1 hold294 (.A(\rf_ram.RAM[5][25] ),
    .X(net1674));
 sg13g2_dlygate4sd3_1 hold295 (.A(_00941_),
    .X(net1675));
 sg13g2_dlygate4sd3_1 hold296 (.A(\rf_ram.RAM[10][31] ),
    .X(net1676));
 sg13g2_dlygate4sd3_1 hold297 (.A(\rf_ram.RAM[28][26] ),
    .X(net1677));
 sg13g2_dlygate4sd3_1 hold298 (.A(\rf_ram.RAM[16][25] ),
    .X(net1678));
 sg13g2_dlygate4sd3_1 hold299 (.A(\rf_ram.RAM[6][25] ),
    .X(net1679));
 sg13g2_dlygate4sd3_1 hold300 (.A(\rf_ram.RAM[12][12] ),
    .X(net1680));
 sg13g2_dlygate4sd3_1 hold301 (.A(\rf_ram.RAM[13][6] ),
    .X(net1681));
 sg13g2_dlygate4sd3_1 hold302 (.A(\rf_ram.RAM[23][10] ),
    .X(net1682));
 sg13g2_dlygate4sd3_1 hold303 (.A(\rf_ram.RAM[3][20] ),
    .X(net1683));
 sg13g2_dlygate4sd3_1 hold304 (.A(\rf_ram.RAM[8][6] ),
    .X(net1684));
 sg13g2_dlygate4sd3_1 hold305 (.A(\rf_ram.RAM[25][0] ),
    .X(net1685));
 sg13g2_dlygate4sd3_1 hold306 (.A(\rf_ram.RAM[26][3] ),
    .X(net1686));
 sg13g2_dlygate4sd3_1 hold307 (.A(\rf_ram.RAM[17][10] ),
    .X(net1687));
 sg13g2_dlygate4sd3_1 hold308 (.A(\rf_ram.RAM[22][16] ),
    .X(net1688));
 sg13g2_dlygate4sd3_1 hold309 (.A(\rf_ram.RAM[2][21] ),
    .X(net1689));
 sg13g2_dlygate4sd3_1 hold310 (.A(\rf_ram.RAM[16][5] ),
    .X(net1690));
 sg13g2_dlygate4sd3_1 hold311 (.A(\rf_ram.RAM[31][18] ),
    .X(net1691));
 sg13g2_dlygate4sd3_1 hold312 (.A(\rf_ram.RAM[22][9] ),
    .X(net1692));
 sg13g2_dlygate4sd3_1 hold313 (.A(\rf_ram.RAM[19][11] ),
    .X(net1693));
 sg13g2_dlygate4sd3_1 hold314 (.A(\rf_ram.RAM[12][23] ),
    .X(net1694));
 sg13g2_dlygate4sd3_1 hold315 (.A(\rf_ram.RAM[7][24] ),
    .X(net1695));
 sg13g2_dlygate4sd3_1 hold316 (.A(\rf_ram.RAM[22][0] ),
    .X(net1696));
 sg13g2_dlygate4sd3_1 hold317 (.A(_00247_),
    .X(net1697));
 sg13g2_dlygate4sd3_1 hold318 (.A(\rf_ram.RAM[19][25] ),
    .X(net1698));
 sg13g2_dlygate4sd3_1 hold319 (.A(\rf_ram.RAM[27][24] ),
    .X(net1699));
 sg13g2_dlygate4sd3_1 hold320 (.A(\rf_ram.RAM[23][2] ),
    .X(net1700));
 sg13g2_dlygate4sd3_1 hold321 (.A(\rf_ram.RAM[17][13] ),
    .X(net1701));
 sg13g2_dlygate4sd3_1 hold322 (.A(\rf_ram.RAM[7][9] ),
    .X(net1702));
 sg13g2_dlygate4sd3_1 hold323 (.A(\rf_ram.RAM[26][13] ),
    .X(net1703));
 sg13g2_dlygate4sd3_1 hold324 (.A(\rf_ram.RAM[12][28] ),
    .X(net1704));
 sg13g2_dlygate4sd3_1 hold325 (.A(\rf_ram.RAM[23][28] ),
    .X(net1705));
 sg13g2_dlygate4sd3_1 hold326 (.A(\rf_ram.RAM[30][16] ),
    .X(net1706));
 sg13g2_dlygate4sd3_1 hold327 (.A(\rf_ram.RAM[26][0] ),
    .X(net1707));
 sg13g2_dlygate4sd3_1 hold328 (.A(\rf_ram.RAM[5][18] ),
    .X(net1708));
 sg13g2_dlygate4sd3_1 hold329 (.A(\rf_ram.RAM[0][1] ),
    .X(net1709));
 sg13g2_dlygate4sd3_1 hold330 (.A(\rf_ram.RAM[15][22] ),
    .X(net1710));
 sg13g2_dlygate4sd3_1 hold331 (.A(\rf_ram.RAM[1][21] ),
    .X(net1711));
 sg13g2_dlygate4sd3_1 hold332 (.A(\rf_ram.RAM[31][11] ),
    .X(net1712));
 sg13g2_dlygate4sd3_1 hold333 (.A(\rf_ram.RAM[1][5] ),
    .X(net1713));
 sg13g2_dlygate4sd3_1 hold334 (.A(\rf_ram.RAM[30][3] ),
    .X(net1714));
 sg13g2_dlygate4sd3_1 hold335 (.A(\rf_ram.RAM[28][18] ),
    .X(net1715));
 sg13g2_dlygate4sd3_1 hold336 (.A(\rf_ram.RAM[7][10] ),
    .X(net1716));
 sg13g2_dlygate4sd3_1 hold337 (.A(\rf_ram.RAM[25][12] ),
    .X(net1717));
 sg13g2_dlygate4sd3_1 hold338 (.A(\rf_ram.RAM[8][4] ),
    .X(net1718));
 sg13g2_dlygate4sd3_1 hold339 (.A(\rf_ram.RAM[3][6] ),
    .X(net1719));
 sg13g2_dlygate4sd3_1 hold340 (.A(\rf_ram.RAM[27][17] ),
    .X(net1720));
 sg13g2_dlygate4sd3_1 hold341 (.A(\rf_ram.RAM[30][9] ),
    .X(net1721));
 sg13g2_dlygate4sd3_1 hold342 (.A(\rf_ram.RAM[14][24] ),
    .X(net1722));
 sg13g2_dlygate4sd3_1 hold343 (.A(\rf_ram.RAM[2][30] ),
    .X(net1723));
 sg13g2_dlygate4sd3_1 hold344 (.A(\rf_ram.RAM[24][19] ),
    .X(net1724));
 sg13g2_dlygate4sd3_1 hold345 (.A(\rf_ram.RAM[6][26] ),
    .X(net1725));
 sg13g2_dlygate4sd3_1 hold346 (.A(\rf_ram.RAM[22][5] ),
    .X(net1726));
 sg13g2_dlygate4sd3_1 hold347 (.A(\rf_ram.RAM[23][22] ),
    .X(net1727));
 sg13g2_dlygate4sd3_1 hold348 (.A(\rf_ram.RAM[31][7] ),
    .X(net1728));
 sg13g2_dlygate4sd3_1 hold349 (.A(\rf_ram.RAM[12][17] ),
    .X(net1729));
 sg13g2_dlygate4sd3_1 hold350 (.A(\rf_ram.RAM[3][2] ),
    .X(net1730));
 sg13g2_dlygate4sd3_1 hold351 (.A(\rf_ram.RAM[27][31] ),
    .X(net1731));
 sg13g2_dlygate4sd3_1 hold352 (.A(\rf_ram.RAM[1][20] ),
    .X(net1732));
 sg13g2_dlygate4sd3_1 hold353 (.A(\rf_ram.RAM[12][10] ),
    .X(net1733));
 sg13g2_dlygate4sd3_1 hold354 (.A(\rf_ram.RAM[1][12] ),
    .X(net1734));
 sg13g2_dlygate4sd3_1 hold355 (.A(\rf_ram.RAM[19][7] ),
    .X(net1735));
 sg13g2_dlygate4sd3_1 hold356 (.A(\rf_ram.RAM[20][14] ),
    .X(net1736));
 sg13g2_dlygate4sd3_1 hold357 (.A(\rf_ram.RAM[19][2] ),
    .X(net1737));
 sg13g2_dlygate4sd3_1 hold358 (.A(\rf_ram.RAM[16][27] ),
    .X(net1738));
 sg13g2_dlygate4sd3_1 hold359 (.A(\rf_ram.RAM[28][6] ),
    .X(net1739));
 sg13g2_dlygate4sd3_1 hold360 (.A(\rf_ram.RAM[21][30] ),
    .X(net1740));
 sg13g2_dlygate4sd3_1 hold361 (.A(\rf_ram.RAM[22][23] ),
    .X(net1741));
 sg13g2_dlygate4sd3_1 hold362 (.A(\rf_ram.RAM[24][21] ),
    .X(net1742));
 sg13g2_dlygate4sd3_1 hold363 (.A(\rf_ram.RAM[9][23] ),
    .X(net1743));
 sg13g2_dlygate4sd3_1 hold364 (.A(\rf_ram.RAM[5][19] ),
    .X(net1744));
 sg13g2_dlygate4sd3_1 hold365 (.A(\rf_ram.RAM[14][18] ),
    .X(net1745));
 sg13g2_dlygate4sd3_1 hold366 (.A(\rf_ram.RAM[16][8] ),
    .X(net1746));
 sg13g2_dlygate4sd3_1 hold367 (.A(\rf_ram.RAM[14][14] ),
    .X(net1747));
 sg13g2_dlygate4sd3_1 hold368 (.A(\rf_ram.RAM[27][18] ),
    .X(net1748));
 sg13g2_dlygate4sd3_1 hold369 (.A(\rf_ram.RAM[6][9] ),
    .X(net2603));
 sg13g2_dlygate4sd3_1 hold370 (.A(\rf_ram.RAM[11][22] ),
    .X(net2604));
 sg13g2_dlygate4sd3_1 hold371 (.A(\rf_ram.RAM[12][6] ),
    .X(net2605));
 sg13g2_dlygate4sd3_1 hold372 (.A(\rf_ram.RAM[2][20] ),
    .X(net2606));
 sg13g2_dlygate4sd3_1 hold373 (.A(\rf_ram.RAM[0][3] ),
    .X(net2607));
 sg13g2_dlygate4sd3_1 hold374 (.A(\rf_ram.RAM[7][18] ),
    .X(net2608));
 sg13g2_dlygate4sd3_1 hold375 (.A(\rf_ram.RAM[7][20] ),
    .X(net2609));
 sg13g2_dlygate4sd3_1 hold376 (.A(\rf_ram.RAM[2][5] ),
    .X(net2610));
 sg13g2_dlygate4sd3_1 hold377 (.A(\rf_ram.RAM[0][29] ),
    .X(net2611));
 sg13g2_dlygate4sd3_1 hold378 (.A(\rf_ram.RAM[24][1] ),
    .X(net2612));
 sg13g2_dlygate4sd3_1 hold379 (.A(\rf_ram.RAM[6][4] ),
    .X(net2613));
 sg13g2_dlygate4sd3_1 hold380 (.A(\rf_ram.RAM[4][28] ),
    .X(net2614));
 sg13g2_dlygate4sd3_1 hold381 (.A(\rf_ram.RAM[21][18] ),
    .X(net2615));
 sg13g2_dlygate4sd3_1 hold382 (.A(\rf_ram.RAM[27][25] ),
    .X(net2616));
 sg13g2_dlygate4sd3_1 hold383 (.A(\rf_ram.RAM[3][28] ),
    .X(net2617));
 sg13g2_dlygate4sd3_1 hold384 (.A(\rf_ram.RAM[4][14] ),
    .X(net2618));
 sg13g2_dlygate4sd3_1 hold385 (.A(\rf_ram.RAM[22][13] ),
    .X(net2619));
 sg13g2_dlygate4sd3_1 hold386 (.A(\rf_ram.RAM[29][1] ),
    .X(net2620));
 sg13g2_dlygate4sd3_1 hold387 (.A(\rf_ram.RAM[17][9] ),
    .X(net2621));
 sg13g2_dlygate4sd3_1 hold388 (.A(\rf_ram.RAM[13][7] ),
    .X(net2622));
 sg13g2_dlygate4sd3_1 hold389 (.A(\rf_ram.RAM[7][21] ),
    .X(net2623));
 sg13g2_dlygate4sd3_1 hold390 (.A(\rf_ram.RAM[29][24] ),
    .X(net2624));
 sg13g2_dlygate4sd3_1 hold391 (.A(\rf_ram.RAM[0][5] ),
    .X(net2625));
 sg13g2_dlygate4sd3_1 hold392 (.A(\rf_ram.RAM[7][19] ),
    .X(net2626));
 sg13g2_dlygate4sd3_1 hold393 (.A(\rf_ram.RAM[14][4] ),
    .X(net2627));
 sg13g2_dlygate4sd3_1 hold394 (.A(\rf_ram.RAM[27][26] ),
    .X(net2628));
 sg13g2_dlygate4sd3_1 hold395 (.A(\rf_ram.RAM[2][9] ),
    .X(net2629));
 sg13g2_dlygate4sd3_1 hold396 (.A(\rf_ram.RAM[17][23] ),
    .X(net2630));
 sg13g2_dlygate4sd3_1 hold397 (.A(\rf_ram.RAM[4][15] ),
    .X(net2631));
 sg13g2_dlygate4sd3_1 hold398 (.A(\rf_ram.RAM[16][16] ),
    .X(net2632));
 sg13g2_dlygate4sd3_1 hold399 (.A(\rf_ram.RAM[14][21] ),
    .X(net2633));
 sg13g2_dlygate4sd3_1 hold400 (.A(\rf_ram.RAM[21][2] ),
    .X(net2634));
 sg13g2_dlygate4sd3_1 hold401 (.A(\rf_ram.RAM[27][11] ),
    .X(net2635));
 sg13g2_dlygate4sd3_1 hold402 (.A(\rf_ram.RAM[29][20] ),
    .X(net2636));
 sg13g2_dlygate4sd3_1 hold403 (.A(\rf_ram.RAM[24][8] ),
    .X(net2637));
 sg13g2_dlygate4sd3_1 hold404 (.A(\rf_ram.RAM[10][19] ),
    .X(net2638));
 sg13g2_dlygate4sd3_1 hold405 (.A(\rf_ram.RAM[14][31] ),
    .X(net2639));
 sg13g2_dlygate4sd3_1 hold406 (.A(\rf_ram.RAM[19][5] ),
    .X(net2640));
 sg13g2_dlygate4sd3_1 hold407 (.A(\rf_ram.RAM[22][22] ),
    .X(net2641));
 sg13g2_dlygate4sd3_1 hold408 (.A(\rf_ram.RAM[10][5] ),
    .X(net2642));
 sg13g2_dlygate4sd3_1 hold409 (.A(\rf_ram.RAM[22][17] ),
    .X(net2643));
 sg13g2_dlygate4sd3_1 hold410 (.A(\rf_ram.RAM[1][8] ),
    .X(net2644));
 sg13g2_dlygate4sd3_1 hold411 (.A(\rf_ram.RAM[18][15] ),
    .X(net2645));
 sg13g2_dlygate4sd3_1 hold412 (.A(\rf_ram.RAM[25][4] ),
    .X(net2646));
 sg13g2_dlygate4sd3_1 hold413 (.A(\rf_ram.RAM[6][11] ),
    .X(net2647));
 sg13g2_dlygate4sd3_1 hold414 (.A(\rf_ram.RAM[25][22] ),
    .X(net2648));
 sg13g2_dlygate4sd3_1 hold415 (.A(\rf_ram.RAM[25][19] ),
    .X(net2649));
 sg13g2_dlygate4sd3_1 hold416 (.A(\rf_ram.RAM[21][4] ),
    .X(net2650));
 sg13g2_dlygate4sd3_1 hold417 (.A(\rf_ram.RAM[7][2] ),
    .X(net2651));
 sg13g2_dlygate4sd3_1 hold418 (.A(\rf_ram.RAM[13][16] ),
    .X(net2652));
 sg13g2_dlygate4sd3_1 hold419 (.A(\rf_ram.RAM[0][16] ),
    .X(net2653));
 sg13g2_dlygate4sd3_1 hold420 (.A(\rf_ram.RAM[22][26] ),
    .X(net2654));
 sg13g2_dlygate4sd3_1 hold421 (.A(\rf_ram.RAM[19][24] ),
    .X(net2655));
 sg13g2_dlygate4sd3_1 hold422 (.A(\rf_ram.RAM[16][24] ),
    .X(net2656));
 sg13g2_dlygate4sd3_1 hold423 (.A(\rf_ram.RAM[27][3] ),
    .X(net2657));
 sg13g2_dlygate4sd3_1 hold424 (.A(\rf_ram.RAM[24][4] ),
    .X(net2658));
 sg13g2_dlygate4sd3_1 hold425 (.A(\rf_ram.RAM[5][3] ),
    .X(net2659));
 sg13g2_dlygate4sd3_1 hold426 (.A(\rf_ram.RAM[4][30] ),
    .X(net2660));
 sg13g2_dlygate4sd3_1 hold427 (.A(\rf_ram.RAM[15][16] ),
    .X(net2661));
 sg13g2_dlygate4sd3_1 hold428 (.A(\rf_ram.RAM[25][1] ),
    .X(net2662));
 sg13g2_dlygate4sd3_1 hold429 (.A(\rf_ram.RAM[1][4] ),
    .X(net2663));
 sg13g2_dlygate4sd3_1 hold430 (.A(\rf_ram.RAM[22][2] ),
    .X(net2664));
 sg13g2_dlygate4sd3_1 hold431 (.A(\rf_ram.RAM[1][3] ),
    .X(net2665));
 sg13g2_dlygate4sd3_1 hold432 (.A(\rf_ram.RAM[24][7] ),
    .X(net2666));
 sg13g2_dlygate4sd3_1 hold433 (.A(\rf_ram.RAM[3][5] ),
    .X(net2667));
 sg13g2_dlygate4sd3_1 hold434 (.A(\rf_ram.RAM[15][26] ),
    .X(net2668));
 sg13g2_dlygate4sd3_1 hold435 (.A(\rf_ram.RAM[7][25] ),
    .X(net2669));
 sg13g2_dlygate4sd3_1 hold436 (.A(\rf_ram.RAM[30][20] ),
    .X(net2670));
 sg13g2_dlygate4sd3_1 hold437 (.A(\rf_ram.RAM[22][12] ),
    .X(net2671));
 sg13g2_dlygate4sd3_1 hold438 (.A(\rf_ram.RAM[7][4] ),
    .X(net2672));
 sg13g2_dlygate4sd3_1 hold439 (.A(\rf_ram.RAM[6][31] ),
    .X(net2673));
 sg13g2_dlygate4sd3_1 hold440 (.A(\rf_ram.RAM[10][22] ),
    .X(net2674));
 sg13g2_dlygate4sd3_1 hold441 (.A(\rf_ram.RAM[22][24] ),
    .X(net2675));
 sg13g2_dlygate4sd3_1 hold442 (.A(\rf_ram.RAM[28][17] ),
    .X(net2676));
 sg13g2_dlygate4sd3_1 hold443 (.A(\rf_ram.RAM[25][10] ),
    .X(net2677));
 sg13g2_dlygate4sd3_1 hold444 (.A(\rf_ram.RAM[18][30] ),
    .X(net2678));
 sg13g2_dlygate4sd3_1 hold445 (.A(\rf_ram.RAM[27][28] ),
    .X(net2679));
 sg13g2_dlygate4sd3_1 hold446 (.A(\rf_ram.RAM[30][14] ),
    .X(net2680));
 sg13g2_dlygate4sd3_1 hold447 (.A(\rf_ram.RAM[2][3] ),
    .X(net2681));
 sg13g2_dlygate4sd3_1 hold448 (.A(\rf_ram.RAM[1][6] ),
    .X(net2682));
 sg13g2_dlygate4sd3_1 hold449 (.A(\rf_ram.RAM[24][0] ),
    .X(net2683));
 sg13g2_dlygate4sd3_1 hold450 (.A(\rf_ram.RAM[12][30] ),
    .X(net2684));
 sg13g2_dlygate4sd3_1 hold451 (.A(\rf_ram.RAM[22][27] ),
    .X(net2685));
 sg13g2_dlygate4sd3_1 hold452 (.A(\rf_ram.RAM[15][7] ),
    .X(net2686));
 sg13g2_dlygate4sd3_1 hold453 (.A(\rf_ram.RAM[28][3] ),
    .X(net2687));
 sg13g2_dlygate4sd3_1 hold454 (.A(\rf_ram.RAM[11][27] ),
    .X(net2688));
 sg13g2_dlygate4sd3_1 hold455 (.A(\rf_ram.RAM[0][28] ),
    .X(net2689));
 sg13g2_dlygate4sd3_1 hold456 (.A(\rf_ram.RAM[5][16] ),
    .X(net2690));
 sg13g2_dlygate4sd3_1 hold457 (.A(\rf_ram.RAM[28][30] ),
    .X(net2691));
 sg13g2_dlygate4sd3_1 hold458 (.A(\rf_ram.RAM[4][20] ),
    .X(net2692));
 sg13g2_dlygate4sd3_1 hold459 (.A(\rf_ram.RAM[26][6] ),
    .X(net2693));
 sg13g2_dlygate4sd3_1 hold460 (.A(\rf_ram.RAM[6][17] ),
    .X(net2694));
 sg13g2_dlygate4sd3_1 hold461 (.A(\rf_ram.RAM[11][14] ),
    .X(net2695));
 sg13g2_dlygate4sd3_1 hold462 (.A(\rf_ram.RAM[14][6] ),
    .X(net2696));
 sg13g2_dlygate4sd3_1 hold463 (.A(\rf_ram.RAM[16][6] ),
    .X(net2697));
 sg13g2_dlygate4sd3_1 hold464 (.A(\rf_ram.RAM[26][31] ),
    .X(net2698));
 sg13g2_dlygate4sd3_1 hold465 (.A(\rf_ram.RAM[31][6] ),
    .X(net2699));
 sg13g2_dlygate4sd3_1 hold466 (.A(\rf_ram.RAM[26][2] ),
    .X(net2700));
 sg13g2_dlygate4sd3_1 hold467 (.A(\rf_ram.RAM[6][10] ),
    .X(net2701));
 sg13g2_dlygate4sd3_1 hold468 (.A(\rf_ram.RAM[9][30] ),
    .X(net2702));
 sg13g2_dlygate4sd3_1 hold469 (.A(\rf_ram.RAM[2][31] ),
    .X(net2703));
 sg13g2_dlygate4sd3_1 hold470 (.A(\rf_ram.RAM[21][7] ),
    .X(net2704));
 sg13g2_dlygate4sd3_1 hold471 (.A(\rf_ram.RAM[31][25] ),
    .X(net2705));
 sg13g2_dlygate4sd3_1 hold472 (.A(\rf_ram.RAM[9][15] ),
    .X(net2706));
 sg13g2_dlygate4sd3_1 hold473 (.A(\rf_ram.RAM[4][1] ),
    .X(net2707));
 sg13g2_dlygate4sd3_1 hold474 (.A(\rf_ram.RAM[18][9] ),
    .X(net2708));
 sg13g2_dlygate4sd3_1 hold475 (.A(\rf_ram.RAM[7][29] ),
    .X(net2709));
 sg13g2_dlygate4sd3_1 hold476 (.A(\rf_ram.RAM[16][1] ),
    .X(net2710));
 sg13g2_dlygate4sd3_1 hold477 (.A(\rf_ram.RAM[13][0] ),
    .X(net2711));
 sg13g2_dlygate4sd3_1 hold478 (.A(_01092_),
    .X(net2712));
 sg13g2_dlygate4sd3_1 hold479 (.A(\rf_ram.RAM[17][5] ),
    .X(net2713));
 sg13g2_dlygate4sd3_1 hold480 (.A(\rf_ram.RAM[14][10] ),
    .X(net2714));
 sg13g2_dlygate4sd3_1 hold481 (.A(\rf_ram.RAM[30][28] ),
    .X(net2715));
 sg13g2_dlygate4sd3_1 hold482 (.A(\rf_ram.RAM[11][9] ),
    .X(net2716));
 sg13g2_dlygate4sd3_1 hold483 (.A(\rf_ram.RAM[5][6] ),
    .X(net2717));
 sg13g2_dlygate4sd3_1 hold484 (.A(\rf_ram.RAM[15][9] ),
    .X(net2718));
 sg13g2_dlygate4sd3_1 hold485 (.A(\rf_ram.RAM[28][0] ),
    .X(net2719));
 sg13g2_dlygate4sd3_1 hold486 (.A(_01060_),
    .X(net2720));
 sg13g2_dlygate4sd3_1 hold487 (.A(\rf_ram.RAM[13][27] ),
    .X(net2721));
 sg13g2_dlygate4sd3_1 hold488 (.A(\rf_ram.RAM[10][15] ),
    .X(net2722));
 sg13g2_dlygate4sd3_1 hold489 (.A(\rf_ram.RAM[5][17] ),
    .X(net2723));
 sg13g2_dlygate4sd3_1 hold490 (.A(\rf_ram.RAM[4][24] ),
    .X(net2724));
 sg13g2_dlygate4sd3_1 hold491 (.A(\rf_ram.RAM[15][23] ),
    .X(net2725));
 sg13g2_dlygate4sd3_1 hold492 (.A(\rf_ram.RAM[26][17] ),
    .X(net2726));
 sg13g2_dlygate4sd3_1 hold493 (.A(\rf_ram.RAM[1][13] ),
    .X(net2727));
 sg13g2_dlygate4sd3_1 hold494 (.A(\rf_ram.RAM[6][19] ),
    .X(net2728));
 sg13g2_dlygate4sd3_1 hold495 (.A(\rf_ram.RAM[18][19] ),
    .X(net2729));
 sg13g2_dlygate4sd3_1 hold496 (.A(\rf_ram.RAM[18][27] ),
    .X(net2730));
 sg13g2_dlygate4sd3_1 hold497 (.A(\rf_ram.RAM[14][27] ),
    .X(net2731));
 sg13g2_dlygate4sd3_1 hold498 (.A(\rf_ram.RAM[4][31] ),
    .X(net2732));
 sg13g2_dlygate4sd3_1 hold499 (.A(\rf_ram.RAM[1][24] ),
    .X(net2733));
 sg13g2_dlygate4sd3_1 hold500 (.A(\rf_ram.RAM[11][15] ),
    .X(net2734));
 sg13g2_dlygate4sd3_1 hold501 (.A(\rf_ram.RAM[1][27] ),
    .X(net2735));
 sg13g2_dlygate4sd3_1 hold502 (.A(\rf_ram.RAM[6][23] ),
    .X(net2736));
 sg13g2_dlygate4sd3_1 hold503 (.A(\rf_ram.RAM[26][15] ),
    .X(net2737));
 sg13g2_dlygate4sd3_1 hold504 (.A(\rf_ram.RAM[1][9] ),
    .X(net2738));
 sg13g2_dlygate4sd3_1 hold505 (.A(\rf_ram.RAM[9][4] ),
    .X(net2739));
 sg13g2_dlygate4sd3_1 hold506 (.A(\rf_ram.RAM[1][0] ),
    .X(net2740));
 sg13g2_dlygate4sd3_1 hold507 (.A(_00151_),
    .X(net2741));
 sg13g2_dlygate4sd3_1 hold508 (.A(\rf_ram.RAM[18][4] ),
    .X(net2742));
 sg13g2_dlygate4sd3_1 hold509 (.A(\rf_ram.RAM[17][25] ),
    .X(net2743));
 sg13g2_dlygate4sd3_1 hold510 (.A(\rf_ram.RAM[3][11] ),
    .X(net2744));
 sg13g2_dlygate4sd3_1 hold511 (.A(\rf_ram.RAM[1][16] ),
    .X(net2745));
 sg13g2_dlygate4sd3_1 hold512 (.A(\rf_ram.RAM[20][24] ),
    .X(net2746));
 sg13g2_dlygate4sd3_1 hold513 (.A(\rf_ram.RAM[23][11] ),
    .X(net2747));
 sg13g2_dlygate4sd3_1 hold514 (.A(\rf_ram.RAM[17][29] ),
    .X(net2748));
 sg13g2_dlygate4sd3_1 hold515 (.A(\rf_ram.RAM[14][2] ),
    .X(net2749));
 sg13g2_dlygate4sd3_1 hold516 (.A(\rf_ram.RAM[23][3] ),
    .X(net2750));
 sg13g2_dlygate4sd3_1 hold517 (.A(\rf_ram.RAM[30][10] ),
    .X(net2751));
 sg13g2_dlygate4sd3_1 hold518 (.A(\rf_ram.RAM[12][25] ),
    .X(net2752));
 sg13g2_dlygate4sd3_1 hold519 (.A(\rf_ram.RAM[6][30] ),
    .X(net2753));
 sg13g2_dlygate4sd3_1 hold520 (.A(\rf_ram.RAM[6][27] ),
    .X(net2754));
 sg13g2_dlygate4sd3_1 hold521 (.A(\rf_ram.RAM[17][24] ),
    .X(net2755));
 sg13g2_dlygate4sd3_1 hold522 (.A(\rf_ram.RAM[20][17] ),
    .X(net2756));
 sg13g2_dlygate4sd3_1 hold523 (.A(\rf_ram.RAM[19][12] ),
    .X(net2757));
 sg13g2_dlygate4sd3_1 hold524 (.A(\rf_ram.RAM[24][16] ),
    .X(net2758));
 sg13g2_dlygate4sd3_1 hold525 (.A(\rf_ram.RAM[10][24] ),
    .X(net2759));
 sg13g2_dlygate4sd3_1 hold526 (.A(\rf_ram.RAM[11][18] ),
    .X(net2760));
 sg13g2_dlygate4sd3_1 hold527 (.A(\rf_ram.RAM[13][12] ),
    .X(net2761));
 sg13g2_dlygate4sd3_1 hold528 (.A(\rf_ram.RAM[6][6] ),
    .X(net2762));
 sg13g2_dlygate4sd3_1 hold529 (.A(\rf_ram.RAM[22][7] ),
    .X(net2763));
 sg13g2_dlygate4sd3_1 hold530 (.A(\rf_ram.RAM[17][27] ),
    .X(net2764));
 sg13g2_dlygate4sd3_1 hold531 (.A(\rf_ram.RAM[8][30] ),
    .X(net2765));
 sg13g2_dlygate4sd3_1 hold532 (.A(\rf_ram.RAM[31][4] ),
    .X(net2766));
 sg13g2_dlygate4sd3_1 hold533 (.A(\rf_ram.RAM[30][27] ),
    .X(net2767));
 sg13g2_dlygate4sd3_1 hold534 (.A(\rf_ram.RAM[27][1] ),
    .X(net2768));
 sg13g2_dlygate4sd3_1 hold535 (.A(\rf_ram.RAM[16][21] ),
    .X(net2769));
 sg13g2_dlygate4sd3_1 hold536 (.A(\rf_ram.RAM[30][4] ),
    .X(net2770));
 sg13g2_dlygate4sd3_1 hold537 (.A(\rf_ram.RAM[17][17] ),
    .X(net2771));
 sg13g2_dlygate4sd3_1 hold538 (.A(\rf_ram.RAM[17][4] ),
    .X(net2772));
 sg13g2_dlygate4sd3_1 hold539 (.A(\rf_ram.RAM[21][16] ),
    .X(net2773));
 sg13g2_dlygate4sd3_1 hold540 (.A(\rf_ram.RAM[6][21] ),
    .X(net2774));
 sg13g2_dlygate4sd3_1 hold541 (.A(\rf_ram.RAM[11][8] ),
    .X(net2775));
 sg13g2_dlygate4sd3_1 hold542 (.A(\rf_ram.RAM[16][2] ),
    .X(net2776));
 sg13g2_dlygate4sd3_1 hold543 (.A(\rf_ram.RAM[13][4] ),
    .X(net2777));
 sg13g2_dlygate4sd3_1 hold544 (.A(\rf_ram.RAM[15][3] ),
    .X(net2778));
 sg13g2_dlygate4sd3_1 hold545 (.A(\rf_ram.RAM[0][27] ),
    .X(net2779));
 sg13g2_dlygate4sd3_1 hold546 (.A(\rf_ram.RAM[0][18] ),
    .X(net2780));
 sg13g2_dlygate4sd3_1 hold547 (.A(\rf_ram.RAM[7][5] ),
    .X(net2781));
 sg13g2_dlygate4sd3_1 hold548 (.A(\rf_ram.RAM[22][28] ),
    .X(net2782));
 sg13g2_dlygate4sd3_1 hold549 (.A(\rf_ram.RAM[31][16] ),
    .X(net2783));
 sg13g2_dlygate4sd3_1 hold550 (.A(\rf_ram.RAM[31][27] ),
    .X(net2784));
 sg13g2_dlygate4sd3_1 hold551 (.A(\rf_ram.RAM[5][1] ),
    .X(net2785));
 sg13g2_dlygate4sd3_1 hold552 (.A(\rf_ram.RAM[0][20] ),
    .X(net2786));
 sg13g2_dlygate4sd3_1 hold553 (.A(\rf_ram.RAM[11][24] ),
    .X(net2787));
 sg13g2_dlygate4sd3_1 hold554 (.A(\rf_ram.RAM[20][5] ),
    .X(net2788));
 sg13g2_dlygate4sd3_1 hold555 (.A(\rf_ram.RAM[31][26] ),
    .X(net2789));
 sg13g2_dlygate4sd3_1 hold556 (.A(\rf_ram.RAM[30][24] ),
    .X(net2790));
 sg13g2_dlygate4sd3_1 hold557 (.A(\rf_ram.RAM[20][2] ),
    .X(net2791));
 sg13g2_dlygate4sd3_1 hold558 (.A(\rf_ram.RAM[29][22] ),
    .X(net2792));
 sg13g2_dlygate4sd3_1 hold559 (.A(\rf_ram.RAM[15][30] ),
    .X(net2793));
 sg13g2_dlygate4sd3_1 hold560 (.A(\rf_ram.RAM[8][8] ),
    .X(net2794));
 sg13g2_dlygate4sd3_1 hold561 (.A(\rf_ram.RAM[30][7] ),
    .X(net2795));
 sg13g2_dlygate4sd3_1 hold562 (.A(\rf_ram.RAM[25][18] ),
    .X(net2796));
 sg13g2_dlygate4sd3_1 hold563 (.A(\rf_ram.RAM[17][21] ),
    .X(net2797));
 sg13g2_dlygate4sd3_1 hold564 (.A(\rf_ram.RAM[28][12] ),
    .X(net2798));
 sg13g2_dlygate4sd3_1 hold565 (.A(\rf_ram.RAM[7][16] ),
    .X(net2799));
 sg13g2_dlygate4sd3_1 hold566 (.A(\rf_ram.RAM[8][1] ),
    .X(net2800));
 sg13g2_dlygate4sd3_1 hold567 (.A(\rf_ram.RAM[21][19] ),
    .X(net2801));
 sg13g2_dlygate4sd3_1 hold568 (.A(\rf_ram.RAM[11][21] ),
    .X(net2802));
 sg13g2_dlygate4sd3_1 hold569 (.A(\rf_ram.RAM[24][3] ),
    .X(net2803));
 sg13g2_dlygate4sd3_1 hold570 (.A(\rf_ram.RAM[5][26] ),
    .X(net2804));
 sg13g2_dlygate4sd3_1 hold571 (.A(\rf_ram.RAM[21][22] ),
    .X(net2805));
 sg13g2_dlygate4sd3_1 hold572 (.A(\rf_ram.RAM[11][16] ),
    .X(net2806));
 sg13g2_dlygate4sd3_1 hold573 (.A(\rf_ram.RAM[17][0] ),
    .X(net2807));
 sg13g2_dlygate4sd3_1 hold574 (.A(\rf_ram.RAM[6][3] ),
    .X(net2808));
 sg13g2_dlygate4sd3_1 hold575 (.A(\rf_ram.RAM[29][12] ),
    .X(net2809));
 sg13g2_dlygate4sd3_1 hold576 (.A(\rf_ram.RAM[31][0] ),
    .X(net2810));
 sg13g2_dlygate4sd3_1 hold577 (.A(_00339_),
    .X(net2811));
 sg13g2_dlygate4sd3_1 hold578 (.A(\rf_ram.RAM[21][6] ),
    .X(net2812));
 sg13g2_dlygate4sd3_1 hold579 (.A(\rf_ram.RAM[16][20] ),
    .X(net2813));
 sg13g2_dlygate4sd3_1 hold580 (.A(\rf_ram.RAM[14][16] ),
    .X(net2814));
 sg13g2_dlygate4sd3_1 hold581 (.A(\rf_ram.RAM[28][27] ),
    .X(net2815));
 sg13g2_dlygate4sd3_1 hold582 (.A(\rf_ram.RAM[4][9] ),
    .X(net2816));
 sg13g2_dlygate4sd3_1 hold583 (.A(\rf_ram.RAM[29][17] ),
    .X(net2817));
 sg13g2_dlygate4sd3_1 hold584 (.A(\rf_ram.RAM[21][27] ),
    .X(net2818));
 sg13g2_dlygate4sd3_1 hold585 (.A(\rf_ram.RAM[9][7] ),
    .X(net2819));
 sg13g2_dlygate4sd3_1 hold586 (.A(\rf_ram.RAM[5][14] ),
    .X(net2820));
 sg13g2_dlygate4sd3_1 hold587 (.A(\rf_ram.RAM[5][22] ),
    .X(net2821));
 sg13g2_dlygate4sd3_1 hold588 (.A(\rf_ram.RAM[20][7] ),
    .X(net2822));
 sg13g2_dlygate4sd3_1 hold589 (.A(\rf_ram.RAM[31][15] ),
    .X(net2823));
 sg13g2_dlygate4sd3_1 hold590 (.A(\rf_ram.RAM[6][0] ),
    .X(net2824));
 sg13g2_dlygate4sd3_1 hold591 (.A(_00852_),
    .X(net2825));
 sg13g2_dlygate4sd3_1 hold592 (.A(\rf_ram.RAM[21][14] ),
    .X(net2826));
 sg13g2_dlygate4sd3_1 hold593 (.A(\rf_ram.RAM[28][25] ),
    .X(net2827));
 sg13g2_dlygate4sd3_1 hold594 (.A(\rf_ram.RAM[8][16] ),
    .X(net2828));
 sg13g2_dlygate4sd3_1 hold595 (.A(\rf_ram.RAM[8][0] ),
    .X(net2829));
 sg13g2_dlygate4sd3_1 hold596 (.A(_01284_),
    .X(net2830));
 sg13g2_dlygate4sd3_1 hold597 (.A(\rf_ram.RAM[0][2] ),
    .X(net2831));
 sg13g2_dlygate4sd3_1 hold598 (.A(\rf_ram.RAM[30][18] ),
    .X(net2832));
 sg13g2_dlygate4sd3_1 hold599 (.A(\rf_ram.RAM[14][12] ),
    .X(net2833));
 sg13g2_dlygate4sd3_1 hold600 (.A(\rf_ram.RAM[27][30] ),
    .X(net2834));
 sg13g2_dlygate4sd3_1 hold601 (.A(\rf_ram.RAM[8][18] ),
    .X(net2835));
 sg13g2_dlygate4sd3_1 hold602 (.A(\rf_ram.RAM[2][4] ),
    .X(net2836));
 sg13g2_dlygate4sd3_1 hold603 (.A(\rf_ram.RAM[10][7] ),
    .X(net2837));
 sg13g2_dlygate4sd3_1 hold604 (.A(\rf_ram.RAM[5][24] ),
    .X(net2838));
 sg13g2_dlygate4sd3_1 hold605 (.A(\rf_ram.RAM[0][0] ),
    .X(net2839));
 sg13g2_dlygate4sd3_1 hold606 (.A(_01220_),
    .X(net2840));
 sg13g2_dlygate4sd3_1 hold607 (.A(\rf_ram.RAM[31][30] ),
    .X(net2841));
 sg13g2_dlygate4sd3_1 hold608 (.A(\rf_ram.RAM[7][28] ),
    .X(net2842));
 sg13g2_dlygate4sd3_1 hold609 (.A(\rf_ram.RAM[31][14] ),
    .X(net2843));
 sg13g2_dlygate4sd3_1 hold610 (.A(\rf_ram.RAM[0][12] ),
    .X(net2844));
 sg13g2_dlygate4sd3_1 hold611 (.A(\rf_ram.RAM[0][7] ),
    .X(net2845));
 sg13g2_dlygate4sd3_1 hold612 (.A(\rf_ram.RAM[6][8] ),
    .X(net2846));
 sg13g2_dlygate4sd3_1 hold613 (.A(\rf_ram.RAM[4][21] ),
    .X(net2847));
 sg13g2_dlygate4sd3_1 hold614 (.A(\rf_ram.RAM[9][10] ),
    .X(net2848));
 sg13g2_dlygate4sd3_1 hold615 (.A(\rf_ram.RAM[10][26] ),
    .X(net2849));
 sg13g2_dlygate4sd3_1 hold616 (.A(\rf_ram.RAM[3][9] ),
    .X(net2850));
 sg13g2_dlygate4sd3_1 hold617 (.A(\rf_ram.RAM[23][6] ),
    .X(net2851));
 sg13g2_dlygate4sd3_1 hold618 (.A(\rf_ram.RAM[30][5] ),
    .X(net2852));
 sg13g2_dlygate4sd3_1 hold619 (.A(\rf_ram.RAM[29][8] ),
    .X(net2853));
 sg13g2_dlygate4sd3_1 hold620 (.A(\rf_ram.RAM[19][13] ),
    .X(net2854));
 sg13g2_dlygate4sd3_1 hold621 (.A(\rf_ram.RAM[23][30] ),
    .X(net2855));
 sg13g2_dlygate4sd3_1 hold622 (.A(\rf_ram.RAM[10][18] ),
    .X(net2856));
 sg13g2_dlygate4sd3_1 hold623 (.A(\rf_ram.RAM[3][24] ),
    .X(net2857));
 sg13g2_dlygate4sd3_1 hold624 (.A(\rf_ram.RAM[7][11] ),
    .X(net2858));
 sg13g2_dlygate4sd3_1 hold625 (.A(\rf_ram.RAM[0][13] ),
    .X(net2859));
 sg13g2_dlygate4sd3_1 hold626 (.A(\rf_ram.RAM[19][19] ),
    .X(net2860));
 sg13g2_dlygate4sd3_1 hold627 (.A(\rf_ram.RAM[12][5] ),
    .X(net2861));
 sg13g2_dlygate4sd3_1 hold628 (.A(\rf_ram.RAM[21][31] ),
    .X(net2862));
 sg13g2_dlygate4sd3_1 hold629 (.A(\rf_ram.RAM[21][23] ),
    .X(net2863));
 sg13g2_dlygate4sd3_1 hold630 (.A(\rf_ram.RAM[31][23] ),
    .X(net2864));
 sg13g2_dlygate4sd3_1 hold631 (.A(\rf_ram.RAM[18][31] ),
    .X(net2865));
 sg13g2_dlygate4sd3_1 hold632 (.A(\rf_ram.RAM[13][8] ),
    .X(net2866));
 sg13g2_dlygate4sd3_1 hold633 (.A(\rf_ram.RAM[8][7] ),
    .X(net2867));
 sg13g2_dlygate4sd3_1 hold634 (.A(\rf_ram.RAM[3][15] ),
    .X(net2868));
 sg13g2_dlygate4sd3_1 hold635 (.A(\rf_ram.RAM[2][29] ),
    .X(net2869));
 sg13g2_dlygate4sd3_1 hold636 (.A(\rf_ram.RAM[19][21] ),
    .X(net2870));
 sg13g2_dlygate4sd3_1 hold637 (.A(\rf_ram.RAM[29][21] ),
    .X(net2871));
 sg13g2_dlygate4sd3_1 hold638 (.A(\rf_ram.RAM[14][25] ),
    .X(net2872));
 sg13g2_dlygate4sd3_1 hold639 (.A(\rf_ram.RAM[21][25] ),
    .X(net2873));
 sg13g2_dlygate4sd3_1 hold640 (.A(\rf_ram.RAM[24][6] ),
    .X(net2874));
 sg13g2_dlygate4sd3_1 hold641 (.A(\rf_ram.RAM[11][25] ),
    .X(net2875));
 sg13g2_dlygate4sd3_1 hold642 (.A(\rf_ram.RAM[18][29] ),
    .X(net2876));
 sg13g2_dlygate4sd3_1 hold643 (.A(\rf_ram.RAM[6][5] ),
    .X(net2877));
 sg13g2_dlygate4sd3_1 hold644 (.A(\rf_ram.RAM[30][11] ),
    .X(net2878));
 sg13g2_dlygate4sd3_1 hold645 (.A(\rf_ram.RAM[8][24] ),
    .X(net2879));
 sg13g2_dlygate4sd3_1 hold646 (.A(\rf_ram.RAM[31][8] ),
    .X(net2880));
 sg13g2_dlygate4sd3_1 hold647 (.A(\rf_ram.RAM[9][8] ),
    .X(net2881));
 sg13g2_dlygate4sd3_1 hold648 (.A(\rf_ram.RAM[14][30] ),
    .X(net2882));
 sg13g2_dlygate4sd3_1 hold649 (.A(\rf_ram.RAM[11][23] ),
    .X(net2883));
 sg13g2_dlygate4sd3_1 hold650 (.A(\rf_ram.RAM[18][18] ),
    .X(net2884));
 sg13g2_dlygate4sd3_1 hold651 (.A(\rf_ram.RAM[16][7] ),
    .X(net2885));
 sg13g2_dlygate4sd3_1 hold652 (.A(\rf_ram.RAM[9][22] ),
    .X(net2886));
 sg13g2_dlygate4sd3_1 hold653 (.A(\rf_ram.RAM[16][29] ),
    .X(net2887));
 sg13g2_dlygate4sd3_1 hold654 (.A(\rf_ram.RAM[11][4] ),
    .X(net2888));
 sg13g2_dlygate4sd3_1 hold655 (.A(\rf_ram.RAM[28][31] ),
    .X(net2889));
 sg13g2_dlygate4sd3_1 hold656 (.A(\rf_ram.RAM[17][6] ),
    .X(net2890));
 sg13g2_dlygate4sd3_1 hold657 (.A(\rf_ram.RAM[13][28] ),
    .X(net2891));
 sg13g2_dlygate4sd3_1 hold658 (.A(\rf_ram.RAM[13][22] ),
    .X(net2892));
 sg13g2_dlygate4sd3_1 hold659 (.A(\rf_ram.RAM[7][3] ),
    .X(net2893));
 sg13g2_dlygate4sd3_1 hold660 (.A(\rf_ram.RAM[24][14] ),
    .X(net2894));
 sg13g2_dlygate4sd3_1 hold661 (.A(\rf_ram.RAM[4][17] ),
    .X(net2895));
 sg13g2_dlygate4sd3_1 hold662 (.A(\rf_ram.RAM[16][10] ),
    .X(net2896));
 sg13g2_dlygate4sd3_1 hold663 (.A(\rf_ram.RAM[2][18] ),
    .X(net2897));
 sg13g2_dlygate4sd3_1 hold664 (.A(\rf_ram.RAM[14][0] ),
    .X(net2898));
 sg13g2_dlygate4sd3_1 hold665 (.A(_00752_),
    .X(net2899));
 sg13g2_dlygate4sd3_1 hold666 (.A(\rf_ram.RAM[5][27] ),
    .X(net2900));
 sg13g2_dlygate4sd3_1 hold667 (.A(\rf_ram.RAM[13][3] ),
    .X(net2901));
 sg13g2_dlygate4sd3_1 hold668 (.A(\rf_ram.RAM[28][28] ),
    .X(net2902));
 sg13g2_dlygate4sd3_1 hold669 (.A(\rf_ram.RAM[22][4] ),
    .X(net2903));
 sg13g2_dlygate4sd3_1 hold670 (.A(\rf_ram.RAM[10][14] ),
    .X(net2904));
 sg13g2_dlygate4sd3_1 hold671 (.A(\rf_ram.RAM[11][20] ),
    .X(net2905));
 sg13g2_dlygate4sd3_1 hold672 (.A(\rf_ram.RAM[24][29] ),
    .X(net2906));
 sg13g2_dlygate4sd3_1 hold673 (.A(\rf_ram.RAM[15][29] ),
    .X(net2907));
 sg13g2_dlygate4sd3_1 hold674 (.A(\rf_ram.RAM[29][25] ),
    .X(net2908));
 sg13g2_dlygate4sd3_1 hold675 (.A(\rf_ram.RAM[19][17] ),
    .X(net2909));
 sg13g2_dlygate4sd3_1 hold676 (.A(\rf_ram.RAM[3][27] ),
    .X(net2910));
 sg13g2_dlygate4sd3_1 hold677 (.A(\rf_ram.RAM[11][13] ),
    .X(net2911));
 sg13g2_dlygate4sd3_1 hold678 (.A(\rf_ram.RAM[26][23] ),
    .X(net2912));
 sg13g2_dlygate4sd3_1 hold679 (.A(\rf_ram.RAM[7][0] ),
    .X(net2913));
 sg13g2_dlygate4sd3_1 hold680 (.A(_00788_),
    .X(net2914));
 sg13g2_dlygate4sd3_1 hold681 (.A(\rf_ram.RAM[2][22] ),
    .X(net2915));
 sg13g2_dlygate4sd3_1 hold682 (.A(\rf_ram.RAM[29][7] ),
    .X(net2916));
 sg13g2_dlygate4sd3_1 hold683 (.A(\rf_ram.RAM[17][2] ),
    .X(net2917));
 sg13g2_dlygate4sd3_1 hold684 (.A(\rf_ram.RAM[9][0] ),
    .X(net2918));
 sg13g2_dlygate4sd3_1 hold685 (.A(_00720_),
    .X(net2919));
 sg13g2_dlygate4sd3_1 hold686 (.A(\rf_ram.RAM[8][28] ),
    .X(net2920));
 sg13g2_dlygate4sd3_1 hold687 (.A(\rf_ram.RAM[16][23] ),
    .X(net2921));
 sg13g2_dlygate4sd3_1 hold688 (.A(\rf_ram.RAM[30][13] ),
    .X(net2922));
 sg13g2_dlygate4sd3_1 hold689 (.A(\rf_ram.RAM[25][15] ),
    .X(net2923));
 sg13g2_dlygate4sd3_1 hold690 (.A(\rf_ram.RAM[21][12] ),
    .X(net2924));
 sg13g2_dlygate4sd3_1 hold691 (.A(\rf_ram.RAM[11][29] ),
    .X(net2925));
 sg13g2_dlygate4sd3_1 hold692 (.A(\rf_ram.RAM[19][16] ),
    .X(net2926));
 sg13g2_dlygate4sd3_1 hold693 (.A(\rf_ram.RAM[5][11] ),
    .X(net2927));
 sg13g2_dlygate4sd3_1 hold694 (.A(\rf_ram.RAM[15][19] ),
    .X(net2928));
 sg13g2_dlygate4sd3_1 hold695 (.A(\rf_ram.RAM[5][2] ),
    .X(net2929));
 sg13g2_dlygate4sd3_1 hold696 (.A(\rf_ram.RAM[19][8] ),
    .X(net2930));
 sg13g2_dlygate4sd3_1 hold697 (.A(\rf_ram.RAM[0][22] ),
    .X(net2931));
 sg13g2_dlygate4sd3_1 hold698 (.A(\rf_ram.RAM[23][26] ),
    .X(net2932));
 sg13g2_dlygate4sd3_1 hold699 (.A(\rf_ram.RAM[31][13] ),
    .X(net2933));
 sg13g2_dlygate4sd3_1 hold700 (.A(\rf_ram.RAM[9][3] ),
    .X(net2934));
 sg13g2_dlygate4sd3_1 hold701 (.A(\rf_ram.RAM[28][20] ),
    .X(net2935));
 sg13g2_dlygate4sd3_1 hold702 (.A(\rf_ram.RAM[28][4] ),
    .X(net2936));
 sg13g2_dlygate4sd3_1 hold703 (.A(\rf_ram.RAM[12][26] ),
    .X(net2937));
 sg13g2_dlygate4sd3_1 hold704 (.A(\rf_ram.RAM[5][30] ),
    .X(net2938));
 sg13g2_dlygate4sd3_1 hold705 (.A(\rf_ram.RAM[31][29] ),
    .X(net2939));
 sg13g2_dlygate4sd3_1 hold706 (.A(\rf_ram.RAM[12][24] ),
    .X(net2940));
 sg13g2_dlygate4sd3_1 hold707 (.A(\rf_ram.RAM[1][19] ),
    .X(net2941));
 sg13g2_dlygate4sd3_1 hold708 (.A(\rf_ram.RAM[4][10] ),
    .X(net2942));
 sg13g2_dlygate4sd3_1 hold709 (.A(\rf_ram.RAM[11][26] ),
    .X(net2943));
 sg13g2_dlygate4sd3_1 hold710 (.A(\rf_ram.RAM[15][14] ),
    .X(net2944));
 sg13g2_dlygate4sd3_1 hold711 (.A(\rf_ram.RAM[22][10] ),
    .X(net2945));
 sg13g2_dlygate4sd3_1 hold712 (.A(\rf_ram.RAM[16][12] ),
    .X(net2946));
 sg13g2_dlygate4sd3_1 hold713 (.A(\rf_ram.RAM[16][11] ),
    .X(net2947));
 sg13g2_dlygate4sd3_1 hold714 (.A(\rf_ram.RAM[17][11] ),
    .X(net2948));
 sg13g2_dlygate4sd3_1 hold715 (.A(\rf_ram.RAM[3][8] ),
    .X(net2949));
 sg13g2_dlygate4sd3_1 hold716 (.A(\rf_ram.RAM[0][25] ),
    .X(net2950));
 sg13g2_dlygate4sd3_1 hold717 (.A(\rf_ram.RAM[5][21] ),
    .X(net2951));
 sg13g2_dlygate4sd3_1 hold718 (.A(\rf_ram.RAM[29][13] ),
    .X(net2952));
 sg13g2_dlygate4sd3_1 hold719 (.A(\rf_ram.RAM[4][8] ),
    .X(net2953));
 sg13g2_dlygate4sd3_1 hold720 (.A(\rf_ram.RAM[24][12] ),
    .X(net2954));
 sg13g2_dlygate4sd3_1 hold721 (.A(\rf_ram.RAM[14][8] ),
    .X(net2955));
 sg13g2_dlygate4sd3_1 hold722 (.A(\rf_ram.RAM[13][13] ),
    .X(net2956));
 sg13g2_dlygate4sd3_1 hold723 (.A(\rf_ram.RAM[4][29] ),
    .X(net2957));
 sg13g2_dlygate4sd3_1 hold724 (.A(\rf_ram.RAM[19][3] ),
    .X(net2958));
 sg13g2_dlygate4sd3_1 hold725 (.A(\rf_ram.RAM[28][10] ),
    .X(net2959));
 sg13g2_dlygate4sd3_1 hold726 (.A(\rf_ram.RAM[26][9] ),
    .X(net2960));
 sg13g2_dlygate4sd3_1 hold727 (.A(\rf_ram.RAM[27][4] ),
    .X(net2961));
 sg13g2_dlygate4sd3_1 hold728 (.A(\rf_ram.RAM[19][15] ),
    .X(net2962));
 sg13g2_dlygate4sd3_1 hold729 (.A(\rf_ram.RAM[23][1] ),
    .X(net2963));
 sg13g2_dlygate4sd3_1 hold730 (.A(\rf_ram.RAM[13][26] ),
    .X(net2964));
 sg13g2_dlygate4sd3_1 hold731 (.A(\rf_ram.RAM[5][7] ),
    .X(net2965));
 sg13g2_dlygate4sd3_1 hold732 (.A(\rf_ram.RAM[21][28] ),
    .X(net2966));
 sg13g2_dlygate4sd3_1 hold733 (.A(\rf_ram.RAM[29][27] ),
    .X(net2967));
 sg13g2_dlygate4sd3_1 hold734 (.A(\rf_ram.RAM[18][5] ),
    .X(net2968));
 sg13g2_dlygate4sd3_1 hold735 (.A(\rf_ram.RAM[16][4] ),
    .X(net2969));
 sg13g2_dlygate4sd3_1 hold736 (.A(\rf_ram.RAM[8][17] ),
    .X(net2970));
 sg13g2_dlygate4sd3_1 hold737 (.A(\rf_ram.RAM[25][29] ),
    .X(net2971));
 sg13g2_dlygate4sd3_1 hold738 (.A(\rf_ram.RAM[16][22] ),
    .X(net2972));
 sg13g2_dlygate4sd3_1 hold739 (.A(\rf_ram.RAM[26][10] ),
    .X(net2973));
 sg13g2_dlygate4sd3_1 hold740 (.A(\rf_ram.RAM[26][25] ),
    .X(net2974));
 sg13g2_dlygate4sd3_1 hold741 (.A(\rf_ram.RAM[11][31] ),
    .X(net2975));
 sg13g2_dlygate4sd3_1 hold742 (.A(\rf_ram.RAM[10][20] ),
    .X(net2976));
 sg13g2_dlygate4sd3_1 hold743 (.A(\rf_ram.RAM[24][28] ),
    .X(net2977));
 sg13g2_dlygate4sd3_1 hold744 (.A(\rf_ram.RAM[8][19] ),
    .X(net2978));
 sg13g2_dlygate4sd3_1 hold745 (.A(\rf_ram.RAM[20][20] ),
    .X(net2979));
 sg13g2_dlygate4sd3_1 hold746 (.A(\rf_ram.RAM[25][17] ),
    .X(net2980));
 sg13g2_dlygate4sd3_1 hold747 (.A(\rf_ram.RAM[12][2] ),
    .X(net2981));
 sg13g2_dlygate4sd3_1 hold748 (.A(\rf_ram.RAM[7][7] ),
    .X(net2982));
 sg13g2_dlygate4sd3_1 hold749 (.A(\rf_ram.RAM[12][18] ),
    .X(net2983));
 sg13g2_dlygate4sd3_1 hold750 (.A(\rf_ram.RAM[19][26] ),
    .X(net2984));
 sg13g2_dlygate4sd3_1 hold751 (.A(\rf_ram.RAM[1][28] ),
    .X(net2985));
 sg13g2_dlygate4sd3_1 hold752 (.A(\rf_ram.RAM[18][25] ),
    .X(net2986));
 sg13g2_dlygate4sd3_1 hold753 (.A(\rf_ram.RAM[25][11] ),
    .X(net2987));
 sg13g2_dlygate4sd3_1 hold754 (.A(\rf_ram.RAM[27][6] ),
    .X(net2988));
 sg13g2_dlygate4sd3_1 hold755 (.A(\rf_ram.RAM[11][17] ),
    .X(net2989));
 sg13g2_dlygate4sd3_1 hold756 (.A(\rf_ram.RAM[15][31] ),
    .X(net2990));
 sg13g2_dlygate4sd3_1 hold757 (.A(\rf_ram.RAM[29][10] ),
    .X(net2991));
 sg13g2_dlygate4sd3_1 hold758 (.A(\rf_ram.RAM[24][5] ),
    .X(net2992));
 sg13g2_dlygate4sd3_1 hold759 (.A(\cpu.cpu.mem_if.signbit ),
    .X(net2993));
 sg13g2_dlygate4sd3_1 hold760 (.A(_01517_),
    .X(net2994));
 sg13g2_dlygate4sd3_1 hold761 (.A(_00473_),
    .X(net2995));
 sg13g2_dlygate4sd3_1 hold762 (.A(\rf_ram.RAM[23][5] ),
    .X(net2996));
 sg13g2_dlygate4sd3_1 hold763 (.A(\rf_ram.RAM[25][16] ),
    .X(net2997));
 sg13g2_dlygate4sd3_1 hold764 (.A(\rf_ram.RAM[8][9] ),
    .X(net2998));
 sg13g2_dlygate4sd3_1 hold765 (.A(\rf_ram.RAM[15][4] ),
    .X(net2999));
 sg13g2_dlygate4sd3_1 hold766 (.A(\rf_ram.RAM[26][19] ),
    .X(net3000));
 sg13g2_dlygate4sd3_1 hold767 (.A(\rf_ram.RAM[6][20] ),
    .X(net3001));
 sg13g2_dlygate4sd3_1 hold768 (.A(\rf_ram.RAM[16][17] ),
    .X(net3002));
 sg13g2_dlygate4sd3_1 hold769 (.A(\rf_ram.RAM[24][17] ),
    .X(net3003));
 sg13g2_dlygate4sd3_1 hold770 (.A(\rf_ram.RAM[7][30] ),
    .X(net3004));
 sg13g2_dlygate4sd3_1 hold771 (.A(\rf_ram.RAM[21][1] ),
    .X(net3005));
 sg13g2_dlygate4sd3_1 hold772 (.A(\rf_ram.RAM[5][23] ),
    .X(net3006));
 sg13g2_dlygate4sd3_1 hold773 (.A(\rf_ram.RAM[15][28] ),
    .X(net3007));
 sg13g2_dlygate4sd3_1 hold774 (.A(\rf_ram.RAM[17][12] ),
    .X(net3008));
 sg13g2_dlygate4sd3_1 hold775 (.A(\rf_ram.RAM[16][19] ),
    .X(net3009));
 sg13g2_dlygate4sd3_1 hold776 (.A(\rf_ram.RAM[25][14] ),
    .X(net3010));
 sg13g2_dlygate4sd3_1 hold777 (.A(\rf_ram.RAM[8][2] ),
    .X(net3011));
 sg13g2_dlygate4sd3_1 hold778 (.A(\rf_ram.RAM[29][19] ),
    .X(net3012));
 sg13g2_dlygate4sd3_1 hold779 (.A(\rf_ram.RAM[31][20] ),
    .X(net3013));
 sg13g2_dlygate4sd3_1 hold780 (.A(\rf_ram.RAM[7][27] ),
    .X(net3014));
 sg13g2_dlygate4sd3_1 hold781 (.A(\rf_ram.RAM[3][14] ),
    .X(net3015));
 sg13g2_dlygate4sd3_1 hold782 (.A(\rf_ram.RAM[26][27] ),
    .X(net3016));
 sg13g2_dlygate4sd3_1 hold783 (.A(\rf_ram.RAM[30][21] ),
    .X(net3017));
 sg13g2_dlygate4sd3_1 hold784 (.A(\rf_ram.RAM[7][13] ),
    .X(net3018));
 sg13g2_dlygate4sd3_1 hold785 (.A(\rf_ram.RAM[11][2] ),
    .X(net3019));
 sg13g2_dlygate4sd3_1 hold786 (.A(\rf_ram.RAM[7][26] ),
    .X(net3020));
 sg13g2_dlygate4sd3_1 hold787 (.A(\rf_ram.RAM[11][0] ),
    .X(net3021));
 sg13g2_dlygate4sd3_1 hold788 (.A(_01188_),
    .X(net3022));
 sg13g2_dlygate4sd3_1 hold789 (.A(\rf_ram.RAM[15][25] ),
    .X(net3023));
 sg13g2_dlygate4sd3_1 hold790 (.A(\rf_ram.RAM[12][22] ),
    .X(net3024));
 sg13g2_dlygate4sd3_1 hold791 (.A(\rf_ram.RAM[23][21] ),
    .X(net3025));
 sg13g2_dlygate4sd3_1 hold792 (.A(\rf_ram.RAM[25][25] ),
    .X(net3026));
 sg13g2_dlygate4sd3_1 hold793 (.A(\rf_ram.RAM[20][22] ),
    .X(net3027));
 sg13g2_dlygate4sd3_1 hold794 (.A(\rf_ram.RAM[13][5] ),
    .X(net3028));
 sg13g2_dlygate4sd3_1 hold795 (.A(\rf_ram.RAM[19][31] ),
    .X(net3029));
 sg13g2_dlygate4sd3_1 hold796 (.A(\rf_ram.RAM[13][21] ),
    .X(net3030));
 sg13g2_dlygate4sd3_1 hold797 (.A(\rf_ram.RAM[0][26] ),
    .X(net3031));
 sg13g2_dlygate4sd3_1 hold798 (.A(\rf_ram.RAM[3][0] ),
    .X(net3032));
 sg13g2_dlygate4sd3_1 hold799 (.A(_00620_),
    .X(net3033));
 sg13g2_dlygate4sd3_1 hold800 (.A(\rf_ram.RAM[6][29] ),
    .X(net3034));
 sg13g2_dlygate4sd3_1 hold801 (.A(\rf_ram.RAM[10][23] ),
    .X(net3035));
 sg13g2_dlygate4sd3_1 hold802 (.A(\rf_ram.RAM[3][4] ),
    .X(net3036));
 sg13g2_dlygate4sd3_1 hold803 (.A(\rf_ram.RAM[3][23] ),
    .X(net3037));
 sg13g2_dlygate4sd3_1 hold804 (.A(\rf_ram.RAM[21][17] ),
    .X(net3038));
 sg13g2_dlygate4sd3_1 hold805 (.A(\rf_ram.RAM[3][30] ),
    .X(net3039));
 sg13g2_dlygate4sd3_1 hold806 (.A(\rf_ram.RAM[22][11] ),
    .X(net3040));
 sg13g2_dlygate4sd3_1 hold807 (.A(\rf_ram.RAM[5][31] ),
    .X(net3041));
 sg13g2_dlygate4sd3_1 hold808 (.A(\rf_ram.RAM[24][9] ),
    .X(net3042));
 sg13g2_dlygate4sd3_1 hold809 (.A(\rf_ram.RAM[10][8] ),
    .X(net3043));
 sg13g2_dlygate4sd3_1 hold810 (.A(\rf_ram.RAM[4][11] ),
    .X(net3044));
 sg13g2_dlygate4sd3_1 hold811 (.A(\rf_ram.RAM[1][2] ),
    .X(net3045));
 sg13g2_dlygate4sd3_1 hold812 (.A(\rf_ram.RAM[16][14] ),
    .X(net3046));
 sg13g2_dlygate4sd3_1 hold813 (.A(\rf_ram.RAM[15][11] ),
    .X(net3047));
 sg13g2_dlygate4sd3_1 hold814 (.A(\rf_ram.RAM[27][27] ),
    .X(net3048));
 sg13g2_dlygate4sd3_1 hold815 (.A(\rf_ram.RAM[9][2] ),
    .X(net3049));
 sg13g2_dlygate4sd3_1 hold816 (.A(\rf_ram.RAM[26][16] ),
    .X(net3050));
 sg13g2_dlygate4sd3_1 hold817 (.A(\rf_ram.RAM[22][31] ),
    .X(net3051));
 sg13g2_dlygate4sd3_1 hold818 (.A(\rf_ram.RAM[1][23] ),
    .X(net3052));
 sg13g2_dlygate4sd3_1 hold819 (.A(\rf_ram.RAM[19][29] ),
    .X(net3053));
 sg13g2_dlygate4sd3_1 hold820 (.A(\rf_ram.RAM[20][6] ),
    .X(net3054));
 sg13g2_dlygate4sd3_1 hold821 (.A(\rf_ram.RAM[6][2] ),
    .X(net3055));
 sg13g2_dlygate4sd3_1 hold822 (.A(\rf_ram.RAM[10][11] ),
    .X(net3056));
 sg13g2_dlygate4sd3_1 hold823 (.A(\rf_ram.RAM[2][24] ),
    .X(net3057));
 sg13g2_dlygate4sd3_1 hold824 (.A(\rf_ram.RAM[24][26] ),
    .X(net3058));
 sg13g2_dlygate4sd3_1 hold825 (.A(\rf_ram.RAM[2][15] ),
    .X(net3059));
 sg13g2_dlygate4sd3_1 hold826 (.A(\rf_ram.RAM[12][1] ),
    .X(net3060));
 sg13g2_dlygate4sd3_1 hold827 (.A(\rf_ram.RAM[26][8] ),
    .X(net3061));
 sg13g2_dlygate4sd3_1 hold828 (.A(\rf_ram.RAM[9][19] ),
    .X(net3062));
 sg13g2_dlygate4sd3_1 hold829 (.A(\rf_ram.RAM[21][11] ),
    .X(net3063));
 sg13g2_dlygate4sd3_1 hold830 (.A(\rf_ram.RAM[6][1] ),
    .X(net3064));
 sg13g2_dlygate4sd3_1 hold831 (.A(\rf_ram.RAM[10][29] ),
    .X(net3065));
 sg13g2_dlygate4sd3_1 hold832 (.A(\rf_ram.RAM[21][29] ),
    .X(net3066));
 sg13g2_dlygate4sd3_1 hold833 (.A(\rf_ram.RAM[21][5] ),
    .X(net3067));
 sg13g2_dlygate4sd3_1 hold834 (.A(\rf_ram.RAM[22][21] ),
    .X(net3068));
 sg13g2_dlygate4sd3_1 hold835 (.A(\rf_ram.RAM[5][8] ),
    .X(net3069));
 sg13g2_dlygate4sd3_1 hold836 (.A(\rf_ram.RAM[15][13] ),
    .X(net3070));
 sg13g2_dlygate4sd3_1 hold837 (.A(\rf_ram.RAM[0][14] ),
    .X(net3071));
 sg13g2_dlygate4sd3_1 hold838 (.A(\rf_ram.RAM[13][25] ),
    .X(net3072));
 sg13g2_dlygate4sd3_1 hold839 (.A(\rf_ram.RAM[7][8] ),
    .X(net3073));
 sg13g2_dlygate4sd3_1 hold840 (.A(\rf_ram.RAM[12][20] ),
    .X(net3074));
 sg13g2_dlygate4sd3_1 hold841 (.A(\rf_ram.RAM[12][7] ),
    .X(net3075));
 sg13g2_dlygate4sd3_1 hold842 (.A(\rf_ram.RAM[19][30] ),
    .X(net3076));
 sg13g2_dlygate4sd3_1 hold843 (.A(\rf_ram.RAM[16][28] ),
    .X(net3077));
 sg13g2_dlygate4sd3_1 hold844 (.A(\rf_ram.RAM[20][25] ),
    .X(net3078));
 sg13g2_dlygate4sd3_1 hold845 (.A(\rf_ram.RAM[27][16] ),
    .X(net3079));
 sg13g2_dlygate4sd3_1 hold846 (.A(\rf_ram.RAM[29][3] ),
    .X(net3080));
 sg13g2_dlygate4sd3_1 hold847 (.A(\rf_ram.RAM[1][14] ),
    .X(net3081));
 sg13g2_dlygate4sd3_1 hold848 (.A(\rf_ram.RAM[22][20] ),
    .X(net3082));
 sg13g2_dlygate4sd3_1 hold849 (.A(\rf_ram.RAM[12][3] ),
    .X(net3083));
 sg13g2_dlygate4sd3_1 hold850 (.A(\rf_ram.RAM[22][14] ),
    .X(net3084));
 sg13g2_dlygate4sd3_1 hold851 (.A(\rf_ram.RAM[10][13] ),
    .X(net3085));
 sg13g2_dlygate4sd3_1 hold852 (.A(\rf_ram.RAM[14][26] ),
    .X(net3086));
 sg13g2_dlygate4sd3_1 hold853 (.A(\rf_ram.RAM[10][3] ),
    .X(net3087));
 sg13g2_dlygate4sd3_1 hold854 (.A(\rf_ram.RAM[17][30] ),
    .X(net3088));
 sg13g2_dlygate4sd3_1 hold855 (.A(\rf_ram.RAM[15][27] ),
    .X(net3089));
 sg13g2_dlygate4sd3_1 hold856 (.A(\rf_ram.RAM[3][26] ),
    .X(net3090));
 sg13g2_dlygate4sd3_1 hold857 (.A(\rf_ram.RAM[28][15] ),
    .X(net3091));
 sg13g2_dlygate4sd3_1 hold858 (.A(\rf_ram.RAM[25][2] ),
    .X(net3092));
 sg13g2_dlygate4sd3_1 hold859 (.A(\rf_ram.RAM[31][1] ),
    .X(net3093));
 sg13g2_dlygate4sd3_1 hold860 (.A(\rf_ram.RAM[24][13] ),
    .X(net3094));
 sg13g2_dlygate4sd3_1 hold861 (.A(\rf_ram.RAM[30][30] ),
    .X(net3095));
 sg13g2_dlygate4sd3_1 hold862 (.A(\rf_ram.RAM[13][2] ),
    .X(net3096));
 sg13g2_dlygate4sd3_1 hold863 (.A(\rf_ram.RAM[25][28] ),
    .X(net3097));
 sg13g2_dlygate4sd3_1 hold864 (.A(\rf_ram.RAM[1][26] ),
    .X(net3098));
 sg13g2_dlygate4sd3_1 hold865 (.A(\rf_ram.RAM[15][8] ),
    .X(net3099));
 sg13g2_dlygate4sd3_1 hold866 (.A(\rf_ram.RAM[5][28] ),
    .X(net3100));
 sg13g2_dlygate4sd3_1 hold867 (.A(\rf_ram.RAM[27][7] ),
    .X(net3101));
 sg13g2_dlygate4sd3_1 hold868 (.A(\rf_ram.RAM[23][14] ),
    .X(net3102));
 sg13g2_dlygate4sd3_1 hold869 (.A(\rf_ram.RAM[23][13] ),
    .X(net3103));
 sg13g2_dlygate4sd3_1 hold870 (.A(\rf_ram.RAM[30][29] ),
    .X(net3104));
 sg13g2_dlygate4sd3_1 hold871 (.A(\rf_ram.RAM[18][23] ),
    .X(net3105));
 sg13g2_dlygate4sd3_1 hold872 (.A(\rf_ram.RAM[13][24] ),
    .X(net3106));
 sg13g2_dlygate4sd3_1 hold873 (.A(\rf_ram.RAM[18][17] ),
    .X(net3107));
 sg13g2_dlygate4sd3_1 hold874 (.A(\rf_ram.RAM[21][9] ),
    .X(net3108));
 sg13g2_dlygate4sd3_1 hold875 (.A(\rf_ram.RAM[1][11] ),
    .X(net3109));
 sg13g2_dlygate4sd3_1 hold876 (.A(\rf_ram.RAM[19][28] ),
    .X(net3110));
 sg13g2_dlygate4sd3_1 hold877 (.A(\rf_ram.RAM[29][30] ),
    .X(net3111));
 sg13g2_dlygate4sd3_1 hold878 (.A(\rf_ram.RAM[19][6] ),
    .X(net3112));
 sg13g2_dlygate4sd3_1 hold879 (.A(\rf_ram.RAM[4][23] ),
    .X(net3113));
 sg13g2_dlygate4sd3_1 hold880 (.A(\rf_ram.RAM[5][29] ),
    .X(net3114));
 sg13g2_dlygate4sd3_1 hold881 (.A(\rf_ram.RAM[29][26] ),
    .X(net3115));
 sg13g2_dlygate4sd3_1 hold882 (.A(\rf_ram.RAM[29][31] ),
    .X(net3116));
 sg13g2_dlygate4sd3_1 hold883 (.A(\rf_ram.RAM[27][13] ),
    .X(net3117));
 sg13g2_dlygate4sd3_1 hold884 (.A(\rf_ram.RAM[18][20] ),
    .X(net3118));
 sg13g2_dlygate4sd3_1 hold885 (.A(\rf_ram.RAM[8][13] ),
    .X(net3119));
 sg13g2_dlygate4sd3_1 hold886 (.A(\rf_ram.RAM[20][27] ),
    .X(net3120));
 sg13g2_dlygate4sd3_1 hold887 (.A(\rf_ram.RAM[3][1] ),
    .X(net3121));
 sg13g2_dlygate4sd3_1 hold888 (.A(\rf_ram.RAM[27][8] ),
    .X(net3122));
 sg13g2_dlygate4sd3_1 hold889 (.A(\rf_ram.RAM[3][22] ),
    .X(net3123));
 sg13g2_dlygate4sd3_1 hold890 (.A(\rf_ram.RAM[20][23] ),
    .X(net3124));
 sg13g2_dlygate4sd3_1 hold891 (.A(\rf_ram.RAM[15][18] ),
    .X(net3125));
 sg13g2_dlygate4sd3_1 hold892 (.A(\rf_ram.RAM[13][31] ),
    .X(net3126));
 sg13g2_dlygate4sd3_1 hold893 (.A(\rf_ram.RAM[29][2] ),
    .X(net3127));
 sg13g2_dlygate4sd3_1 hold894 (.A(\rf_ram.RAM[17][1] ),
    .X(net3128));
 sg13g2_dlygate4sd3_1 hold895 (.A(\rf_ram.RAM[28][16] ),
    .X(net3129));
 sg13g2_dlygate4sd3_1 hold896 (.A(\rf_ram.RAM[31][31] ),
    .X(net3130));
 sg13g2_dlygate4sd3_1 hold897 (.A(\rf_ram.RAM[22][30] ),
    .X(net3131));
 sg13g2_dlygate4sd3_1 hold898 (.A(\rf_ram.RAM[6][7] ),
    .X(net3132));
 sg13g2_dlygate4sd3_1 hold899 (.A(\rf_ram.RAM[20][3] ),
    .X(net3133));
 sg13g2_dlygate4sd3_1 hold900 (.A(\rf_ram.RAM[9][16] ),
    .X(net3134));
 sg13g2_dlygate4sd3_1 hold901 (.A(\rf_ram.RAM[5][15] ),
    .X(net3135));
 sg13g2_dlygate4sd3_1 hold902 (.A(\rf_ram.RAM[9][14] ),
    .X(net3136));
 sg13g2_dlygate4sd3_1 hold903 (.A(\rf_ram.RAM[31][10] ),
    .X(net3137));
 sg13g2_dlygate4sd3_1 hold904 (.A(\rf_ram.RAM[17][18] ),
    .X(net3138));
 sg13g2_dlygate4sd3_1 hold905 (.A(\rf_ram.RAM[31][12] ),
    .X(net3139));
 sg13g2_dlygate4sd3_1 hold906 (.A(\rf_ram.RAM[10][16] ),
    .X(net3140));
 sg13g2_dlygate4sd3_1 hold907 (.A(\rf_ram.RAM[0][15] ),
    .X(net3141));
 sg13g2_dlygate4sd3_1 hold908 (.A(\rf_ram.RAM[5][0] ),
    .X(net3142));
 sg13g2_dlygate4sd3_1 hold909 (.A(_00916_),
    .X(net3143));
 sg13g2_dlygate4sd3_1 hold910 (.A(\rf_ram.RAM[10][0] ),
    .X(net3144));
 sg13g2_dlygate4sd3_1 hold911 (.A(_00550_),
    .X(net3145));
 sg13g2_dlygate4sd3_1 hold912 (.A(\rf_ram.RAM[4][7] ),
    .X(net3146));
 sg13g2_dlygate4sd3_1 hold913 (.A(\rf_ram.RAM[29][9] ),
    .X(net3147));
 sg13g2_dlygate4sd3_1 hold914 (.A(\rf_ram.RAM[25][13] ),
    .X(net3148));
 sg13g2_dlygate4sd3_1 hold915 (.A(\rf_ram.RAM[21][10] ),
    .X(net3149));
 sg13g2_dlygate4sd3_1 hold916 (.A(\rf_ram.RAM[12][13] ),
    .X(net3150));
 sg13g2_dlygate4sd3_1 hold917 (.A(\rf_ram.RAM[19][14] ),
    .X(net3151));
 sg13g2_dlygate4sd3_1 hold918 (.A(\rf_ram.RAM[21][3] ),
    .X(net3152));
 sg13g2_dlygate4sd3_1 hold919 (.A(\rf_ram.RAM[31][3] ),
    .X(net3153));
 sg13g2_dlygate4sd3_1 hold920 (.A(\rf_ram.RAM[15][20] ),
    .X(net3154));
 sg13g2_dlygate4sd3_1 hold921 (.A(\rf_ram.RAM[30][1] ),
    .X(net3155));
 sg13g2_dlygate4sd3_1 hold922 (.A(\rf_ram.RAM[15][0] ),
    .X(net3156));
 sg13g2_dlygate4sd3_1 hold923 (.A(_00688_),
    .X(net3157));
 sg13g2_dlygate4sd3_1 hold924 (.A(\rf_ram.RAM[3][19] ),
    .X(net3158));
 sg13g2_dlygate4sd3_1 hold925 (.A(\rf_ram.RAM[23][24] ),
    .X(net3159));
 sg13g2_dlygate4sd3_1 hold926 (.A(\rf_ram.RAM[2][12] ),
    .X(net3160));
 sg13g2_dlygate4sd3_1 hold927 (.A(\rf_ram.RAM[20][26] ),
    .X(net3161));
 sg13g2_dlygate4sd3_1 hold928 (.A(\rf_ram.RAM[6][16] ),
    .X(net3162));
 sg13g2_dlygate4sd3_1 hold929 (.A(\rf_ram.RAM[7][1] ),
    .X(net3163));
 sg13g2_dlygate4sd3_1 hold930 (.A(\rf_ram.RAM[3][31] ),
    .X(net3164));
 sg13g2_dlygate4sd3_1 hold931 (.A(\rf_ram.RAM[3][12] ),
    .X(net3165));
 sg13g2_dlygate4sd3_1 hold932 (.A(\rf_ram.RAM[29][16] ),
    .X(net3166));
 sg13g2_dlygate4sd3_1 hold933 (.A(\rf_ram.RAM[9][21] ),
    .X(net3167));
 sg13g2_dlygate4sd3_1 hold934 (.A(\rf_ram.RAM[9][12] ),
    .X(net3168));
 sg13g2_dlygate4sd3_1 hold935 (.A(\rf_ram.RAM[4][6] ),
    .X(net3169));
 sg13g2_dlygate4sd3_1 hold936 (.A(\rf_ram.RAM[0][11] ),
    .X(net3170));
 sg13g2_dlygate4sd3_1 hold937 (.A(\rf_ram.RAM[8][15] ),
    .X(net3171));
 sg13g2_dlygate4sd3_1 hold938 (.A(\rf_ram.RAM[1][31] ),
    .X(net3172));
 sg13g2_dlygate4sd3_1 hold939 (.A(\rf_ram.RAM[18][7] ),
    .X(net3173));
 sg13g2_dlygate4sd3_1 hold940 (.A(\rf_ram.RAM[11][11] ),
    .X(net3174));
 sg13g2_dlygate4sd3_1 hold941 (.A(\rf_ram.RAM[22][1] ),
    .X(net3175));
 sg13g2_dlygate4sd3_1 hold942 (.A(\rf_ram.RAM[26][24] ),
    .X(net3176));
 sg13g2_dlygate4sd3_1 hold943 (.A(\rf_ram.RAM[21][21] ),
    .X(net3177));
 sg13g2_dlygate4sd3_1 hold944 (.A(\rf_ram.RAM[1][18] ),
    .X(net3178));
 sg13g2_dlygate4sd3_1 hold945 (.A(\rf_ram.RAM[14][17] ),
    .X(net3179));
 sg13g2_dlygate4sd3_1 hold946 (.A(\rf_ram.RAM[1][7] ),
    .X(net3180));
 sg13g2_dlygate4sd3_1 hold947 (.A(\rf_ram.RAM[20][16] ),
    .X(net3181));
 sg13g2_dlygate4sd3_1 hold948 (.A(\rf_ram.RAM[15][15] ),
    .X(net3182));
 sg13g2_dlygate4sd3_1 hold949 (.A(\rf_ram.RAM[11][28] ),
    .X(net3183));
 sg13g2_dlygate4sd3_1 hold950 (.A(\rf_ram.RAM[22][3] ),
    .X(net3184));
 sg13g2_dlygate4sd3_1 hold951 (.A(\rf_ram.RAM[2][2] ),
    .X(net3185));
 sg13g2_dlygate4sd3_1 hold952 (.A(\rf_ram.RAM[6][12] ),
    .X(net3186));
 sg13g2_dlygate4sd3_1 hold953 (.A(\rf_ram.RAM[23][8] ),
    .X(net3187));
 sg13g2_dlygate4sd3_1 hold954 (.A(\rf_ram.RAM[28][9] ),
    .X(net3188));
 sg13g2_dlygate4sd3_1 hold955 (.A(\rf_ram.RAM[25][27] ),
    .X(net3189));
 sg13g2_dlygate4sd3_1 hold956 (.A(\rf_ram.RAM[2][16] ),
    .X(net3190));
 sg13g2_dlygate4sd3_1 hold957 (.A(\rf_ram.RAM[1][15] ),
    .X(net3191));
 sg13g2_dlygate4sd3_1 hold958 (.A(\rf_ram.RAM[30][12] ),
    .X(net3192));
 sg13g2_dlygate4sd3_1 hold959 (.A(\rf_ram.RAM[24][25] ),
    .X(net3193));
 sg13g2_dlygate4sd3_1 hold960 (.A(\rf_ram.RAM[8][21] ),
    .X(net3194));
 sg13g2_dlygate4sd3_1 hold961 (.A(\rf_ram.RAM[23][18] ),
    .X(net3195));
 sg13g2_dlygate4sd3_1 hold962 (.A(\rf_ram.RAM[1][10] ),
    .X(net3196));
 sg13g2_dlygate4sd3_1 hold963 (.A(\rf_ram.RAM[30][0] ),
    .X(net3197));
 sg13g2_dlygate4sd3_1 hold964 (.A(_00980_),
    .X(net3198));
 sg13g2_dlygate4sd3_1 hold965 (.A(\rf_ram.RAM[28][13] ),
    .X(net3199));
 sg13g2_dlygate4sd3_1 hold966 (.A(\rf_ram.RAM[20][13] ),
    .X(net3200));
 sg13g2_dlygate4sd3_1 hold967 (.A(\rf_ram.RAM[27][14] ),
    .X(net3201));
 sg13g2_dlygate4sd3_1 hold968 (.A(\rf_ram.RAM[27][0] ),
    .X(net3202));
 sg13g2_dlygate4sd3_1 hold969 (.A(\rf_ram.RAM[28][8] ),
    .X(net3203));
 sg13g2_dlygate4sd3_1 hold970 (.A(\rf_ram.RAM[28][24] ),
    .X(net3204));
 sg13g2_dlygate4sd3_1 hold971 (.A(\rf_ram.RAM[2][26] ),
    .X(net3205));
 sg13g2_dlygate4sd3_1 hold972 (.A(\rf_ram.RAM[11][3] ),
    .X(net3206));
 sg13g2_dlygate4sd3_1 hold973 (.A(\rf_ram.RAM[27][5] ),
    .X(net3207));
 sg13g2_dlygate4sd3_1 hold974 (.A(\rf_ram.RAM[9][25] ),
    .X(net3208));
 sg13g2_dlygate4sd3_1 hold975 (.A(\rf_ram.RAM[24][31] ),
    .X(net3209));
 sg13g2_dlygate4sd3_1 hold976 (.A(\rf_ram.RAM[30][22] ),
    .X(net3210));
 sg13g2_dlygate4sd3_1 hold977 (.A(\rf_ram.RAM[3][3] ),
    .X(net3211));
 sg13g2_dlygate4sd3_1 hold978 (.A(\rf_ram.RAM[12][19] ),
    .X(net3212));
 sg13g2_dlygate4sd3_1 hold979 (.A(\rf_ram.RAM[5][13] ),
    .X(net3213));
 sg13g2_dlygate4sd3_1 hold980 (.A(\rf_ram.RAM[9][27] ),
    .X(net3214));
 sg13g2_dlygate4sd3_1 hold981 (.A(\rf_ram.RAM[13][10] ),
    .X(net3215));
 sg13g2_dlygate4sd3_1 hold982 (.A(\rf_ram.RAM[31][17] ),
    .X(net3216));
 sg13g2_dlygate4sd3_1 hold983 (.A(\rf_ram.RAM[23][4] ),
    .X(net3217));
 sg13g2_dlygate4sd3_1 hold984 (.A(\rf_ram.RAM[17][16] ),
    .X(net3218));
 sg13g2_dlygate4sd3_1 hold985 (.A(\rf_ram.RAM[8][22] ),
    .X(net3219));
 sg13g2_dlygate4sd3_1 hold986 (.A(\rf_ram.RAM[25][24] ),
    .X(net3220));
 sg13g2_dlygate4sd3_1 hold987 (.A(\rf_ram.RAM[15][6] ),
    .X(net3221));
 sg13g2_dlygate4sd3_1 hold988 (.A(\rf_ram.RAM[12][9] ),
    .X(net3222));
 sg13g2_dlygate4sd3_1 hold989 (.A(\rf_ram.RAM[1][1] ),
    .X(net3223));
 sg13g2_dlygate4sd3_1 hold990 (.A(\rf_ram.RAM[8][23] ),
    .X(net3224));
 sg13g2_dlygate4sd3_1 hold991 (.A(\rf_ram.RAM[15][1] ),
    .X(net3225));
 sg13g2_dlygate4sd3_1 hold992 (.A(\rf_ram.RAM[18][6] ),
    .X(net3226));
 sg13g2_dlygate4sd3_1 hold993 (.A(\rf_ram.RAM[6][24] ),
    .X(net3227));
 sg13g2_dlygate4sd3_1 hold994 (.A(\rf_ram.RAM[8][27] ),
    .X(net3228));
 sg13g2_dlygate4sd3_1 hold995 (.A(\rf_ram.RAM[2][23] ),
    .X(net3229));
 sg13g2_dlygate4sd3_1 hold996 (.A(\rf_ram.RAM[15][2] ),
    .X(net3230));
 sg13g2_dlygate4sd3_1 hold997 (.A(\rf_ram.RAM[17][20] ),
    .X(net3231));
 sg13g2_dlygate4sd3_1 hold998 (.A(\rf_ram.RAM[20][29] ),
    .X(net3232));
 sg13g2_dlygate4sd3_1 hold999 (.A(\rf_ram.RAM[23][12] ),
    .X(net3233));
 sg13g2_dlygate4sd3_1 hold1000 (.A(\rf_ram.RAM[29][29] ),
    .X(net3234));
 sg13g2_dlygate4sd3_1 hold1001 (.A(\rf_ram.RAM[17][31] ),
    .X(net3235));
 sg13g2_dlygate4sd3_1 hold1002 (.A(\rf_ram.RAM[9][17] ),
    .X(net3236));
 sg13g2_dlygate4sd3_1 hold1003 (.A(\rf_ram.RAM[28][5] ),
    .X(net3237));
 sg13g2_dlygate4sd3_1 hold1004 (.A(\rf_ram.RAM[4][22] ),
    .X(net3238));
 sg13g2_dlygate4sd3_1 hold1005 (.A(\rf_ram.RAM[27][20] ),
    .X(net3239));
 sg13g2_dlygate4sd3_1 hold1006 (.A(\rf_ram.RAM[4][13] ),
    .X(net3240));
 sg13g2_dlygate4sd3_1 hold1007 (.A(\rf_ram.RAM[13][23] ),
    .X(net3241));
 sg13g2_dlygate4sd3_1 hold1008 (.A(\rf_ram.RAM[1][17] ),
    .X(net3242));
 sg13g2_dlygate4sd3_1 hold1009 (.A(\rf_ram.RAM[16][3] ),
    .X(net3243));
 sg13g2_dlygate4sd3_1 hold1010 (.A(\rf_ram.RAM[21][20] ),
    .X(net3244));
 sg13g2_dlygate4sd3_1 hold1011 (.A(\rf_ram.RAM[21][13] ),
    .X(net3245));
 sg13g2_dlygate4sd3_1 hold1012 (.A(\rf_ram.RAM[25][3] ),
    .X(net3246));
 sg13g2_dlygate4sd3_1 hold1013 (.A(\rf_ram.RAM[14][23] ),
    .X(net3247));
 sg13g2_dlygate4sd3_1 hold1014 (.A(\rf_ram.RAM[19][18] ),
    .X(net3248));
 sg13g2_dlygate4sd3_1 hold1015 (.A(\rf_ram.RAM[15][24] ),
    .X(net3249));
 sg13g2_dlygate4sd3_1 hold1016 (.A(\rf_ram.RAM[2][11] ),
    .X(net3250));
 sg13g2_dlygate4sd3_1 hold1017 (.A(\rf_ram.RAM[16][0] ),
    .X(net3251));
 sg13g2_dlygate4sd3_1 hold1018 (.A(\rf_ram.RAM[31][21] ),
    .X(net3252));
 sg13g2_dlygate4sd3_1 hold1019 (.A(\rf_ram.RAM[7][31] ),
    .X(net3253));
 sg13g2_dlygate4sd3_1 hold1020 (.A(\cpu.cpu.immdec.gen_immdec_w_eq_1.imm7 ),
    .X(net3254));
 sg13g2_dlygate4sd3_1 hold1021 (.A(_00527_),
    .X(net3255));
 sg13g2_dlygate4sd3_1 hold1022 (.A(\rf_ram.RAM[20][10] ),
    .X(net3256));
 sg13g2_dlygate4sd3_1 hold1023 (.A(\rf_ram.RAM[23][7] ),
    .X(net3257));
 sg13g2_dlygate4sd3_1 hold1024 (.A(\rf_ram.RAM[31][5] ),
    .X(net3258));
 sg13g2_dlygate4sd3_1 hold1025 (.A(\rf_ram.RAM[12][21] ),
    .X(net3259));
 sg13g2_dlygate4sd3_1 hold1026 (.A(\rf_ram.RAM[17][22] ),
    .X(net3260));
 sg13g2_dlygate4sd3_1 hold1027 (.A(\cpu.rf_ram_if.rcnt[2] ),
    .X(net3261));
 sg13g2_dlygate4sd3_1 hold1028 (.A(_02686_),
    .X(net3262));
 sg13g2_dlygate4sd3_1 hold1029 (.A(_00312_),
    .X(net3263));
 sg13g2_dlygate4sd3_1 hold1030 (.A(\rf_ram.RAM[17][3] ),
    .X(net3264));
 sg13g2_dlygate4sd3_1 hold1031 (.A(\rf_ram.RAM[3][29] ),
    .X(net3265));
 sg13g2_dlygate4sd3_1 hold1032 (.A(\rf_ram.RAM[4][2] ),
    .X(net3266));
 sg13g2_dlygate4sd3_1 hold1033 (.A(\rf_ram.RAM[26][11] ),
    .X(net3267));
 sg13g2_dlygate4sd3_1 hold1034 (.A(\rf_ram.RAM[19][1] ),
    .X(net3268));
 sg13g2_dlygate4sd3_1 hold1035 (.A(\rf_ram.RAM[17][14] ),
    .X(net3269));
 sg13g2_dlygate4sd3_1 hold1036 (.A(\rf_ram.RAM[27][15] ),
    .X(net3270));
 sg13g2_dlygate4sd3_1 hold1037 (.A(\rf_ram.RAM[21][0] ),
    .X(net3271));
 sg13g2_dlygate4sd3_1 hold1038 (.A(_00215_),
    .X(net3272));
 sg13g2_dlygate4sd3_1 hold1039 (.A(uo_out[6]),
    .X(net3273));
 sg13g2_dlygate4sd3_1 hold1040 (.A(\rf_ram.RAM[14][7] ),
    .X(net3274));
 sg13g2_dlygate4sd3_1 hold1041 (.A(\rf_ram.RAM[24][15] ),
    .X(net3275));
 sg13g2_dlygate4sd3_1 hold1042 (.A(\rf_ram.RAM[9][11] ),
    .X(net3276));
 sg13g2_dlygate4sd3_1 hold1043 (.A(\rf_ram.RAM[29][5] ),
    .X(net3277));
 sg13g2_dlygate4sd3_1 hold1044 (.A(\rf_ram.RAM[15][21] ),
    .X(net3278));
 sg13g2_dlygate4sd3_1 hold1045 (.A(\rf_ram.RAM[11][10] ),
    .X(net3279));
 sg13g2_dlygate4sd3_1 hold1046 (.A(\rf_ram.RAM[4][27] ),
    .X(net3280));
 sg13g2_dlygate4sd3_1 hold1047 (.A(\rf_ram.RAM[29][0] ),
    .X(net3281));
 sg13g2_dlygate4sd3_1 hold1048 (.A(_00371_),
    .X(net3282));
 sg13g2_dlygate4sd3_1 hold1049 (.A(\rf_ram.RAM[24][20] ),
    .X(net3283));
 sg13g2_dlygate4sd3_1 hold1050 (.A(uo_out[7]),
    .X(net3284));
 sg13g2_dlygate4sd3_1 hold1051 (.A(\rf_ram.RAM[24][10] ),
    .X(net3285));
 sg13g2_dlygate4sd3_1 hold1052 (.A(\rf_ram.RAM[23][19] ),
    .X(net3286));
 sg13g2_dlygate4sd3_1 hold1053 (.A(\rf_ram.RAM[29][14] ),
    .X(net3287));
 sg13g2_dlygate4sd3_1 hold1054 (.A(\rf_ram.RAM[9][29] ),
    .X(net3288));
 sg13g2_dlygate4sd3_1 hold1055 (.A(\rf_ram.RAM[28][14] ),
    .X(net3289));
 sg13g2_dlygate4sd3_1 hold1056 (.A(\rf_ram.RAM[13][11] ),
    .X(net3290));
 sg13g2_dlygate4sd3_1 hold1057 (.A(\rf_ram.RAM[24][24] ),
    .X(net3291));
 sg13g2_dlygate4sd3_1 hold1058 (.A(\rf_ram.RAM[23][9] ),
    .X(net3292));
 sg13g2_dlygate4sd3_1 hold1059 (.A(\rf_ram.RAM[2][7] ),
    .X(net3293));
 sg13g2_dlygate4sd3_1 hold1060 (.A(\rf_ram.RAM[18][13] ),
    .X(net3294));
 sg13g2_dlygate4sd3_1 hold1061 (.A(\rf_ram.RAM[24][22] ),
    .X(net3295));
 sg13g2_dlygate4sd3_1 hold1062 (.A(\rf_ram.RAM[25][21] ),
    .X(net3296));
 sg13g2_dlygate4sd3_1 hold1063 (.A(\rf_ram.RAM[18][22] ),
    .X(net3297));
 sg13g2_dlygate4sd3_1 hold1064 (.A(\rf_ram.RAM[3][17] ),
    .X(net3298));
 sg13g2_dlygate4sd3_1 hold1065 (.A(\rf_ram.RAM[27][2] ),
    .X(net3299));
 sg13g2_dlygate4sd3_1 hold1066 (.A(\rf_ram.RAM[25][20] ),
    .X(net3300));
 sg13g2_dlygate4sd3_1 hold1067 (.A(\rf_ram.RAM[25][23] ),
    .X(net3301));
 sg13g2_dlygate4sd3_1 hold1068 (.A(\rf_ram.RAM[27][22] ),
    .X(net3302));
 sg13g2_dlygate4sd3_1 hold1069 (.A(\rf_ram.RAM[2][1] ),
    .X(net3303));
 sg13g2_dlygate4sd3_1 hold1070 (.A(\cpu.rf_ram_if.rdata1[21] ),
    .X(net3304));
 sg13g2_dlygate4sd3_1 hold1071 (.A(_00043_),
    .X(net3305));
 sg13g2_dlygate4sd3_1 hold1072 (.A(\rf_ram.RAM[23][20] ),
    .X(net3306));
 sg13g2_dlygate4sd3_1 hold1073 (.A(\rf_ram.RAM[17][15] ),
    .X(net3307));
 sg13g2_dlygate4sd3_1 hold1074 (.A(\rf_ram.RAM[4][12] ),
    .X(net3308));
 sg13g2_dlygate4sd3_1 hold1075 (.A(\rf_ram.RAM[24][2] ),
    .X(net3309));
 sg13g2_dlygate4sd3_1 hold1076 (.A(\rf_ram.RAM[23][31] ),
    .X(net3310));
 sg13g2_dlygate4sd3_1 hold1077 (.A(\rf_ram.RAM[13][19] ),
    .X(net3311));
 sg13g2_dlygate4sd3_1 hold1078 (.A(\rf_ram.RAM[25][5] ),
    .X(net3312));
 sg13g2_dlygate4sd3_1 hold1079 (.A(\rf_ram.RAM[23][27] ),
    .X(net3313));
 sg13g2_dlygate4sd3_1 hold1080 (.A(\cpu.arbiter.i_wb_cpu_ibus_adr[23] ),
    .X(net3314));
 sg13g2_dlygate4sd3_1 hold1081 (.A(_03907_),
    .X(net3315));
 sg13g2_dlygate4sd3_1 hold1082 (.A(\rf_ram.RAM[20][1] ),
    .X(net3316));
 sg13g2_dlygate4sd3_1 hold1083 (.A(\rf_ram.RAM[27][23] ),
    .X(net3317));
 sg13g2_dlygate4sd3_1 hold1084 (.A(\rf_ram.RAM[5][12] ),
    .X(net3318));
 sg13g2_dlygate4sd3_1 hold1085 (.A(\rf_ram.RAM[31][2] ),
    .X(net3319));
 sg13g2_dlygate4sd3_1 hold1086 (.A(\rf_ram.RAM[27][10] ),
    .X(net3320));
 sg13g2_dlygate4sd3_1 hold1087 (.A(\rf_ram.RAM[19][9] ),
    .X(net3321));
 sg13g2_dlygate4sd3_1 hold1088 (.A(\rf_ram.RAM[1][22] ),
    .X(net3322));
 sg13g2_dlygate4sd3_1 hold1089 (.A(\rf_ram.RAM[24][27] ),
    .X(net3323));
 sg13g2_dlygate4sd3_1 hold1090 (.A(\rf_ram.RAM[28][21] ),
    .X(net3324));
 sg13g2_dlygate4sd3_1 hold1091 (.A(\cpu.arbiter.i_wb_cpu_ibus_adr[17] ),
    .X(net3325));
 sg13g2_dlygate4sd3_1 hold1092 (.A(_03901_),
    .X(net3326));
 sg13g2_dlygate4sd3_1 hold1093 (.A(\cpu.rf_ram_if.rdata0[7] ),
    .X(net3327));
 sg13g2_dlygate4sd3_1 hold1094 (.A(_00027_),
    .X(net3328));
 sg13g2_dlygate4sd3_1 hold1095 (.A(\rf_ram.RAM[26][5] ),
    .X(net3329));
 sg13g2_dlygate4sd3_1 hold1096 (.A(\cpu.rf_ram_if.rdata0[14] ),
    .X(net3330));
 sg13g2_dlygate4sd3_1 hold1097 (.A(_00004_),
    .X(net3331));
 sg13g2_dlygate4sd3_1 hold1098 (.A(\cpu.rf_ram_if.rdata0[25] ),
    .X(net3332));
 sg13g2_dlygate4sd3_1 hold1099 (.A(_00016_),
    .X(net3333));
 sg13g2_dlygate4sd3_1 hold1100 (.A(\cpu.cpu.state.cnt_r[2] ),
    .X(net3334));
 sg13g2_dlygate4sd3_1 hold1101 (.A(\rf_ram.RAM[18][3] ),
    .X(net3335));
 sg13g2_dlygate4sd3_1 hold1102 (.A(\rf_ram.RAM[23][17] ),
    .X(net3336));
 sg13g2_dlygate4sd3_1 hold1103 (.A(\rf_ram.RAM[19][0] ),
    .X(net3337));
 sg13g2_dlygate4sd3_1 hold1104 (.A(\cpu.rf_ram_if.rdata1[18] ),
    .X(net3338));
 sg13g2_dlygate4sd3_1 hold1105 (.A(_00039_),
    .X(net3339));
 sg13g2_dlygate4sd3_1 hold1106 (.A(\cpu.rf_ram_if.rcnt[0] ),
    .X(net3340));
 sg13g2_dlygate4sd3_1 hold1107 (.A(\ram_spi_if.cycle_counter[2] ),
    .X(net3341));
 sg13g2_dlygate4sd3_1 hold1108 (.A(_01410_),
    .X(net3342));
 sg13g2_dlygate4sd3_1 hold1109 (.A(_00067_),
    .X(net3343));
 sg13g2_dlygate4sd3_1 hold1110 (.A(\rf_ram.RAM[22][8] ),
    .X(net3344));
 sg13g2_dlygate4sd3_1 hold1111 (.A(\cpu.rf_ram_if.rdata0[29] ),
    .X(net3345));
 sg13g2_dlygate4sd3_1 hold1112 (.A(_00020_),
    .X(net3346));
 sg13g2_dlygate4sd3_1 hold1113 (.A(\cpu.rf_ram_if.rdata0[18] ),
    .X(net3347));
 sg13g2_dlygate4sd3_1 hold1114 (.A(_00008_),
    .X(net3348));
 sg13g2_dlygate4sd3_1 hold1115 (.A(\cpu.rf_ram_if.rdata0[19] ),
    .X(net3349));
 sg13g2_dlygate4sd3_1 hold1116 (.A(_00009_),
    .X(net3350));
 sg13g2_dlygate4sd3_1 hold1117 (.A(\cpu.rf_ram_if.rdata1[13] ),
    .X(net3351));
 sg13g2_dlygate4sd3_1 hold1118 (.A(_00034_),
    .X(net3352));
 sg13g2_dlygate4sd3_1 hold1119 (.A(\cpu.rf_ram_if.rdata1[16] ),
    .X(net3353));
 sg13g2_dlygate4sd3_1 hold1120 (.A(_00037_),
    .X(net3354));
 sg13g2_dlygate4sd3_1 hold1121 (.A(\cpu.rf_ram_if.rdata1[10] ),
    .X(net3355));
 sg13g2_dlygate4sd3_1 hold1122 (.A(_00060_),
    .X(net3356));
 sg13g2_dlygate4sd3_1 hold1123 (.A(\cpu.rf_ram_if.rdata1[4] ),
    .X(net3357));
 sg13g2_dlygate4sd3_1 hold1124 (.A(_00054_),
    .X(net3358));
 sg13g2_dlygate4sd3_1 hold1125 (.A(\cpu.rf_ram_if.rdata0[5] ),
    .X(net3359));
 sg13g2_dlygate4sd3_1 hold1126 (.A(_00025_),
    .X(net3360));
 sg13g2_dlygate4sd3_1 hold1127 (.A(uo_out[4]),
    .X(net3361));
 sg13g2_dlygate4sd3_1 hold1128 (.A(\cpu.cpu.immdec.gen_immdec_w_eq_1.imm30_25[2] ),
    .X(net3362));
 sg13g2_dlygate4sd3_1 hold1129 (.A(_00523_),
    .X(net3363));
 sg13g2_dlygate4sd3_1 hold1130 (.A(\cpu.cpu.state.cnt_r[1] ),
    .X(net3364));
 sg13g2_dlygate4sd3_1 hold1131 (.A(\cpu.rf_ram_if.rdata1[6] ),
    .X(net3365));
 sg13g2_dlygate4sd3_1 hold1132 (.A(_00056_),
    .X(net3366));
 sg13g2_dlygate4sd3_1 hold1133 (.A(\cpu.arbiter.i_wb_cpu_ibus_adr[26] ),
    .X(net3367));
 sg13g2_dlygate4sd3_1 hold1134 (.A(_03910_),
    .X(net3368));
 sg13g2_dlygate4sd3_1 hold1135 (.A(\cpu.rf_ram_if.rdata1[17] ),
    .X(net3369));
 sg13g2_dlygate4sd3_1 hold1136 (.A(_00038_),
    .X(net3370));
 sg13g2_dlygate4sd3_1 hold1137 (.A(\cpu.rf_ram_if.rdata1[24] ),
    .X(net3371));
 sg13g2_dlygate4sd3_1 hold1138 (.A(_00046_),
    .X(net3372));
 sg13g2_dlygate4sd3_1 hold1139 (.A(\cpu.cpu.immdec.gen_immdec_w_eq_1.imm30_25[3] ),
    .X(net3373));
 sg13g2_dlygate4sd3_1 hold1140 (.A(_00524_),
    .X(net3374));
 sg13g2_dlygate4sd3_1 hold1141 (.A(\cpu.rf_ram_if.rdata0[6] ),
    .X(net3375));
 sg13g2_dlygate4sd3_1 hold1142 (.A(_00026_),
    .X(net3376));
 sg13g2_dlygate4sd3_1 hold1143 (.A(\rf_ram.RAM[7][12] ),
    .X(net3377));
 sg13g2_dlygate4sd3_1 hold1144 (.A(\cpu.rf_ram_if.rdata1[11] ),
    .X(net3378));
 sg13g2_dlygate4sd3_1 hold1145 (.A(_00032_),
    .X(net3379));
 sg13g2_dlygate4sd3_1 hold1146 (.A(\cpu.arbiter.i_wb_cpu_ibus_adr[19] ),
    .X(net3380));
 sg13g2_dlygate4sd3_1 hold1147 (.A(_03903_),
    .X(net3381));
 sg13g2_dlygate4sd3_1 hold1148 (.A(\cpu.arbiter.i_wb_cpu_ibus_adr[29] ),
    .X(net3382));
 sg13g2_dlygate4sd3_1 hold1149 (.A(_03913_),
    .X(net3383));
 sg13g2_dlygate4sd3_1 hold1150 (.A(\cpu.rf_ram_if.rdata0[17] ),
    .X(net3384));
 sg13g2_dlygate4sd3_1 hold1151 (.A(_00007_),
    .X(net3385));
 sg13g2_dlygate4sd3_1 hold1152 (.A(\cpu.arbiter.i_wb_cpu_ibus_adr[30] ),
    .X(net3386));
 sg13g2_dlygate4sd3_1 hold1153 (.A(\rf_ram.RAM[21][8] ),
    .X(net3387));
 sg13g2_dlygate4sd3_1 hold1154 (.A(\rf_ram.RAM[8][10] ),
    .X(net3388));
 sg13g2_dlygate4sd3_1 hold1155 (.A(\cpu.rf_ram_if.rdata0[30] ),
    .X(net3389));
 sg13g2_dlygate4sd3_1 hold1156 (.A(_00021_),
    .X(net3390));
 sg13g2_dlygate4sd3_1 hold1157 (.A(uo_out[5]),
    .X(net3391));
 sg13g2_dlygate4sd3_1 hold1158 (.A(\cpu.arbiter.i_wb_cpu_dbus_adr[2] ),
    .X(net3392));
 sg13g2_dlygate4sd3_1 hold1159 (.A(_00403_),
    .X(net3393));
 sg13g2_dlygate4sd3_1 hold1160 (.A(\cpu.rf_ram_if.rdata0[11] ),
    .X(net3394));
 sg13g2_dlygate4sd3_1 hold1161 (.A(_00001_),
    .X(net3395));
 sg13g2_dlygate4sd3_1 hold1162 (.A(\cpu.rf_ram_if.rdata1[15] ),
    .X(net3396));
 sg13g2_dlygate4sd3_1 hold1163 (.A(_00036_),
    .X(net3397));
 sg13g2_dlygate4sd3_1 hold1164 (.A(\cpu.cpu.immdec.gen_immdec_w_eq_1.imm30_25[1] ),
    .X(net3398));
 sg13g2_dlygate4sd3_1 hold1165 (.A(_00522_),
    .X(net3399));
 sg13g2_dlygate4sd3_1 hold1166 (.A(\cpu.arbiter.i_wb_cpu_ibus_adr[24] ),
    .X(net3400));
 sg13g2_dlygate4sd3_1 hold1167 (.A(\cpu.rf_ram_if.rdata1[22] ),
    .X(net3401));
 sg13g2_dlygate4sd3_1 hold1168 (.A(_00044_),
    .X(net3402));
 sg13g2_dlygate4sd3_1 hold1169 (.A(\cpu.rf_ram_if.rdata0[31] ),
    .X(net3403));
 sg13g2_dlygate4sd3_1 hold1170 (.A(_00023_),
    .X(net3404));
 sg13g2_dlygate4sd3_1 hold1171 (.A(\cpu.rf_ram_if.rdata1[25] ),
    .X(net3405));
 sg13g2_dlygate4sd3_1 hold1172 (.A(_00047_),
    .X(net3406));
 sg13g2_dlygate4sd3_1 hold1173 (.A(\rf_ram.RAM[23][29] ),
    .X(net3407));
 sg13g2_dlygate4sd3_1 hold1174 (.A(\cpu.rf_ram_if.rdata1[5] ),
    .X(net3408));
 sg13g2_dlygate4sd3_1 hold1175 (.A(_00055_),
    .X(net3409));
 sg13g2_dlygate4sd3_1 hold1176 (.A(\cpu.rf_ram_if.rdata0[26] ),
    .X(net3410));
 sg13g2_dlygate4sd3_1 hold1177 (.A(_00017_),
    .X(net3411));
 sg13g2_dlygate4sd3_1 hold1178 (.A(\cpu.rf_ram_if.rdata1[29] ),
    .X(net3412));
 sg13g2_dlygate4sd3_1 hold1179 (.A(_00051_),
    .X(net3413));
 sg13g2_dlygate4sd3_1 hold1180 (.A(\cpu.rf_ram_if.rdata1[30] ),
    .X(net3414));
 sg13g2_dlygate4sd3_1 hold1181 (.A(_00052_),
    .X(net3415));
 sg13g2_dlygate4sd3_1 hold1182 (.A(\cpu.rf_ram_if.rdata0[13] ),
    .X(net3416));
 sg13g2_dlygate4sd3_1 hold1183 (.A(_00003_),
    .X(net3417));
 sg13g2_dlygate4sd3_1 hold1184 (.A(\cpu.cpu.csr_imm [0]),
    .X(net3418));
 sg13g2_dlygate4sd3_1 hold1185 (.A(_00532_),
    .X(net3419));
 sg13g2_dlygate4sd3_1 hold1186 (.A(\cpu.cpu.immdec.gen_immdec_w_eq_1.imm30_25[5] ),
    .X(net3420));
 sg13g2_dlygate4sd3_1 hold1187 (.A(_00526_),
    .X(net3421));
 sg13g2_dlygate4sd3_1 hold1188 (.A(\cpu.rf_ram_if.rdata0[10] ),
    .X(net3422));
 sg13g2_dlygate4sd3_1 hold1189 (.A(_00030_),
    .X(net3423));
 sg13g2_dlygate4sd3_1 hold1190 (.A(\cpu.rf_ram_if.rdata1[28] ),
    .X(net3424));
 sg13g2_dlygate4sd3_1 hold1191 (.A(_00050_),
    .X(net3425));
 sg13g2_dlygate4sd3_1 hold1192 (.A(\cpu.arbiter.i_wb_cpu_ibus_adr[31] ),
    .X(net3426));
 sg13g2_dlygate4sd3_1 hold1193 (.A(\cpu.rf_ram_if.rdata0[23] ),
    .X(net3427));
 sg13g2_dlygate4sd3_1 hold1194 (.A(_00014_),
    .X(net3428));
 sg13g2_dlygate4sd3_1 hold1195 (.A(\cpu.arbiter.i_wb_cpu_ibus_adr[18] ),
    .X(net3429));
 sg13g2_dlygate4sd3_1 hold1196 (.A(\cpu.rf_ram_if.rdata1[12] ),
    .X(net3430));
 sg13g2_dlygate4sd3_1 hold1197 (.A(_00033_),
    .X(net3431));
 sg13g2_dlygate4sd3_1 hold1198 (.A(\cpu.cpu.ctrl.pc_plus_4_cy_r_w [0]),
    .X(net3432));
 sg13g2_dlygate4sd3_1 hold1199 (.A(_01500_),
    .X(net3433));
 sg13g2_dlygate4sd3_1 hold1200 (.A(_00063_),
    .X(net3434));
 sg13g2_dlygate4sd3_1 hold1201 (.A(\cpu.cpu.immdec.gen_immdec_w_eq_1.imm19_12_20[3] ),
    .X(net3435));
 sg13g2_dlygate4sd3_1 hold1202 (.A(_00531_),
    .X(net3436));
 sg13g2_dlygate4sd3_1 hold1203 (.A(\cpu.arbiter.i_wb_cpu_ibus_adr[28] ),
    .X(net3437));
 sg13g2_dlygate4sd3_1 hold1204 (.A(_03912_),
    .X(net3438));
 sg13g2_dlygate4sd3_1 hold1205 (.A(\cpu.cpu.state.cnt_r[0] ),
    .X(net3439));
 sg13g2_dlygate4sd3_1 hold1206 (.A(\cpu.cpu.immdec.gen_immdec_w_eq_1.imm19_12_20[1] ),
    .X(net3440));
 sg13g2_dlygate4sd3_1 hold1207 (.A(_00529_),
    .X(net3441));
 sg13g2_dlygate4sd3_1 hold1208 (.A(\cpu.rf_ram_if.rdata0[28] ),
    .X(net3442));
 sg13g2_dlygate4sd3_1 hold1209 (.A(_00019_),
    .X(net3443));
 sg13g2_dlygate4sd3_1 hold1210 (.A(\cpu.rf_ram_if.rdata1[7] ),
    .X(net3444));
 sg13g2_dlygate4sd3_1 hold1211 (.A(_00057_),
    .X(net3445));
 sg13g2_dlygate4sd3_1 hold1212 (.A(\cpu.rf_ram_if.rdata1[26] ),
    .X(net3446));
 sg13g2_dlygate4sd3_1 hold1213 (.A(_00048_),
    .X(net3447));
 sg13g2_dlygate4sd3_1 hold1214 (.A(\cpu.rf_ram_if.rdata0[12] ),
    .X(net3448));
 sg13g2_dlygate4sd3_1 hold1215 (.A(_00002_),
    .X(net3449));
 sg13g2_dlygate4sd3_1 hold1216 (.A(\cpu.arbiter.i_wb_cpu_dbus_dat[30] ),
    .X(net3450));
 sg13g2_dlygate4sd3_1 hold1217 (.A(_00546_),
    .X(net3451));
 sg13g2_dlygate4sd3_1 hold1218 (.A(\cpu.rf_ram_if.rdata0[9] ),
    .X(net3452));
 sg13g2_dlygate4sd3_1 hold1219 (.A(_00029_),
    .X(net3453));
 sg13g2_dlygate4sd3_1 hold1220 (.A(\cpu.arbiter.i_wb_cpu_ibus_adr[27] ),
    .X(net3454));
 sg13g2_dlygate4sd3_1 hold1221 (.A(\cpu.arbiter.i_wb_cpu_ibus_adr[16] ),
    .X(net3455));
 sg13g2_dlygate4sd3_1 hold1222 (.A(_03900_),
    .X(net3456));
 sg13g2_dlygate4sd3_1 hold1223 (.A(\cpu.cpu.immdec.gen_immdec_w_eq_1.imm30_25[4] ),
    .X(net3457));
 sg13g2_dlygate4sd3_1 hold1224 (.A(_00525_),
    .X(net3458));
 sg13g2_dlygate4sd3_1 hold1225 (.A(\cpu.rf_ram_if.rdata0[27] ),
    .X(net3459));
 sg13g2_dlygate4sd3_1 hold1226 (.A(_00018_),
    .X(net3460));
 sg13g2_dlygate4sd3_1 hold1227 (.A(\ram_spi_if.cycle_counter[4] ),
    .X(net3461));
 sg13g2_dlygate4sd3_1 hold1228 (.A(_01414_),
    .X(net3462));
 sg13g2_dlygate4sd3_1 hold1229 (.A(_00069_),
    .X(net3463));
 sg13g2_dlygate4sd3_1 hold1230 (.A(\cpu.arbiter.i_wb_cpu_dbus_dat[31] ),
    .X(net3464));
 sg13g2_dlygate4sd3_1 hold1231 (.A(_00547_),
    .X(net3465));
 sg13g2_dlygate4sd3_1 hold1232 (.A(\cpu.rf_ram_if.rdata0[16] ),
    .X(net3466));
 sg13g2_dlygate4sd3_1 hold1233 (.A(_00006_),
    .X(net3467));
 sg13g2_dlygate4sd3_1 hold1234 (.A(\cpu.rf_ram_if.rdata1[27] ),
    .X(net3468));
 sg13g2_dlygate4sd3_1 hold1235 (.A(_00049_),
    .X(net3469));
 sg13g2_dlygate4sd3_1 hold1236 (.A(\cpu.rf_ram_if.rdata1[9] ),
    .X(net3470));
 sg13g2_dlygate4sd3_1 hold1237 (.A(_00059_),
    .X(net3471));
 sg13g2_dlygate4sd3_1 hold1238 (.A(\cpu.arbiter.i_wb_cpu_ibus_adr[1] ),
    .X(net3472));
 sg13g2_dlygate4sd3_1 hold1239 (.A(_03885_),
    .X(net3473));
 sg13g2_dlygate4sd3_1 hold1240 (.A(\cpu.arbiter.i_wb_cpu_ibus_adr[21] ),
    .X(net3474));
 sg13g2_dlygate4sd3_1 hold1241 (.A(_03905_),
    .X(net3475));
 sg13g2_dlygate4sd3_1 hold1242 (.A(\ram_spi_if.spi_mosi ),
    .X(net3476));
 sg13g2_dlygate4sd3_1 hold1243 (.A(\cpu.cpu.immdec.gen_immdec_w_eq_1.imm11_7[0] ),
    .X(net3477));
 sg13g2_dlygate4sd3_1 hold1244 (.A(_00614_),
    .X(net3478));
 sg13g2_dlygate4sd3_1 hold1245 (.A(\cpu.arbiter.i_wb_cpu_ibus_adr[14] ),
    .X(net3479));
 sg13g2_dlygate4sd3_1 hold1246 (.A(_03898_),
    .X(net3480));
 sg13g2_dlygate4sd3_1 hold1247 (.A(\cpu.arbiter.i_wb_cpu_ibus_adr[22] ),
    .X(net3481));
 sg13g2_dlygate4sd3_1 hold1248 (.A(\cpu.rf_ram_if.rdata1[8] ),
    .X(net3482));
 sg13g2_dlygate4sd3_1 hold1249 (.A(_00058_),
    .X(net3483));
 sg13g2_dlygate4sd3_1 hold1250 (.A(\cpu.arbiter.i_wb_cpu_ibus_adr[25] ),
    .X(net3484));
 sg13g2_dlygate4sd3_1 hold1251 (.A(\cpu.arbiter.i_wb_mem_rdt[17] ),
    .X(net3485));
 sg13g2_dlygate4sd3_1 hold1252 (.A(_00317_),
    .X(net3486));
 sg13g2_dlygate4sd3_1 hold1253 (.A(\cpu.cpu.immdec.gen_immdec_w_eq_1.imm19_12_20[2] ),
    .X(net3487));
 sg13g2_dlygate4sd3_1 hold1254 (.A(_00530_),
    .X(net3488));
 sg13g2_dlygate4sd3_1 hold1255 (.A(\cpu.cpu.ctrl.i_jump ),
    .X(net3489));
 sg13g2_dlygate4sd3_1 hold1256 (.A(\cpu.arbiter.i_wb_cpu_ibus_adr[13] ),
    .X(net3490));
 sg13g2_dlygate4sd3_1 hold1257 (.A(_03897_),
    .X(net3491));
 sg13g2_dlygate4sd3_1 hold1258 (.A(\cpu.cpu.state.cnt_r[3] ),
    .X(net3492));
 sg13g2_dlygate4sd3_1 hold1259 (.A(_00474_),
    .X(net3493));
 sg13g2_dlygate4sd3_1 hold1260 (.A(\cpu.arbiter.i_wb_mem_rdt[16] ),
    .X(net3494));
 sg13g2_dlygate4sd3_1 hold1261 (.A(_00316_),
    .X(net3495));
 sg13g2_dlygate4sd3_1 hold1262 (.A(\ram_spi_if.cycle_counter[3] ),
    .X(net3496));
 sg13g2_dlygate4sd3_1 hold1263 (.A(_00068_),
    .X(net3497));
 sg13g2_dlygate4sd3_1 hold1264 (.A(\cpu.rf_ram_if.rdata0[4] ),
    .X(net3498));
 sg13g2_dlygate4sd3_1 hold1265 (.A(_00024_),
    .X(net3499));
 sg13g2_dlygate4sd3_1 hold1266 (.A(\cpu.arbiter.i_wb_cpu_ibus_adr[7] ),
    .X(net3500));
 sg13g2_dlygate4sd3_1 hold1267 (.A(_03891_),
    .X(net3501));
 sg13g2_dlygate4sd3_1 hold1268 (.A(\cpu.i_rf_rdata[20] ),
    .X(net3502));
 sg13g2_dlygate4sd3_1 hold1269 (.A(_00041_),
    .X(net3503));
 sg13g2_dlygate4sd3_1 hold1270 (.A(\cpu.rf_ram_if.rdata0[8] ),
    .X(net3504));
 sg13g2_dlygate4sd3_1 hold1271 (.A(_00028_),
    .X(net3505));
 sg13g2_dlygate4sd3_1 hold1272 (.A(\cpu.arbiter.i_wb_cpu_dbus_adr[24] ),
    .X(net3506));
 sg13g2_dlygate4sd3_1 hold1273 (.A(_00424_),
    .X(net3507));
 sg13g2_dlygate4sd3_1 hold1274 (.A(\cpu.arbiter.i_wb_cpu_dbus_adr[29] ),
    .X(net3508));
 sg13g2_dlygate4sd3_1 hold1275 (.A(_00429_),
    .X(net3509));
 sg13g2_dlygate4sd3_1 hold1276 (.A(\cpu.cpu.immdec.gen_immdec_w_eq_1.imm19_12_20[0] ),
    .X(net3510));
 sg13g2_dlygate4sd3_1 hold1277 (.A(_00528_),
    .X(net3511));
 sg13g2_dlygate4sd3_1 hold1278 (.A(\cpu.rf_ram_if.rdata1[19] ),
    .X(net3512));
 sg13g2_dlygate4sd3_1 hold1279 (.A(_00040_),
    .X(net3513));
 sg13g2_dlygate4sd3_1 hold1280 (.A(\cpu.arbiter.i_wb_cpu_dbus_adr[17] ),
    .X(net3514));
 sg13g2_dlygate4sd3_1 hold1281 (.A(_00417_),
    .X(net3515));
 sg13g2_dlygate4sd3_1 hold1282 (.A(\cpu.cpu.decode.co_ebreak ),
    .X(net3516));
 sg13g2_dlygate4sd3_1 hold1283 (.A(_00515_),
    .X(net3517));
 sg13g2_dlygate4sd3_1 hold1284 (.A(\cpu.arbiter.i_wb_cpu_ibus_adr[20] ),
    .X(net3518));
 sg13g2_dlygate4sd3_1 hold1285 (.A(\cpu.arbiter.i_wb_cpu_dbus_dat[21] ),
    .X(net3519));
 sg13g2_dlygate4sd3_1 hold1286 (.A(_00504_),
    .X(net3520));
 sg13g2_dlygate4sd3_1 hold1287 (.A(\cpu.arbiter.i_wb_cpu_dbus_dat[20] ),
    .X(net3521));
 sg13g2_dlygate4sd3_1 hold1288 (.A(_00503_),
    .X(net3522));
 sg13g2_dlygate4sd3_1 hold1289 (.A(\cpu.rf_ram_if.rdata1[14] ),
    .X(net3523));
 sg13g2_dlygate4sd3_1 hold1290 (.A(_00035_),
    .X(net3524));
 sg13g2_dlygate4sd3_1 hold1291 (.A(\cpu.rf_ram_if.rdata0[20] ),
    .X(net3525));
 sg13g2_dlygate4sd3_1 hold1292 (.A(_00010_),
    .X(net3526));
 sg13g2_dlygate4sd3_1 hold1293 (.A(\cpu.arbiter.i_wb_cpu_ibus_adr[8] ),
    .X(net3527));
 sg13g2_dlygate4sd3_1 hold1294 (.A(\cpu.arbiter.i_wb_cpu_dbus_adr[16] ),
    .X(net3528));
 sg13g2_dlygate4sd3_1 hold1295 (.A(_00416_),
    .X(net3529));
 sg13g2_dlygate4sd3_1 hold1296 (.A(\cpu.rf_ram_if.rdata0[15] ),
    .X(net3530));
 sg13g2_dlygate4sd3_1 hold1297 (.A(_00005_),
    .X(net3531));
 sg13g2_dlygate4sd3_1 hold1298 (.A(\cpu.rf_ram_if.rgnt ),
    .X(net3532));
 sg13g2_dlygate4sd3_1 hold1299 (.A(_03670_),
    .X(net3533));
 sg13g2_dlygate4sd3_1 hold1300 (.A(\cpu.arbiter.i_wb_cpu_ibus_adr[3] ),
    .X(net3534));
 sg13g2_dlygate4sd3_1 hold1301 (.A(_03887_),
    .X(net3535));
 sg13g2_dlygate4sd3_1 hold1302 (.A(\cpu.arbiter.i_wb_mem_rdt[26] ),
    .X(net3536));
 sg13g2_dlygate4sd3_1 hold1303 (.A(_00326_),
    .X(net3537));
 sg13g2_dlygate4sd3_1 hold1304 (.A(\cpu.rf_ram_if.rdata1[3] ),
    .X(net3538));
 sg13g2_dlygate4sd3_1 hold1305 (.A(_00053_),
    .X(net3539));
 sg13g2_dlygate4sd3_1 hold1306 (.A(\cpu.arbiter.i_wb_cpu_dbus_adr[30] ),
    .X(net3540));
 sg13g2_dlygate4sd3_1 hold1307 (.A(\cpu.arbiter.i_wb_cpu_dbus_adr[18] ),
    .X(net3541));
 sg13g2_dlygate4sd3_1 hold1308 (.A(\cpu.arbiter.i_wb_cpu_ibus_adr[12] ),
    .X(net3542));
 sg13g2_dlygate4sd3_1 hold1309 (.A(_03896_),
    .X(net3543));
 sg13g2_dlygate4sd3_1 hold1310 (.A(\cpu.arbiter.i_wb_cpu_ibus_adr[2] ),
    .X(net3544));
 sg13g2_dlygate4sd3_1 hold1311 (.A(\cpu.arbiter.i_wb_cpu_dbus_adr[25] ),
    .X(net3545));
 sg13g2_dlygate4sd3_1 hold1312 (.A(\cpu.arbiter.i_wb_cpu_dbus_dat[10] ),
    .X(net3546));
 sg13g2_dlygate4sd3_1 hold1313 (.A(_00493_),
    .X(net3547));
 sg13g2_dlygate4sd3_1 hold1314 (.A(\cpu.arbiter.i_wb_cpu_dbus_dat[12] ),
    .X(net3548));
 sg13g2_dlygate4sd3_1 hold1315 (.A(_00495_),
    .X(net3549));
 sg13g2_dlygate4sd3_1 hold1316 (.A(\cpu.arbiter.i_wb_cpu_dbus_dat[22] ),
    .X(net3550));
 sg13g2_dlygate4sd3_1 hold1317 (.A(_00505_),
    .X(net3551));
 sg13g2_dlygate4sd3_1 hold1318 (.A(\cpu.arbiter.i_wb_cpu_dbus_dat[9] ),
    .X(net3552));
 sg13g2_dlygate4sd3_1 hold1319 (.A(_00492_),
    .X(net3553));
 sg13g2_dlygate4sd3_1 hold1320 (.A(\cpu.arbiter.i_wb_cpu_dbus_adr[27] ),
    .X(net3554));
 sg13g2_dlygate4sd3_1 hold1321 (.A(_00428_),
    .X(net3555));
 sg13g2_dlygate4sd3_1 hold1322 (.A(\cpu.arbiter.i_wb_mem_rdt[25] ),
    .X(net3556));
 sg13g2_dlygate4sd3_1 hold1323 (.A(_00325_),
    .X(net3557));
 sg13g2_dlygate4sd3_1 hold1324 (.A(\cpu.arbiter.i_wb_mem_rdt[20] ),
    .X(net3558));
 sg13g2_dlygate4sd3_1 hold1325 (.A(_00320_),
    .X(net3559));
 sg13g2_dlygate4sd3_1 hold1326 (.A(\cpu.arbiter.i_wb_cpu_dbus_adr[26] ),
    .X(net3560));
 sg13g2_dlygate4sd3_1 hold1327 (.A(\cpu.arbiter.i_wb_cpu_dbus_adr[22] ),
    .X(net3561));
 sg13g2_dlygate4sd3_1 hold1328 (.A(_00423_),
    .X(net3562));
 sg13g2_dlygate4sd3_1 hold1329 (.A(\cpu.arbiter.i_wb_cpu_dbus_adr[21] ),
    .X(net3563));
 sg13g2_dlygate4sd3_1 hold1330 (.A(\cpu.arbiter.i_wb_cpu_dbus_adr[19] ),
    .X(net3564));
 sg13g2_dlygate4sd3_1 hold1331 (.A(\cpu.arbiter.i_wb_mem_rdt[18] ),
    .X(net3565));
 sg13g2_dlygate4sd3_1 hold1332 (.A(_00318_),
    .X(net3566));
 sg13g2_dlygate4sd3_1 hold1333 (.A(\cpu.arbiter.i_wb_cpu_ibus_adr[11] ),
    .X(net3567));
 sg13g2_dlygate4sd3_1 hold1334 (.A(_03895_),
    .X(net3568));
 sg13g2_dlygate4sd3_1 hold1335 (.A(\cpu.arbiter.i_wb_cpu_ibus_adr[10] ),
    .X(net3569));
 sg13g2_dlygate4sd3_1 hold1336 (.A(_03894_),
    .X(net3570));
 sg13g2_dlygate4sd3_1 hold1337 (.A(\cpu.cpu.alu.cmp_r ),
    .X(net3571));
 sg13g2_dlygate4sd3_1 hold1338 (.A(\cpu.rf_ram_if.rdata0[24] ),
    .X(net3572));
 sg13g2_dlygate4sd3_1 hold1339 (.A(_00015_),
    .X(net3573));
 sg13g2_dlygate4sd3_1 hold1340 (.A(\cpu.i_rf_rdata[2] ),
    .X(net3574));
 sg13g2_dlygate4sd3_1 hold1341 (.A(_00022_),
    .X(net3575));
 sg13g2_dlygate4sd3_1 hold1342 (.A(\cpu.arbiter.i_wb_cpu_dbus_dat[2] ),
    .X(net3576));
 sg13g2_dlygate4sd3_1 hold1343 (.A(_00485_),
    .X(net3577));
 sg13g2_dlygate4sd3_1 hold1344 (.A(\cpu.cpu.immdec.gen_immdec_w_eq_1.imm19_12_20[7] ),
    .X(net3578));
 sg13g2_dlygate4sd3_1 hold1345 (.A(_00535_),
    .X(net3579));
 sg13g2_dlygate4sd3_1 hold1346 (.A(\cpu.arbiter.i_wb_cpu_dbus_dat[19] ),
    .X(net3580));
 sg13g2_dlygate4sd3_1 hold1347 (.A(_00502_),
    .X(net3581));
 sg13g2_dlygate4sd3_1 hold1348 (.A(\cpu.cpu.immdec.gen_immdec_w_eq_1.imm11_7[1] ),
    .X(net3582));
 sg13g2_dlygate4sd3_1 hold1349 (.A(_00615_),
    .X(net3583));
 sg13g2_dlygate4sd3_1 hold1350 (.A(\cpu.arbiter.i_wb_mem_rdt[24] ),
    .X(net3584));
 sg13g2_dlygate4sd3_1 hold1351 (.A(_00324_),
    .X(net3585));
 sg13g2_dlygate4sd3_1 hold1352 (.A(\cpu.arbiter.i_wb_cpu_dbus_dat[16] ),
    .X(net3586));
 sg13g2_dlygate4sd3_1 hold1353 (.A(_02693_),
    .X(net3587));
 sg13g2_dlygate4sd3_1 hold1354 (.A(\cpu.arbiter.i_wb_cpu_dbus_dat[17] ),
    .X(net3588));
 sg13g2_dlygate4sd3_1 hold1355 (.A(_00500_),
    .X(net3589));
 sg13g2_dlygate4sd3_1 hold1356 (.A(\cpu.arbiter.i_wb_cpu_dbus_we ),
    .X(net3590));
 sg13g2_dlygate4sd3_1 hold1357 (.A(\cpu.arbiter.i_wb_mem_rdt[29] ),
    .X(net3591));
 sg13g2_dlygate4sd3_1 hold1358 (.A(_02731_),
    .X(net3592));
 sg13g2_dlygate4sd3_1 hold1359 (.A(_00329_),
    .X(net3593));
 sg13g2_dlygate4sd3_1 hold1360 (.A(\cpu.arbiter.i_wb_mem_rdt[0] ),
    .X(net3594));
 sg13g2_dlygate4sd3_1 hold1361 (.A(_01012_),
    .X(net3595));
 sg13g2_dlygate4sd3_1 hold1362 (.A(\cpu.arbiter.i_wb_cpu_ibus_adr[6] ),
    .X(net3596));
 sg13g2_dlygate4sd3_1 hold1363 (.A(_03890_),
    .X(net3597));
 sg13g2_dlygate4sd3_1 hold1364 (.A(\cpu.arbiter.i_wb_cpu_dbus_dat[15] ),
    .X(net3598));
 sg13g2_dlygate4sd3_1 hold1365 (.A(_00498_),
    .X(net3599));
 sg13g2_dlygate4sd3_1 hold1366 (.A(\cpu.cpu.bufreg.c_r [0]),
    .X(net3600));
 sg13g2_dlygate4sd3_1 hold1367 (.A(_01476_),
    .X(net3601));
 sg13g2_dlygate4sd3_1 hold1368 (.A(\cpu.arbiter.i_wb_mem_rdt[27] ),
    .X(net3602));
 sg13g2_dlygate4sd3_1 hold1369 (.A(_00327_),
    .X(net3603));
 sg13g2_dlygate4sd3_1 hold1370 (.A(\cpu.rf_ram_if.rdata1[23] ),
    .X(net3604));
 sg13g2_dlygate4sd3_1 hold1371 (.A(_00045_),
    .X(net3605));
 sg13g2_dlygate4sd3_1 hold1372 (.A(\cpu.rf_ram_if.wen0_r ),
    .X(net3606));
 sg13g2_dlygate4sd3_1 hold1373 (.A(_00472_),
    .X(net3607));
 sg13g2_dlygate4sd3_1 hold1374 (.A(\cpu.arbiter.i_wb_cpu_ibus_adr[15] ),
    .X(net3608));
 sg13g2_dlygate4sd3_1 hold1375 (.A(\cpu.cpu.state.ibus_cyc ),
    .X(net3609));
 sg13g2_dlygate4sd3_1 hold1376 (.A(\cpu.arbiter.i_wb_cpu_dbus_dat[11] ),
    .X(net3610));
 sg13g2_dlygate4sd3_1 hold1377 (.A(_00494_),
    .X(net3611));
 sg13g2_dlygate4sd3_1 hold1378 (.A(\cpu.arbiter.i_wb_cpu_dbus_dat[0] ),
    .X(net3612));
 sg13g2_dlygate4sd3_1 hold1379 (.A(\cpu.arbiter.i_wb_mem_rdt[28] ),
    .X(net3613));
 sg13g2_dlygate4sd3_1 hold1380 (.A(_00328_),
    .X(net3614));
 sg13g2_dlygate4sd3_1 hold1381 (.A(\cpu.cpu.immdec.gen_immdec_w_eq_1.imm19_12_20[6] ),
    .X(net3615));
 sg13g2_dlygate4sd3_1 hold1382 (.A(\cpu.cpu.immdec.gen_immdec_w_eq_1.imm19_12_20[5] ),
    .X(net3616));
 sg13g2_dlygate4sd3_1 hold1383 (.A(\cpu.arbiter.i_wb_cpu_dbus_dat[13] ),
    .X(net3617));
 sg13g2_dlygate4sd3_1 hold1384 (.A(_00496_),
    .X(net3618));
 sg13g2_dlygate4sd3_1 hold1385 (.A(\cpu.rf_ram_if.rcnt[3] ),
    .X(net3619));
 sg13g2_dlygate4sd3_1 hold1386 (.A(_02688_),
    .X(net3620));
 sg13g2_dlygate4sd3_1 hold1387 (.A(\cpu.arbiter.i_wb_cpu_dbus_dat[3] ),
    .X(net3621));
 sg13g2_dlygate4sd3_1 hold1388 (.A(\cpu.arbiter.i_wb_cpu_dbus_adr[20] ),
    .X(net3622));
 sg13g2_dlygate4sd3_1 hold1389 (.A(\cpu.cpu.immdec.gen_immdec_w_eq_1.imm19_12_20[8] ),
    .X(net3623));
 sg13g2_dlygate4sd3_1 hold1390 (.A(_03815_),
    .X(net3624));
 sg13g2_dlygate4sd3_1 hold1391 (.A(_00536_),
    .X(net3625));
 sg13g2_dlygate4sd3_1 hold1392 (.A(\cpu.arbiter.i_wb_mem_rdt[10] ),
    .X(net3626));
 sg13g2_dlygate4sd3_1 hold1393 (.A(_01022_),
    .X(net3627));
 sg13g2_dlygate4sd3_1 hold1394 (.A(\cpu.arbiter.i_wb_mem_rdt[14] ),
    .X(net3628));
 sg13g2_dlygate4sd3_1 hold1395 (.A(_01026_),
    .X(net3629));
 sg13g2_dlygate4sd3_1 hold1396 (.A(\cpu.arbiter.i_wb_cpu_ibus_adr[4] ),
    .X(net3630));
 sg13g2_dlygate4sd3_1 hold1397 (.A(\cpu.arbiter.i_wb_cpu_dbus_dat[18] ),
    .X(net3631));
 sg13g2_dlygate4sd3_1 hold1398 (.A(\cpu.arbiter.i_wb_cpu_dbus_dat[6] ),
    .X(net3632));
 sg13g2_dlygate4sd3_1 hold1399 (.A(_00489_),
    .X(net3633));
 sg13g2_dlygate4sd3_1 hold1400 (.A(\cpu.arbiter.i_wb_cpu_ibus_adr[5] ),
    .X(net3634));
 sg13g2_dlygate4sd3_1 hold1401 (.A(\cpu.arbiter.i_wb_cpu_dbus_dat[4] ),
    .X(net3635));
 sg13g2_dlygate4sd3_1 hold1402 (.A(_00487_),
    .X(net3636));
 sg13g2_dlygate4sd3_1 hold1403 (.A(\cpu.arbiter.i_wb_mem_rdt[2] ),
    .X(net3637));
 sg13g2_dlygate4sd3_1 hold1404 (.A(_01014_),
    .X(net3638));
 sg13g2_dlygate4sd3_1 hold1405 (.A(\cpu.arbiter.i_wb_cpu_dbus_dat[14] ),
    .X(net3639));
 sg13g2_dlygate4sd3_1 hold1406 (.A(\cpu.cpu.immdec.gen_immdec_w_eq_1.imm31 ),
    .X(net3640));
 sg13g2_dlygate4sd3_1 hold1407 (.A(_00537_),
    .X(net3641));
 sg13g2_dlygate4sd3_1 hold1408 (.A(\cpu.i_wb_ext_rdt[3] ),
    .X(net3642));
 sg13g2_dlygate4sd3_1 hold1409 (.A(_03695_),
    .X(net3643));
 sg13g2_dlygate4sd3_1 hold1410 (.A(\cpu.i_rf_rdata[0] ),
    .X(net3644));
 sg13g2_dlygate4sd3_1 hold1411 (.A(_00000_),
    .X(net3645));
 sg13g2_dlygate4sd3_1 hold1412 (.A(\cpu.rf_ram_if.rdata1[1] ),
    .X(net3646));
 sg13g2_dlygate4sd3_1 hold1413 (.A(_00031_),
    .X(net3647));
 sg13g2_dlygate4sd3_1 hold1414 (.A(\cpu.arbiter.i_wb_cpu_dbus_dat[7] ),
    .X(net3648));
 sg13g2_dlygate4sd3_1 hold1415 (.A(_00490_),
    .X(net3649));
 sg13g2_dlygate4sd3_1 hold1416 (.A(\cpu.arbiter.i_wb_cpu_dbus_dat[23] ),
    .X(net3650));
 sg13g2_dlygate4sd3_1 hold1417 (.A(_00506_),
    .X(net3651));
 sg13g2_dlygate4sd3_1 hold1418 (.A(\cpu.arbiter.i_wb_cpu_dbus_dat[1] ),
    .X(net3652));
 sg13g2_dlygate4sd3_1 hold1419 (.A(\cpu.arbiter.i_wb_mem_rdt[19] ),
    .X(net3653));
 sg13g2_dlygate4sd3_1 hold1420 (.A(\cpu.arbiter.i_wb_cpu_dbus_adr[6] ),
    .X(net3654));
 sg13g2_dlygate4sd3_1 hold1421 (.A(_00407_),
    .X(net3655));
 sg13g2_dlygate4sd3_1 hold1422 (.A(\cpu.rf_ram_if.rdata0[2] ),
    .X(net3656));
 sg13g2_dlygate4sd3_1 hold1423 (.A(_00011_),
    .X(net3657));
 sg13g2_dlygate4sd3_1 hold1424 (.A(\cpu.i_wb_ext_rdt[1] ),
    .X(net3658));
 sg13g2_dlygate4sd3_1 hold1425 (.A(_03685_),
    .X(net3659));
 sg13g2_dlygate4sd3_1 hold1426 (.A(\cpu.cpu.bne_or_bge ),
    .X(net3660));
 sg13g2_dlygate4sd3_1 hold1427 (.A(_03667_),
    .X(net3661));
 sg13g2_dlygate4sd3_1 hold1428 (.A(\cpu.arbiter.i_wb_cpu_dbus_adr[11] ),
    .X(net3662));
 sg13g2_dlygate4sd3_1 hold1429 (.A(_00411_),
    .X(net3663));
 sg13g2_dlygate4sd3_1 hold1430 (.A(\cpu.arbiter.i_wb_cpu_dbus_adr[8] ),
    .X(net3664));
 sg13g2_dlygate4sd3_1 hold1431 (.A(_00408_),
    .X(net3665));
 sg13g2_dlygate4sd3_1 hold1432 (.A(\cpu.arbiter.i_wb_cpu_ibus_adr[9] ),
    .X(net3666));
 sg13g2_dlygate4sd3_1 hold1433 (.A(\cpu.arbiter.i_wb_cpu_dbus_adr[9] ),
    .X(net3667));
 sg13g2_dlygate4sd3_1 hold1434 (.A(\cpu.arbiter.i_wb_mem_rdt[1] ),
    .X(net3668));
 sg13g2_dlygate4sd3_1 hold1435 (.A(\cpu.arbiter.i_wb_mem_rdt[12] ),
    .X(net3669));
 sg13g2_dlygate4sd3_1 hold1436 (.A(\cpu.arbiter.i_wb_cpu_dbus_adr[5] ),
    .X(net3670));
 sg13g2_dlygate4sd3_1 hold1437 (.A(\cpu.arbiter.i_wb_cpu_dbus_adr[14] ),
    .X(net3671));
 sg13g2_dlygate4sd3_1 hold1438 (.A(_00414_),
    .X(net3672));
 sg13g2_dlygate4sd3_1 hold1439 (.A(\cpu.rf_ram_if.rdata1[2] ),
    .X(net3673));
 sg13g2_dlygate4sd3_1 hold1440 (.A(\cpu.arbiter.i_wb_cpu_dbus_dat[27] ),
    .X(net3674));
 sg13g2_dlygate4sd3_1 hold1441 (.A(_00543_),
    .X(net3675));
 sg13g2_dlygate4sd3_1 hold1442 (.A(\cpu.arbiter.i_wb_cpu_dbus_adr[3] ),
    .X(net3676));
 sg13g2_dlygate4sd3_1 hold1443 (.A(_00404_),
    .X(net3677));
 sg13g2_dlygate4sd3_1 hold1444 (.A(\cpu.arbiter.i_wb_mem_rdt[5] ),
    .X(net3678));
 sg13g2_dlygate4sd3_1 hold1445 (.A(_01017_),
    .X(net3679));
 sg13g2_dlygate4sd3_1 hold1446 (.A(\cpu.arbiter.i_wb_mem_rdt[22] ),
    .X(net3680));
 sg13g2_dlygate4sd3_1 hold1447 (.A(_02711_),
    .X(net3681));
 sg13g2_dlygate4sd3_1 hold1448 (.A(_00322_),
    .X(net3682));
 sg13g2_dlygate4sd3_1 hold1449 (.A(\cpu.arbiter.i_wb_mem_rdt[6] ),
    .X(net3683));
 sg13g2_dlygate4sd3_1 hold1450 (.A(\cpu.arbiter.i_wb_cpu_dbus_adr[15] ),
    .X(net3684));
 sg13g2_dlygate4sd3_1 hold1451 (.A(\cpu.arbiter.i_wb_cpu_dbus_adr[12] ),
    .X(net3685));
 sg13g2_dlygate4sd3_1 hold1452 (.A(\cpu.arbiter.i_wb_cpu_dbus_dat[5] ),
    .X(net3686));
 sg13g2_dlygate4sd3_1 hold1453 (.A(_00488_),
    .X(net3687));
 sg13g2_dlygate4sd3_1 hold1454 (.A(\cpu.arbiter.i_wb_mem_rdt[31] ),
    .X(net3688));
 sg13g2_dlygate4sd3_1 hold1455 (.A(_00330_),
    .X(net3689));
 sg13g2_dlygate4sd3_1 hold1456 (.A(\cpu.arbiter.i_wb_mem_rdt[3] ),
    .X(net3690));
 sg13g2_dlygate4sd3_1 hold1457 (.A(\ram_spi_if.cycle_counter[1] ),
    .X(net3691));
 sg13g2_dlygate4sd3_1 hold1458 (.A(\cpu.arbiter.i_wb_mem_rdt[8] ),
    .X(net3692));
 sg13g2_dlygate4sd3_1 hold1459 (.A(_01020_),
    .X(net3693));
 sg13g2_dlygate4sd3_1 hold1460 (.A(\cpu.arbiter.i_wb_mem_rdt[13] ),
    .X(net3694));
 sg13g2_dlygate4sd3_1 hold1461 (.A(_01025_),
    .X(net3695));
 sg13g2_dlygate4sd3_1 hold1462 (.A(\cpu.cpu.immdec.gen_immdec_w_eq_1.imm30_25[0] ),
    .X(net3696));
 sg13g2_dlygate4sd3_1 hold1463 (.A(\cpu.cpu.bufreg2.i_bytecnt[0] ),
    .X(net3697));
 sg13g2_dlygate4sd3_1 hold1464 (.A(_03654_),
    .X(net3698));
 sg13g2_dlygate4sd3_1 hold1465 (.A(_00475_),
    .X(net3699));
 sg13g2_dlygate4sd3_1 hold1466 (.A(\cpu.arbiter.i_wb_cpu_dbus_adr[10] ),
    .X(net3700));
 sg13g2_dlygate4sd3_1 hold1467 (.A(\cpu.cpu.immdec.gen_immdec_w_eq_1.imm24_20[3] ),
    .X(net3701));
 sg13g2_dlygate4sd3_1 hold1468 (.A(_03762_),
    .X(net3702));
 sg13g2_dlygate4sd3_1 hold1469 (.A(\cpu.arbiter.i_wb_cpu_dbus_adr[4] ),
    .X(net3703));
 sg13g2_dlygate4sd3_1 hold1470 (.A(\ram_spi_if.state_reg[2] ),
    .X(net3704));
 sg13g2_dlygate4sd3_1 hold1471 (.A(_01675_),
    .X(net3705));
 sg13g2_dlygate4sd3_1 hold1472 (.A(_00686_),
    .X(net3706));
 sg13g2_dlygate4sd3_1 hold1473 (.A(\cpu.arbiter.i_wb_mem_rdt[21] ),
    .X(net3707));
 sg13g2_dlygate4sd3_1 hold1474 (.A(_00517_),
    .X(net3708));
 sg13g2_dlygate4sd3_1 hold1475 (.A(\cpu.cpu.immdec.gen_immdec_w_eq_1.imm11_7[2] ),
    .X(net3709));
 sg13g2_dlygate4sd3_1 hold1476 (.A(_03924_),
    .X(net3710));
 sg13g2_dlygate4sd3_1 hold1477 (.A(_00616_),
    .X(net3711));
 sg13g2_dlygate4sd3_1 hold1478 (.A(\cpu.arbiter.i_wb_cpu_dbus_adr[13] ),
    .X(net3712));
 sg13g2_dlygate4sd3_1 hold1479 (.A(\cpu.arbiter.i_wb_mem_rdt[11] ),
    .X(net3713));
 sg13g2_dlygate4sd3_1 hold1480 (.A(\cpu.cpu.immdec.gen_immdec_w_eq_1.imm11_7[3] ),
    .X(net3714));
 sg13g2_dlygate4sd3_1 hold1481 (.A(_03925_),
    .X(net3715));
 sg13g2_dlygate4sd3_1 hold1482 (.A(\cpu.cpu.decode.opcode[0] ),
    .X(net3716));
 sg13g2_dlygate4sd3_1 hold1483 (.A(\ram_spi_if.cycle_counter[5] ),
    .X(net3717));
 sg13g2_dlygate4sd3_1 hold1484 (.A(\cpu.arbiter.i_wb_mem_rdt[4] ),
    .X(net3718));
 sg13g2_dlygate4sd3_1 hold1485 (.A(\cpu.cpu.immdec.gen_immdec_w_eq_1.imm24_20[4] ),
    .X(net3719));
 sg13g2_dlygate4sd3_1 hold1486 (.A(\cpu.cpu.state.init_done ),
    .X(net3720));
 sg13g2_dlygate4sd3_1 hold1487 (.A(\cpu.i_wb_ext_rdt[0] ),
    .X(net3721));
 sg13g2_dlygate4sd3_1 hold1488 (.A(\cpu.cpu.immdec.gen_immdec_w_eq_1.imm11_7[4] ),
    .X(net3722));
 sg13g2_dlygate4sd3_1 hold1489 (.A(\cpu.rf_ram_if.rcnt[4] ),
    .X(net3723));
 sg13g2_dlygate4sd3_1 hold1490 (.A(\cpu.arbiter.i_wb_mem_rdt[9] ),
    .X(net3724));
 sg13g2_dlygate4sd3_1 hold1491 (.A(\ram_spi_if.state_reg[1] ),
    .X(net3725));
 sg13g2_dlygate4sd3_1 hold1492 (.A(\ram_spi_if.state_reg[3] ),
    .X(net3726));
 sg13g2_dlygate4sd3_1 hold1493 (.A(_00687_),
    .X(net3727));
 sg13g2_dlygate4sd3_1 hold1494 (.A(\cpu.arbiter.i_wb_mem_rdt[23] ),
    .X(net3728));
 sg13g2_dlygate4sd3_1 hold1495 (.A(_02714_),
    .X(net3729));
 sg13g2_dlygate4sd3_1 hold1496 (.A(\cpu.cpu.decode.opcode[1] ),
    .X(net3730));
 sg13g2_dlygate4sd3_1 hold1497 (.A(\ram_spi_if.state_reg[0] ),
    .X(net3731));
 sg13g2_dlygate4sd3_1 hold1498 (.A(\cpu.arbiter.i_wb_mem_rdt[30] ),
    .X(net3732));
 sg13g2_dlygate4sd3_1 hold1499 (.A(_00538_),
    .X(net3733));
 sg13g2_dlygate4sd3_1 hold1500 (.A(\cpu.arbiter.i_wb_cpu_dbus_dat[25] ),
    .X(net3734));
 sg13g2_dlygate4sd3_1 hold1501 (.A(_00541_),
    .X(net3735));
 sg13g2_dlygate4sd3_1 hold1502 (.A(\cpu.cpu.decode.opcode[2] ),
    .X(net3736));
 sg13g2_dlygate4sd3_1 hold1503 (.A(\cpu.cpu.branch_op ),
    .X(net3737));
 sg13g2_dlygate4sd3_1 hold1504 (.A(\cpu.arbiter.i_wb_cpu_dbus_dat[8] ),
    .X(net3738));
 sg13g2_dlygate4sd3_1 hold1505 (.A(\cpu.arbiter.i_wb_cpu_dbus_dat[28] ),
    .X(net3739));
 sg13g2_dlygate4sd3_1 hold1506 (.A(_00544_),
    .X(net3740));
 sg13g2_dlygate4sd3_1 hold1507 (.A(\cpu.arbiter.i_wb_mem_rdt[15] ),
    .X(net3741));
 sg13g2_dlygate4sd3_1 hold1508 (.A(\cpu.arbiter.i_wb_cpu_dbus_dat[29] ),
    .X(net3742));
 sg13g2_dlygate4sd3_1 hold1509 (.A(_00545_),
    .X(net3743));
 sg13g2_dlygate4sd3_1 hold1510 (.A(\cpu.arbiter.i_wb_cpu_dbus_adr[31] ),
    .X(net3744));
 sg13g2_dlygate4sd3_1 hold1511 (.A(_00432_),
    .X(net3745));
 sg13g2_dlygate4sd3_1 hold1512 (.A(\cpu.cpu.bufreg.i_right_shift_op ),
    .X(net3746));
 sg13g2_dlygate4sd3_1 hold1513 (.A(\cpu.cpu.bufreg.data[1] ),
    .X(net3747));
 sg13g2_dlygate4sd3_1 hold1514 (.A(_00548_),
    .X(net3748));
 sg13g2_dlygate4sd3_1 hold1515 (.A(\cpu.arbiter.i_wb_mem_rdt[7] ),
    .X(net3749));
 sg13g2_dlygate4sd3_1 hold1516 (.A(_01019_),
    .X(net3750));
 sg13g2_dlygate4sd3_1 hold1517 (.A(\cpu.arbiter.i_wb_cpu_dbus_dat[24] ),
    .X(net3751));
 sg13g2_dlygate4sd3_1 hold1518 (.A(\cpu.arbiter.i_wb_cpu_dbus_dat[26] ),
    .X(net3752));
 sg13g2_dlygate4sd3_1 hold1519 (.A(\cpu.cpu.immdec.gen_immdec_w_eq_1.imm24_20[1] ),
    .X(net3753));
 sg13g2_dlygate4sd3_1 hold1520 (.A(_03760_),
    .X(net3754));
 sg13g2_dlygate4sd3_1 hold1521 (.A(\cpu.rf_ram_if.rgate ),
    .X(net3755));
 sg13g2_dlygate4sd3_1 hold1522 (.A(\ram_spi_if.state_reg[1] ),
    .X(net3756));
 sg13g2_dlygate4sd3_1 hold1523 (.A(\cpu.cpu.bufreg2.i_bytecnt[1] ),
    .X(net3757));
 sg13g2_dlygate4sd3_1 hold1524 (.A(_00476_),
    .X(net3758));
 sg13g2_dlygate4sd3_1 hold1525 (.A(\cpu.rf_ram_if.rcnt[1] ),
    .X(net3759));
 sg13g2_dlygate4sd3_1 hold1526 (.A(\cpu.rf_ram_if.rdata0[22] ),
    .X(net3760));
 sg13g2_dlygate4sd3_1 hold1527 (.A(_00013_),
    .X(net3761));
 sg13g2_dlygate4sd3_1 hold1528 (.A(\cpu.cpu.ctrl.pc_plus_offset_cy_r_w [0]),
    .X(net3762));
 sg13g2_dlygate4sd3_1 hold1529 (.A(_01499_),
    .X(net3763));
 sg13g2_dlygate4sd3_1 hold1530 (.A(\cpu.cpu.alu.add_cy_r [0]),
    .X(net3764));
 sg13g2_dlygate4sd3_1 hold1531 (.A(_01421_),
    .X(net3765));
 sg13g2_dlygate4sd3_1 hold1532 (.A(_00061_),
    .X(net3766));
 sg13g2_dlygate4sd3_1 hold1533 (.A(\cpu.rf_ram_if.rcnt[4] ),
    .X(net3767));
 sg13g2_dlygate4sd3_1 hold1534 (.A(_01402_),
    .X(net3768));
 sg13g2_dlygate4sd3_1 hold1535 (.A(_02808_),
    .X(net3769));
 sg13g2_dlygate4sd3_1 hold1536 (.A(\rf_ram.RAM[19][6] ),
    .X(net3770));
 sg13g2_dlygate4sd3_1 hold1537 (.A(\rf_ram.RAM[11][12] ),
    .X(net3771));
 sg13g2_dlygate4sd3_1 hold1538 (.A(_03146_),
    .X(net3772));
 sg13g2_dlygate4sd3_1 hold1539 (.A(\rf_ram.RAM[23][1] ),
    .X(net3773));
 sg13g2_dlygate4sd3_1 hold1540 (.A(\rf_ram.RAM[7][8] ),
    .X(net3774));
 sg13g2_dlygate4sd3_1 hold1541 (.A(\rf_ram.RAM[7][25] ),
    .X(net3775));
 sg13g2_dlygate4sd3_1 hold1542 (.A(\rf_ram.RAM[7][17] ),
    .X(net3776));
 sg13g2_dlygate4sd3_1 hold1543 (.A(\rf_ram.RAM[7][10] ),
    .X(net3777));
 sg13g2_dlygate4sd3_1 hold1544 (.A(_03094_),
    .X(net3778));
 sg13g2_dlygate4sd3_1 hold1545 (.A(\rf_ram.RAM[27][7] ),
    .X(net3779));
 sg13g2_dlygate4sd3_1 hold1546 (.A(_03016_),
    .X(net3780));
 sg13g2_dlygate4sd3_1 hold1547 (.A(\rf_ram.RAM[25][23] ),
    .X(net3781));
 sg13g2_dlygate4sd3_1 hold1548 (.A(\rf_ram.RAM[11][16] ),
    .X(net3782));
 sg13g2_dlygate4sd3_1 hold1549 (.A(_03249_),
    .X(net3783));
 sg13g2_dlygate4sd3_1 hold1550 (.A(_00449_),
    .X(net3784));
 sg13g2_dlygate4sd3_1 hold1551 (.A(\rf_ram.RAM[3][4] ),
    .X(net3785));
 sg13g2_dlygate4sd3_1 hold1552 (.A(_02938_),
    .X(net3786));
 sg13g2_dlygate4sd3_1 hold1553 (.A(_00437_),
    .X(net3787));
 sg13g2_dlygate4sd3_1 hold1554 (.A(\rf_ram.RAM[15][28] ),
    .X(net3788));
 sg13g2_dlygate4sd3_1 hold1555 (.A(\rf_ram.RAM[19][22] ),
    .X(net3789));
 sg13g2_dlygate4sd3_1 hold1556 (.A(\rf_ram.RAM[23][18] ),
    .X(net3790));
 sg13g2_dlygate4sd3_1 hold1557 (.A(_03302_),
    .X(net3791));
 sg13g2_dlygate4sd3_1 hold1558 (.A(_00451_),
    .X(net3792));
 sg13g2_dlygate4sd3_1 hold1559 (.A(\rf_ram.RAM[31][0] ),
    .X(net3793));
 sg13g2_dlygate4sd3_1 hold1560 (.A(\rf_ram.RAM[7][26] ),
    .X(net3794));
 sg13g2_dlygate4sd3_1 hold1561 (.A(_00459_),
    .X(net3795));
 sg13g2_dlygate4sd3_1 hold1562 (.A(\rf_ram.RAM[15][3] ),
    .X(net3796));
 sg13g2_dlygate4sd3_1 hold1563 (.A(_00436_),
    .X(net3797));
 sg13g2_dlygate4sd3_1 hold1564 (.A(\rf_ram.RAM[15][5] ),
    .X(net3798));
 sg13g2_dlygate4sd3_1 hold1565 (.A(_02964_),
    .X(net3799));
 sg13g2_dlygate4sd3_1 hold1566 (.A(\rf_ram.RAM[9][9] ),
    .X(net3800));
 sg13g2_dlygate4sd3_1 hold1567 (.A(_03068_),
    .X(net3801));
 sg13g2_dlygate4sd3_1 hold1568 (.A(_00442_),
    .X(net3802));
 sg13g2_dlygate4sd3_1 hold1569 (.A(\rf_ram.RAM[3][31] ),
    .X(net3803));
 sg13g2_dlygate4sd3_1 hold1570 (.A(_03629_),
    .X(net3804));
 sg13g2_dlygate4sd3_1 hold1571 (.A(_03639_),
    .X(net3805));
 sg13g2_dlygate4sd3_1 hold1572 (.A(_00464_),
    .X(net3806));
 sg13g2_dlygate4sd3_1 hold1573 (.A(\rf_ram.RAM[30][19] ),
    .X(net3807));
 sg13g2_dlygate4sd3_1 hold1574 (.A(_03327_),
    .X(net3808));
 sg13g2_dlygate4sd3_1 hold1575 (.A(_00452_),
    .X(net3809));
 sg13g2_dlygate4sd3_1 hold1576 (.A(\rf_ram.RAM[8][2] ),
    .X(net3810));
 sg13g2_dlygate4sd3_1 hold1577 (.A(_02884_),
    .X(net3811));
 sg13g2_dlygate4sd3_1 hold1578 (.A(_02885_),
    .X(net3812));
 sg13g2_dlygate4sd3_1 hold1579 (.A(\rf_ram.RAM[25][30] ),
    .X(net3813));
 sg13g2_dlygate4sd3_1 hold1580 (.A(_03609_),
    .X(net3814));
 sg13g2_dlygate4sd3_1 hold1581 (.A(_03613_),
    .X(net3815));
 sg13g2_dlygate4sd3_1 hold1582 (.A(\rf_ram.RAM[22][14] ),
    .X(net3816));
 sg13g2_dlygate4sd3_1 hold1583 (.A(_03197_),
    .X(net3817));
 sg13g2_dlygate4sd3_1 hold1584 (.A(\cpu.rf_ram_if.rcnt[1] ),
    .X(net3818));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_fill_2 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_71 ();
 sg13g2_decap_8 FILLER_0_78 ();
 sg13g2_fill_2 FILLER_0_85 ();
 sg13g2_fill_1 FILLER_0_87 ();
 sg13g2_fill_1 FILLER_0_92 ();
 sg13g2_fill_1 FILLER_0_112 ();
 sg13g2_fill_2 FILLER_0_122 ();
 sg13g2_decap_8 FILLER_0_143 ();
 sg13g2_decap_8 FILLER_0_150 ();
 sg13g2_decap_8 FILLER_0_157 ();
 sg13g2_decap_8 FILLER_0_164 ();
 sg13g2_decap_8 FILLER_0_171 ();
 sg13g2_decap_4 FILLER_0_178 ();
 sg13g2_fill_1 FILLER_0_182 ();
 sg13g2_fill_1 FILLER_0_187 ();
 sg13g2_decap_8 FILLER_0_201 ();
 sg13g2_decap_8 FILLER_0_208 ();
 sg13g2_fill_2 FILLER_0_215 ();
 sg13g2_fill_2 FILLER_0_221 ();
 sg13g2_fill_1 FILLER_0_223 ();
 sg13g2_decap_4 FILLER_0_246 ();
 sg13g2_decap_8 FILLER_0_254 ();
 sg13g2_decap_8 FILLER_0_261 ();
 sg13g2_decap_8 FILLER_0_268 ();
 sg13g2_decap_8 FILLER_0_275 ();
 sg13g2_fill_2 FILLER_0_282 ();
 sg13g2_decap_8 FILLER_0_288 ();
 sg13g2_decap_8 FILLER_0_295 ();
 sg13g2_decap_8 FILLER_0_302 ();
 sg13g2_decap_8 FILLER_0_340 ();
 sg13g2_decap_8 FILLER_0_347 ();
 sg13g2_decap_8 FILLER_0_354 ();
 sg13g2_decap_4 FILLER_0_361 ();
 sg13g2_fill_2 FILLER_0_369 ();
 sg13g2_fill_1 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_381 ();
 sg13g2_decap_8 FILLER_0_415 ();
 sg13g2_fill_2 FILLER_0_422 ();
 sg13g2_decap_4 FILLER_0_428 ();
 sg13g2_fill_1 FILLER_0_432 ();
 sg13g2_decap_8 FILLER_0_445 ();
 sg13g2_decap_8 FILLER_0_452 ();
 sg13g2_decap_8 FILLER_0_459 ();
 sg13g2_decap_8 FILLER_0_466 ();
 sg13g2_decap_8 FILLER_0_473 ();
 sg13g2_decap_4 FILLER_0_480 ();
 sg13g2_decap_4 FILLER_0_489 ();
 sg13g2_fill_1 FILLER_0_493 ();
 sg13g2_decap_8 FILLER_0_498 ();
 sg13g2_decap_8 FILLER_0_505 ();
 sg13g2_decap_8 FILLER_0_512 ();
 sg13g2_decap_8 FILLER_0_519 ();
 sg13g2_decap_8 FILLER_0_526 ();
 sg13g2_decap_8 FILLER_0_533 ();
 sg13g2_decap_8 FILLER_0_540 ();
 sg13g2_decap_4 FILLER_0_547 ();
 sg13g2_fill_1 FILLER_0_551 ();
 sg13g2_fill_2 FILLER_0_565 ();
 sg13g2_fill_1 FILLER_0_567 ();
 sg13g2_decap_8 FILLER_0_591 ();
 sg13g2_fill_1 FILLER_0_598 ();
 sg13g2_fill_1 FILLER_0_615 ();
 sg13g2_decap_8 FILLER_0_625 ();
 sg13g2_decap_8 FILLER_0_632 ();
 sg13g2_decap_8 FILLER_0_639 ();
 sg13g2_decap_8 FILLER_0_646 ();
 sg13g2_decap_8 FILLER_0_653 ();
 sg13g2_decap_8 FILLER_0_660 ();
 sg13g2_decap_8 FILLER_0_667 ();
 sg13g2_decap_8 FILLER_0_674 ();
 sg13g2_decap_8 FILLER_0_681 ();
 sg13g2_decap_8 FILLER_0_688 ();
 sg13g2_decap_8 FILLER_0_695 ();
 sg13g2_decap_4 FILLER_0_702 ();
 sg13g2_fill_1 FILLER_0_706 ();
 sg13g2_decap_8 FILLER_0_711 ();
 sg13g2_decap_8 FILLER_0_718 ();
 sg13g2_decap_8 FILLER_0_725 ();
 sg13g2_decap_8 FILLER_0_732 ();
 sg13g2_decap_8 FILLER_0_743 ();
 sg13g2_decap_8 FILLER_0_750 ();
 sg13g2_decap_8 FILLER_0_757 ();
 sg13g2_decap_8 FILLER_0_764 ();
 sg13g2_decap_8 FILLER_0_771 ();
 sg13g2_decap_8 FILLER_0_778 ();
 sg13g2_decap_8 FILLER_0_785 ();
 sg13g2_decap_8 FILLER_0_792 ();
 sg13g2_decap_8 FILLER_0_799 ();
 sg13g2_decap_8 FILLER_0_806 ();
 sg13g2_decap_8 FILLER_0_813 ();
 sg13g2_decap_4 FILLER_0_820 ();
 sg13g2_fill_2 FILLER_0_824 ();
 sg13g2_decap_8 FILLER_0_830 ();
 sg13g2_decap_8 FILLER_0_837 ();
 sg13g2_decap_8 FILLER_0_844 ();
 sg13g2_decap_8 FILLER_0_851 ();
 sg13g2_decap_8 FILLER_0_858 ();
 sg13g2_decap_4 FILLER_0_865 ();
 sg13g2_fill_2 FILLER_0_869 ();
 sg13g2_decap_4 FILLER_0_898 ();
 sg13g2_fill_2 FILLER_0_902 ();
 sg13g2_decap_8 FILLER_0_908 ();
 sg13g2_decap_8 FILLER_0_915 ();
 sg13g2_decap_8 FILLER_0_922 ();
 sg13g2_decap_8 FILLER_0_929 ();
 sg13g2_decap_8 FILLER_0_936 ();
 sg13g2_decap_8 FILLER_0_943 ();
 sg13g2_decap_4 FILLER_0_950 ();
 sg13g2_fill_2 FILLER_0_954 ();
 sg13g2_decap_4 FILLER_0_960 ();
 sg13g2_fill_2 FILLER_0_964 ();
 sg13g2_decap_8 FILLER_0_970 ();
 sg13g2_decap_8 FILLER_0_977 ();
 sg13g2_decap_8 FILLER_0_984 ();
 sg13g2_decap_8 FILLER_0_991 ();
 sg13g2_fill_2 FILLER_0_998 ();
 sg13g2_fill_1 FILLER_0_1000 ();
 sg13g2_fill_2 FILLER_0_1019 ();
 sg13g2_fill_1 FILLER_0_1021 ();
 sg13g2_fill_2 FILLER_0_1036 ();
 sg13g2_fill_1 FILLER_0_1038 ();
 sg13g2_decap_8 FILLER_0_1061 ();
 sg13g2_decap_8 FILLER_0_1068 ();
 sg13g2_decap_8 FILLER_0_1075 ();
 sg13g2_decap_8 FILLER_0_1082 ();
 sg13g2_fill_2 FILLER_0_1089 ();
 sg13g2_decap_8 FILLER_0_1096 ();
 sg13g2_decap_8 FILLER_0_1103 ();
 sg13g2_decap_8 FILLER_0_1110 ();
 sg13g2_decap_4 FILLER_0_1117 ();
 sg13g2_fill_1 FILLER_0_1121 ();
 sg13g2_fill_1 FILLER_0_1126 ();
 sg13g2_decap_8 FILLER_0_1131 ();
 sg13g2_decap_8 FILLER_0_1138 ();
 sg13g2_decap_4 FILLER_0_1145 ();
 sg13g2_fill_2 FILLER_0_1149 ();
 sg13g2_decap_4 FILLER_0_1155 ();
 sg13g2_fill_2 FILLER_0_1159 ();
 sg13g2_decap_8 FILLER_0_1174 ();
 sg13g2_decap_8 FILLER_0_1181 ();
 sg13g2_decap_8 FILLER_0_1188 ();
 sg13g2_decap_8 FILLER_0_1195 ();
 sg13g2_decap_8 FILLER_0_1202 ();
 sg13g2_decap_8 FILLER_0_1209 ();
 sg13g2_decap_8 FILLER_0_1216 ();
 sg13g2_decap_8 FILLER_0_1223 ();
 sg13g2_decap_8 FILLER_0_1230 ();
 sg13g2_decap_8 FILLER_0_1237 ();
 sg13g2_decap_8 FILLER_0_1244 ();
 sg13g2_decap_8 FILLER_0_1251 ();
 sg13g2_decap_8 FILLER_0_1258 ();
 sg13g2_decap_8 FILLER_0_1265 ();
 sg13g2_decap_8 FILLER_0_1272 ();
 sg13g2_decap_8 FILLER_0_1279 ();
 sg13g2_decap_8 FILLER_0_1286 ();
 sg13g2_decap_8 FILLER_0_1293 ();
 sg13g2_decap_8 FILLER_0_1300 ();
 sg13g2_decap_8 FILLER_0_1307 ();
 sg13g2_fill_1 FILLER_0_1314 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_fill_1 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_73 ();
 sg13g2_fill_2 FILLER_1_80 ();
 sg13g2_fill_1 FILLER_1_82 ();
 sg13g2_decap_8 FILLER_1_146 ();
 sg13g2_decap_8 FILLER_1_153 ();
 sg13g2_decap_8 FILLER_1_160 ();
 sg13g2_fill_2 FILLER_1_194 ();
 sg13g2_fill_1 FILLER_1_200 ();
 sg13g2_fill_1 FILLER_1_273 ();
 sg13g2_fill_2 FILLER_1_310 ();
 sg13g2_fill_1 FILLER_1_312 ();
 sg13g2_fill_2 FILLER_1_376 ();
 sg13g2_fill_2 FILLER_1_405 ();
 sg13g2_fill_2 FILLER_1_461 ();
 sg13g2_fill_1 FILLER_1_463 ();
 sg13g2_fill_1 FILLER_1_469 ();
 sg13g2_decap_4 FILLER_1_474 ();
 sg13g2_fill_2 FILLER_1_478 ();
 sg13g2_decap_4 FILLER_1_520 ();
 sg13g2_fill_2 FILLER_1_524 ();
 sg13g2_fill_1 FILLER_1_589 ();
 sg13g2_fill_2 FILLER_1_631 ();
 sg13g2_decap_8 FILLER_1_660 ();
 sg13g2_decap_4 FILLER_1_671 ();
 sg13g2_fill_1 FILLER_1_675 ();
 sg13g2_fill_2 FILLER_1_724 ();
 sg13g2_fill_1 FILLER_1_726 ();
 sg13g2_fill_1 FILLER_1_763 ();
 sg13g2_decap_8 FILLER_1_795 ();
 sg13g2_decap_8 FILLER_1_802 ();
 sg13g2_fill_1 FILLER_1_809 ();
 sg13g2_decap_8 FILLER_1_854 ();
 sg13g2_fill_2 FILLER_1_861 ();
 sg13g2_fill_2 FILLER_1_890 ();
 sg13g2_fill_2 FILLER_1_901 ();
 sg13g2_fill_1 FILLER_1_903 ();
 sg13g2_decap_8 FILLER_1_935 ();
 sg13g2_fill_1 FILLER_1_982 ();
 sg13g2_decap_8 FILLER_1_992 ();
 sg13g2_fill_2 FILLER_1_999 ();
 sg13g2_fill_2 FILLER_1_1028 ();
 sg13g2_decap_4 FILLER_1_1079 ();
 sg13g2_fill_2 FILLER_1_1083 ();
 sg13g2_decap_4 FILLER_1_1094 ();
 sg13g2_decap_8 FILLER_1_1138 ();
 sg13g2_fill_2 FILLER_1_1145 ();
 sg13g2_decap_8 FILLER_1_1178 ();
 sg13g2_decap_8 FILLER_1_1185 ();
 sg13g2_decap_8 FILLER_1_1192 ();
 sg13g2_decap_8 FILLER_1_1199 ();
 sg13g2_decap_8 FILLER_1_1206 ();
 sg13g2_decap_8 FILLER_1_1213 ();
 sg13g2_decap_8 FILLER_1_1220 ();
 sg13g2_decap_8 FILLER_1_1227 ();
 sg13g2_decap_8 FILLER_1_1234 ();
 sg13g2_decap_8 FILLER_1_1241 ();
 sg13g2_decap_8 FILLER_1_1248 ();
 sg13g2_decap_8 FILLER_1_1255 ();
 sg13g2_decap_8 FILLER_1_1262 ();
 sg13g2_decap_8 FILLER_1_1269 ();
 sg13g2_decap_8 FILLER_1_1276 ();
 sg13g2_decap_8 FILLER_1_1283 ();
 sg13g2_decap_8 FILLER_1_1290 ();
 sg13g2_decap_8 FILLER_1_1297 ();
 sg13g2_decap_8 FILLER_1_1304 ();
 sg13g2_decap_4 FILLER_1_1311 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_4 FILLER_2_21 ();
 sg13g2_fill_2 FILLER_2_25 ();
 sg13g2_fill_1 FILLER_2_68 ();
 sg13g2_fill_2 FILLER_2_78 ();
 sg13g2_fill_2 FILLER_2_117 ();
 sg13g2_fill_1 FILLER_2_133 ();
 sg13g2_fill_2 FILLER_2_161 ();
 sg13g2_fill_1 FILLER_2_163 ();
 sg13g2_fill_1 FILLER_2_260 ();
 sg13g2_fill_2 FILLER_2_302 ();
 sg13g2_fill_1 FILLER_2_326 ();
 sg13g2_fill_2 FILLER_2_344 ();
 sg13g2_fill_1 FILLER_2_377 ();
 sg13g2_fill_1 FILLER_2_387 ();
 sg13g2_fill_1 FILLER_2_397 ();
 sg13g2_fill_1 FILLER_2_402 ();
 sg13g2_fill_2 FILLER_2_416 ();
 sg13g2_fill_1 FILLER_2_418 ();
 sg13g2_fill_2 FILLER_2_433 ();
 sg13g2_fill_1 FILLER_2_435 ();
 sg13g2_fill_2 FILLER_2_458 ();
 sg13g2_fill_1 FILLER_2_460 ();
 sg13g2_fill_2 FILLER_2_515 ();
 sg13g2_fill_1 FILLER_2_526 ();
 sg13g2_fill_2 FILLER_2_556 ();
 sg13g2_fill_1 FILLER_2_558 ();
 sg13g2_fill_2 FILLER_2_599 ();
 sg13g2_fill_2 FILLER_2_628 ();
 sg13g2_fill_1 FILLER_2_730 ();
 sg13g2_fill_1 FILLER_2_758 ();
 sg13g2_fill_2 FILLER_2_885 ();
 sg13g2_fill_1 FILLER_2_928 ();
 sg13g2_fill_2 FILLER_2_1010 ();
 sg13g2_fill_1 FILLER_2_1012 ();
 sg13g2_fill_1 FILLER_2_1055 ();
 sg13g2_decap_8 FILLER_2_1186 ();
 sg13g2_fill_2 FILLER_2_1193 ();
 sg13g2_fill_1 FILLER_2_1195 ();
 sg13g2_decap_8 FILLER_2_1204 ();
 sg13g2_decap_8 FILLER_2_1211 ();
 sg13g2_decap_8 FILLER_2_1218 ();
 sg13g2_decap_8 FILLER_2_1225 ();
 sg13g2_decap_8 FILLER_2_1232 ();
 sg13g2_decap_8 FILLER_2_1239 ();
 sg13g2_decap_8 FILLER_2_1246 ();
 sg13g2_decap_8 FILLER_2_1253 ();
 sg13g2_decap_8 FILLER_2_1260 ();
 sg13g2_decap_8 FILLER_2_1267 ();
 sg13g2_decap_8 FILLER_2_1274 ();
 sg13g2_decap_8 FILLER_2_1281 ();
 sg13g2_decap_8 FILLER_2_1288 ();
 sg13g2_decap_8 FILLER_2_1295 ();
 sg13g2_decap_8 FILLER_2_1302 ();
 sg13g2_decap_4 FILLER_2_1309 ();
 sg13g2_fill_2 FILLER_2_1313 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_4 FILLER_3_14 ();
 sg13g2_fill_2 FILLER_3_202 ();
 sg13g2_fill_2 FILLER_3_272 ();
 sg13g2_fill_1 FILLER_3_274 ();
 sg13g2_fill_1 FILLER_3_284 ();
 sg13g2_fill_1 FILLER_3_291 ();
 sg13g2_fill_2 FILLER_3_305 ();
 sg13g2_fill_2 FILLER_3_344 ();
 sg13g2_fill_1 FILLER_3_346 ();
 sg13g2_fill_1 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_fill_2 FILLER_3_385 ();
 sg13g2_fill_2 FILLER_3_396 ();
 sg13g2_fill_1 FILLER_3_398 ();
 sg13g2_fill_2 FILLER_3_463 ();
 sg13g2_fill_1 FILLER_3_465 ();
 sg13g2_fill_2 FILLER_3_493 ();
 sg13g2_fill_1 FILLER_3_495 ();
 sg13g2_fill_2 FILLER_3_502 ();
 sg13g2_fill_1 FILLER_3_504 ();
 sg13g2_decap_4 FILLER_3_524 ();
 sg13g2_fill_1 FILLER_3_528 ();
 sg13g2_decap_4 FILLER_3_533 ();
 sg13g2_fill_2 FILLER_3_587 ();
 sg13g2_fill_1 FILLER_3_589 ();
 sg13g2_fill_2 FILLER_3_623 ();
 sg13g2_fill_1 FILLER_3_625 ();
 sg13g2_fill_2 FILLER_3_679 ();
 sg13g2_fill_1 FILLER_3_686 ();
 sg13g2_fill_2 FILLER_3_742 ();
 sg13g2_fill_1 FILLER_3_772 ();
 sg13g2_fill_1 FILLER_3_786 ();
 sg13g2_fill_2 FILLER_3_823 ();
 sg13g2_fill_1 FILLER_3_875 ();
 sg13g2_fill_2 FILLER_3_880 ();
 sg13g2_fill_2 FILLER_3_905 ();
 sg13g2_fill_1 FILLER_3_1064 ();
 sg13g2_fill_1 FILLER_3_1106 ();
 sg13g2_decap_8 FILLER_3_1234 ();
 sg13g2_decap_8 FILLER_3_1241 ();
 sg13g2_decap_8 FILLER_3_1248 ();
 sg13g2_decap_4 FILLER_3_1255 ();
 sg13g2_fill_1 FILLER_3_1259 ();
 sg13g2_decap_8 FILLER_3_1268 ();
 sg13g2_decap_8 FILLER_3_1275 ();
 sg13g2_decap_8 FILLER_3_1282 ();
 sg13g2_decap_8 FILLER_3_1289 ();
 sg13g2_decap_8 FILLER_3_1296 ();
 sg13g2_decap_8 FILLER_3_1303 ();
 sg13g2_decap_4 FILLER_3_1310 ();
 sg13g2_fill_1 FILLER_3_1314 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_fill_2 FILLER_4_7 ();
 sg13g2_fill_1 FILLER_4_9 ();
 sg13g2_decap_4 FILLER_4_79 ();
 sg13g2_fill_1 FILLER_4_83 ();
 sg13g2_fill_2 FILLER_4_107 ();
 sg13g2_decap_4 FILLER_4_161 ();
 sg13g2_fill_2 FILLER_4_192 ();
 sg13g2_fill_2 FILLER_4_230 ();
 sg13g2_fill_1 FILLER_4_232 ();
 sg13g2_fill_1 FILLER_4_242 ();
 sg13g2_fill_2 FILLER_4_256 ();
 sg13g2_fill_2 FILLER_4_282 ();
 sg13g2_fill_1 FILLER_4_284 ();
 sg13g2_decap_4 FILLER_4_289 ();
 sg13g2_fill_2 FILLER_4_293 ();
 sg13g2_decap_8 FILLER_4_304 ();
 sg13g2_fill_2 FILLER_4_347 ();
 sg13g2_decap_4 FILLER_4_353 ();
 sg13g2_fill_2 FILLER_4_357 ();
 sg13g2_fill_2 FILLER_4_386 ();
 sg13g2_fill_1 FILLER_4_388 ();
 sg13g2_fill_1 FILLER_4_426 ();
 sg13g2_fill_2 FILLER_4_454 ();
 sg13g2_fill_1 FILLER_4_456 ();
 sg13g2_fill_2 FILLER_4_466 ();
 sg13g2_fill_1 FILLER_4_468 ();
 sg13g2_fill_1 FILLER_4_539 ();
 sg13g2_fill_2 FILLER_4_567 ();
 sg13g2_decap_4 FILLER_4_582 ();
 sg13g2_fill_2 FILLER_4_627 ();
 sg13g2_fill_1 FILLER_4_629 ();
 sg13g2_fill_2 FILLER_4_677 ();
 sg13g2_fill_1 FILLER_4_771 ();
 sg13g2_fill_1 FILLER_4_777 ();
 sg13g2_fill_2 FILLER_4_793 ();
 sg13g2_fill_2 FILLER_4_805 ();
 sg13g2_fill_1 FILLER_4_807 ();
 sg13g2_fill_2 FILLER_4_828 ();
 sg13g2_fill_2 FILLER_4_949 ();
 sg13g2_fill_2 FILLER_4_971 ();
 sg13g2_fill_1 FILLER_4_1023 ();
 sg13g2_fill_1 FILLER_4_1050 ();
 sg13g2_decap_8 FILLER_4_1055 ();
 sg13g2_decap_4 FILLER_4_1062 ();
 sg13g2_fill_1 FILLER_4_1094 ();
 sg13g2_fill_2 FILLER_4_1099 ();
 sg13g2_fill_1 FILLER_4_1190 ();
 sg13g2_fill_2 FILLER_4_1196 ();
 sg13g2_fill_1 FILLER_4_1198 ();
 sg13g2_decap_4 FILLER_4_1240 ();
 sg13g2_fill_2 FILLER_4_1244 ();
 sg13g2_fill_2 FILLER_4_1250 ();
 sg13g2_fill_1 FILLER_4_1252 ();
 sg13g2_decap_8 FILLER_4_1280 ();
 sg13g2_decap_8 FILLER_4_1287 ();
 sg13g2_decap_8 FILLER_4_1294 ();
 sg13g2_decap_8 FILLER_4_1301 ();
 sg13g2_decap_8 FILLER_4_1308 ();
 sg13g2_fill_1 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_85 ();
 sg13g2_decap_8 FILLER_5_92 ();
 sg13g2_fill_1 FILLER_5_99 ();
 sg13g2_decap_4 FILLER_5_158 ();
 sg13g2_fill_2 FILLER_5_162 ();
 sg13g2_fill_2 FILLER_5_251 ();
 sg13g2_decap_4 FILLER_5_262 ();
 sg13g2_fill_2 FILLER_5_266 ();
 sg13g2_decap_4 FILLER_5_301 ();
 sg13g2_fill_1 FILLER_5_305 ();
 sg13g2_decap_4 FILLER_5_351 ();
 sg13g2_fill_1 FILLER_5_355 ();
 sg13g2_decap_4 FILLER_5_396 ();
 sg13g2_fill_2 FILLER_5_432 ();
 sg13g2_fill_2 FILLER_5_444 ();
 sg13g2_fill_1 FILLER_5_446 ();
 sg13g2_decap_4 FILLER_5_460 ();
 sg13g2_fill_1 FILLER_5_464 ();
 sg13g2_fill_1 FILLER_5_469 ();
 sg13g2_decap_4 FILLER_5_483 ();
 sg13g2_fill_2 FILLER_5_487 ();
 sg13g2_decap_8 FILLER_5_498 ();
 sg13g2_fill_1 FILLER_5_505 ();
 sg13g2_fill_1 FILLER_5_549 ();
 sg13g2_fill_1 FILLER_5_563 ();
 sg13g2_decap_8 FILLER_5_573 ();
 sg13g2_decap_8 FILLER_5_580 ();
 sg13g2_decap_8 FILLER_5_623 ();
 sg13g2_fill_2 FILLER_5_630 ();
 sg13g2_fill_1 FILLER_5_632 ();
 sg13g2_decap_4 FILLER_5_669 ();
 sg13g2_decap_4 FILLER_5_682 ();
 sg13g2_fill_1 FILLER_5_690 ();
 sg13g2_fill_2 FILLER_5_723 ();
 sg13g2_fill_1 FILLER_5_725 ();
 sg13g2_fill_1 FILLER_5_766 ();
 sg13g2_fill_1 FILLER_5_871 ();
 sg13g2_fill_2 FILLER_5_899 ();
 sg13g2_fill_2 FILLER_5_918 ();
 sg13g2_fill_2 FILLER_5_933 ();
 sg13g2_fill_2 FILLER_5_961 ();
 sg13g2_fill_1 FILLER_5_963 ();
 sg13g2_fill_2 FILLER_5_968 ();
 sg13g2_fill_2 FILLER_5_975 ();
 sg13g2_fill_1 FILLER_5_977 ();
 sg13g2_fill_2 FILLER_5_999 ();
 sg13g2_fill_1 FILLER_5_1001 ();
 sg13g2_fill_2 FILLER_5_1024 ();
 sg13g2_fill_1 FILLER_5_1026 ();
 sg13g2_decap_8 FILLER_5_1044 ();
 sg13g2_decap_8 FILLER_5_1051 ();
 sg13g2_decap_8 FILLER_5_1058 ();
 sg13g2_decap_8 FILLER_5_1065 ();
 sg13g2_decap_4 FILLER_5_1072 ();
 sg13g2_fill_2 FILLER_5_1076 ();
 sg13g2_decap_8 FILLER_5_1091 ();
 sg13g2_decap_4 FILLER_5_1098 ();
 sg13g2_fill_2 FILLER_5_1102 ();
 sg13g2_decap_4 FILLER_5_1108 ();
 sg13g2_fill_2 FILLER_5_1116 ();
 sg13g2_fill_1 FILLER_5_1118 ();
 sg13g2_fill_1 FILLER_5_1128 ();
 sg13g2_fill_2 FILLER_5_1149 ();
 sg13g2_fill_2 FILLER_5_1183 ();
 sg13g2_fill_1 FILLER_5_1185 ();
 sg13g2_fill_1 FILLER_5_1213 ();
 sg13g2_fill_1 FILLER_5_1254 ();
 sg13g2_decap_8 FILLER_5_1291 ();
 sg13g2_decap_8 FILLER_5_1298 ();
 sg13g2_decap_8 FILLER_5_1305 ();
 sg13g2_fill_2 FILLER_5_1312 ();
 sg13g2_fill_1 FILLER_5_1314 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_fill_1 FILLER_6_38 ();
 sg13g2_fill_1 FILLER_6_83 ();
 sg13g2_fill_2 FILLER_6_121 ();
 sg13g2_decap_8 FILLER_6_145 ();
 sg13g2_decap_8 FILLER_6_152 ();
 sg13g2_decap_8 FILLER_6_159 ();
 sg13g2_decap_8 FILLER_6_166 ();
 sg13g2_fill_1 FILLER_6_173 ();
 sg13g2_decap_8 FILLER_6_178 ();
 sg13g2_fill_2 FILLER_6_185 ();
 sg13g2_fill_1 FILLER_6_187 ();
 sg13g2_decap_4 FILLER_6_207 ();
 sg13g2_fill_1 FILLER_6_211 ();
 sg13g2_decap_8 FILLER_6_256 ();
 sg13g2_decap_4 FILLER_6_263 ();
 sg13g2_fill_2 FILLER_6_267 ();
 sg13g2_decap_4 FILLER_6_305 ();
 sg13g2_fill_2 FILLER_6_309 ();
 sg13g2_fill_1 FILLER_6_348 ();
 sg13g2_fill_1 FILLER_6_353 ();
 sg13g2_fill_1 FILLER_6_371 ();
 sg13g2_fill_2 FILLER_6_395 ();
 sg13g2_decap_8 FILLER_6_468 ();
 sg13g2_decap_4 FILLER_6_488 ();
 sg13g2_fill_1 FILLER_6_538 ();
 sg13g2_decap_8 FILLER_6_566 ();
 sg13g2_decap_8 FILLER_6_573 ();
 sg13g2_fill_1 FILLER_6_580 ();
 sg13g2_decap_8 FILLER_6_608 ();
 sg13g2_decap_4 FILLER_6_615 ();
 sg13g2_fill_2 FILLER_6_619 ();
 sg13g2_decap_8 FILLER_6_625 ();
 sg13g2_fill_2 FILLER_6_632 ();
 sg13g2_fill_2 FILLER_6_651 ();
 sg13g2_fill_1 FILLER_6_653 ();
 sg13g2_decap_8 FILLER_6_659 ();
 sg13g2_decap_8 FILLER_6_666 ();
 sg13g2_fill_2 FILLER_6_673 ();
 sg13g2_decap_8 FILLER_6_679 ();
 sg13g2_fill_1 FILLER_6_735 ();
 sg13g2_fill_1 FILLER_6_760 ();
 sg13g2_fill_2 FILLER_6_770 ();
 sg13g2_fill_1 FILLER_6_772 ();
 sg13g2_fill_2 FILLER_6_809 ();
 sg13g2_fill_2 FILLER_6_860 ();
 sg13g2_fill_2 FILLER_6_866 ();
 sg13g2_decap_4 FILLER_6_872 ();
 sg13g2_fill_2 FILLER_6_876 ();
 sg13g2_fill_2 FILLER_6_888 ();
 sg13g2_fill_1 FILLER_6_890 ();
 sg13g2_fill_2 FILLER_6_897 ();
 sg13g2_fill_1 FILLER_6_908 ();
 sg13g2_fill_2 FILLER_6_945 ();
 sg13g2_decap_8 FILLER_6_960 ();
 sg13g2_decap_4 FILLER_6_967 ();
 sg13g2_decap_4 FILLER_6_998 ();
 sg13g2_decap_8 FILLER_6_1011 ();
 sg13g2_fill_1 FILLER_6_1050 ();
 sg13g2_fill_2 FILLER_6_1115 ();
 sg13g2_fill_1 FILLER_6_1117 ();
 sg13g2_decap_8 FILLER_6_1145 ();
 sg13g2_fill_2 FILLER_6_1152 ();
 sg13g2_fill_2 FILLER_6_1185 ();
 sg13g2_fill_1 FILLER_6_1191 ();
 sg13g2_fill_1 FILLER_6_1225 ();
 sg13g2_decap_4 FILLER_6_1241 ();
 sg13g2_fill_1 FILLER_6_1255 ();
 sg13g2_fill_2 FILLER_6_1261 ();
 sg13g2_fill_1 FILLER_6_1263 ();
 sg13g2_decap_8 FILLER_6_1291 ();
 sg13g2_decap_8 FILLER_6_1298 ();
 sg13g2_decap_8 FILLER_6_1305 ();
 sg13g2_fill_2 FILLER_6_1312 ();
 sg13g2_fill_1 FILLER_6_1314 ();
 sg13g2_fill_1 FILLER_7_26 ();
 sg13g2_fill_2 FILLER_7_45 ();
 sg13g2_fill_2 FILLER_7_105 ();
 sg13g2_fill_1 FILLER_7_107 ();
 sg13g2_fill_1 FILLER_7_122 ();
 sg13g2_fill_2 FILLER_7_127 ();
 sg13g2_fill_2 FILLER_7_143 ();
 sg13g2_fill_1 FILLER_7_145 ();
 sg13g2_decap_8 FILLER_7_151 ();
 sg13g2_decap_4 FILLER_7_158 ();
 sg13g2_fill_2 FILLER_7_162 ();
 sg13g2_fill_1 FILLER_7_191 ();
 sg13g2_decap_4 FILLER_7_196 ();
 sg13g2_fill_2 FILLER_7_200 ();
 sg13g2_fill_2 FILLER_7_273 ();
 sg13g2_fill_1 FILLER_7_275 ();
 sg13g2_fill_1 FILLER_7_310 ();
 sg13g2_fill_2 FILLER_7_319 ();
 sg13g2_fill_1 FILLER_7_321 ();
 sg13g2_decap_8 FILLER_7_358 ();
 sg13g2_fill_2 FILLER_7_365 ();
 sg13g2_fill_1 FILLER_7_390 ();
 sg13g2_fill_1 FILLER_7_397 ();
 sg13g2_fill_2 FILLER_7_419 ();
 sg13g2_fill_1 FILLER_7_421 ();
 sg13g2_fill_2 FILLER_7_426 ();
 sg13g2_fill_2 FILLER_7_475 ();
 sg13g2_fill_2 FILLER_7_504 ();
 sg13g2_fill_2 FILLER_7_519 ();
 sg13g2_decap_4 FILLER_7_571 ();
 sg13g2_fill_2 FILLER_7_615 ();
 sg13g2_fill_1 FILLER_7_644 ();
 sg13g2_decap_8 FILLER_7_649 ();
 sg13g2_fill_2 FILLER_7_665 ();
 sg13g2_fill_1 FILLER_7_667 ();
 sg13g2_fill_2 FILLER_7_704 ();
 sg13g2_fill_1 FILLER_7_706 ();
 sg13g2_decap_4 FILLER_7_718 ();
 sg13g2_fill_2 FILLER_7_722 ();
 sg13g2_fill_1 FILLER_7_748 ();
 sg13g2_decap_4 FILLER_7_757 ();
 sg13g2_fill_2 FILLER_7_761 ();
 sg13g2_fill_1 FILLER_7_772 ();
 sg13g2_fill_1 FILLER_7_810 ();
 sg13g2_decap_4 FILLER_7_852 ();
 sg13g2_fill_1 FILLER_7_856 ();
 sg13g2_fill_1 FILLER_7_923 ();
 sg13g2_decap_4 FILLER_7_956 ();
 sg13g2_fill_2 FILLER_7_1009 ();
 sg13g2_fill_2 FILLER_7_1044 ();
 sg13g2_fill_1 FILLER_7_1078 ();
 sg13g2_decap_8 FILLER_7_1151 ();
 sg13g2_decap_8 FILLER_7_1158 ();
 sg13g2_decap_4 FILLER_7_1165 ();
 sg13g2_fill_2 FILLER_7_1169 ();
 sg13g2_fill_2 FILLER_7_1184 ();
 sg13g2_decap_4 FILLER_7_1217 ();
 sg13g2_fill_1 FILLER_7_1221 ();
 sg13g2_fill_1 FILLER_7_1226 ();
 sg13g2_fill_1 FILLER_7_1254 ();
 sg13g2_fill_1 FILLER_7_1260 ();
 sg13g2_fill_1 FILLER_7_1296 ();
 sg13g2_decap_8 FILLER_7_1306 ();
 sg13g2_fill_2 FILLER_7_1313 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_fill_2 FILLER_8_7 ();
 sg13g2_fill_1 FILLER_8_48 ();
 sg13g2_fill_2 FILLER_8_55 ();
 sg13g2_fill_1 FILLER_8_97 ();
 sg13g2_decap_4 FILLER_8_164 ();
 sg13g2_fill_1 FILLER_8_168 ();
 sg13g2_decap_8 FILLER_8_200 ();
 sg13g2_fill_1 FILLER_8_207 ();
 sg13g2_decap_8 FILLER_8_212 ();
 sg13g2_decap_4 FILLER_8_223 ();
 sg13g2_fill_2 FILLER_8_307 ();
 sg13g2_fill_1 FILLER_8_318 ();
 sg13g2_decap_4 FILLER_8_405 ();
 sg13g2_fill_2 FILLER_8_409 ();
 sg13g2_fill_1 FILLER_8_425 ();
 sg13g2_fill_1 FILLER_8_446 ();
 sg13g2_fill_1 FILLER_8_469 ();
 sg13g2_fill_1 FILLER_8_524 ();
 sg13g2_fill_2 FILLER_8_530 ();
 sg13g2_fill_1 FILLER_8_532 ();
 sg13g2_fill_2 FILLER_8_584 ();
 sg13g2_fill_2 FILLER_8_595 ();
 sg13g2_fill_1 FILLER_8_660 ();
 sg13g2_decap_4 FILLER_8_697 ();
 sg13g2_fill_2 FILLER_8_701 ();
 sg13g2_fill_1 FILLER_8_713 ();
 sg13g2_fill_2 FILLER_8_741 ();
 sg13g2_fill_1 FILLER_8_743 ();
 sg13g2_decap_8 FILLER_8_771 ();
 sg13g2_fill_2 FILLER_8_778 ();
 sg13g2_fill_1 FILLER_8_790 ();
 sg13g2_decap_4 FILLER_8_795 ();
 sg13g2_decap_8 FILLER_8_808 ();
 sg13g2_decap_4 FILLER_8_815 ();
 sg13g2_fill_1 FILLER_8_819 ();
 sg13g2_decap_4 FILLER_8_825 ();
 sg13g2_fill_2 FILLER_8_852 ();
 sg13g2_fill_2 FILLER_8_863 ();
 sg13g2_fill_2 FILLER_8_874 ();
 sg13g2_fill_1 FILLER_8_898 ();
 sg13g2_decap_8 FILLER_8_955 ();
 sg13g2_decap_8 FILLER_8_962 ();
 sg13g2_fill_1 FILLER_8_974 ();
 sg13g2_fill_1 FILLER_8_980 ();
 sg13g2_decap_8 FILLER_8_1041 ();
 sg13g2_decap_4 FILLER_8_1048 ();
 sg13g2_fill_1 FILLER_8_1052 ();
 sg13g2_fill_2 FILLER_8_1070 ();
 sg13g2_fill_2 FILLER_8_1104 ();
 sg13g2_fill_1 FILLER_8_1112 ();
 sg13g2_fill_2 FILLER_8_1158 ();
 sg13g2_fill_2 FILLER_8_1173 ();
 sg13g2_fill_1 FILLER_8_1175 ();
 sg13g2_fill_2 FILLER_8_1216 ();
 sg13g2_fill_2 FILLER_8_1251 ();
 sg13g2_fill_1 FILLER_8_1253 ();
 sg13g2_fill_1 FILLER_8_1286 ();
 sg13g2_fill_1 FILLER_8_1314 ();
 sg13g2_decap_4 FILLER_9_0 ();
 sg13g2_fill_2 FILLER_9_4 ();
 sg13g2_fill_1 FILLER_9_82 ();
 sg13g2_fill_2 FILLER_9_124 ();
 sg13g2_fill_2 FILLER_9_149 ();
 sg13g2_fill_2 FILLER_9_156 ();
 sg13g2_fill_1 FILLER_9_158 ();
 sg13g2_fill_1 FILLER_9_168 ();
 sg13g2_decap_4 FILLER_9_316 ();
 sg13g2_fill_2 FILLER_9_320 ();
 sg13g2_fill_2 FILLER_9_335 ();
 sg13g2_decap_8 FILLER_9_361 ();
 sg13g2_fill_2 FILLER_9_368 ();
 sg13g2_fill_2 FILLER_9_383 ();
 sg13g2_fill_1 FILLER_9_402 ();
 sg13g2_fill_2 FILLER_9_416 ();
 sg13g2_fill_1 FILLER_9_418 ();
 sg13g2_fill_1 FILLER_9_463 ();
 sg13g2_fill_2 FILLER_9_481 ();
 sg13g2_fill_2 FILLER_9_582 ();
 sg13g2_fill_2 FILLER_9_598 ();
 sg13g2_fill_1 FILLER_9_606 ();
 sg13g2_decap_4 FILLER_9_634 ();
 sg13g2_fill_2 FILLER_9_665 ();
 sg13g2_fill_1 FILLER_9_667 ();
 sg13g2_fill_2 FILLER_9_705 ();
 sg13g2_fill_1 FILLER_9_707 ();
 sg13g2_fill_1 FILLER_9_739 ();
 sg13g2_decap_8 FILLER_9_772 ();
 sg13g2_fill_2 FILLER_9_779 ();
 sg13g2_fill_2 FILLER_9_813 ();
 sg13g2_decap_4 FILLER_9_820 ();
 sg13g2_decap_4 FILLER_9_856 ();
 sg13g2_fill_2 FILLER_9_919 ();
 sg13g2_fill_1 FILLER_9_946 ();
 sg13g2_fill_2 FILLER_9_983 ();
 sg13g2_decap_8 FILLER_9_990 ();
 sg13g2_decap_4 FILLER_9_997 ();
 sg13g2_fill_1 FILLER_9_1001 ();
 sg13g2_decap_4 FILLER_9_1015 ();
 sg13g2_fill_2 FILLER_9_1019 ();
 sg13g2_decap_8 FILLER_9_1047 ();
 sg13g2_fill_2 FILLER_9_1054 ();
 sg13g2_fill_1 FILLER_9_1056 ();
 sg13g2_fill_2 FILLER_9_1091 ();
 sg13g2_fill_1 FILLER_9_1093 ();
 sg13g2_fill_2 FILLER_9_1098 ();
 sg13g2_fill_1 FILLER_9_1100 ();
 sg13g2_fill_2 FILLER_9_1114 ();
 sg13g2_fill_1 FILLER_9_1116 ();
 sg13g2_decap_8 FILLER_9_1148 ();
 sg13g2_fill_1 FILLER_9_1155 ();
 sg13g2_fill_2 FILLER_9_1220 ();
 sg13g2_fill_1 FILLER_9_1222 ();
 sg13g2_fill_2 FILLER_9_1241 ();
 sg13g2_decap_8 FILLER_9_1304 ();
 sg13g2_decap_4 FILLER_9_1311 ();
 sg13g2_decap_4 FILLER_10_0 ();
 sg13g2_fill_1 FILLER_10_4 ();
 sg13g2_decap_8 FILLER_10_171 ();
 sg13g2_decap_4 FILLER_10_178 ();
 sg13g2_fill_1 FILLER_10_240 ();
 sg13g2_fill_2 FILLER_10_281 ();
 sg13g2_fill_1 FILLER_10_283 ();
 sg13g2_decap_8 FILLER_10_316 ();
 sg13g2_decap_8 FILLER_10_323 ();
 sg13g2_decap_4 FILLER_10_357 ();
 sg13g2_fill_1 FILLER_10_361 ();
 sg13g2_decap_4 FILLER_10_403 ();
 sg13g2_decap_4 FILLER_10_411 ();
 sg13g2_fill_1 FILLER_10_415 ();
 sg13g2_fill_2 FILLER_10_452 ();
 sg13g2_fill_1 FILLER_10_454 ();
 sg13g2_fill_1 FILLER_10_516 ();
 sg13g2_fill_2 FILLER_10_540 ();
 sg13g2_fill_1 FILLER_10_542 ();
 sg13g2_fill_1 FILLER_10_547 ();
 sg13g2_decap_8 FILLER_10_593 ();
 sg13g2_fill_1 FILLER_10_600 ();
 sg13g2_decap_8 FILLER_10_606 ();
 sg13g2_fill_2 FILLER_10_613 ();
 sg13g2_fill_1 FILLER_10_647 ();
 sg13g2_fill_2 FILLER_10_654 ();
 sg13g2_fill_2 FILLER_10_669 ();
 sg13g2_fill_2 FILLER_10_683 ();
 sg13g2_fill_1 FILLER_10_685 ();
 sg13g2_fill_1 FILLER_10_717 ();
 sg13g2_fill_1 FILLER_10_728 ();
 sg13g2_fill_1 FILLER_10_755 ();
 sg13g2_fill_1 FILLER_10_782 ();
 sg13g2_decap_8 FILLER_10_864 ();
 sg13g2_fill_1 FILLER_10_895 ();
 sg13g2_fill_2 FILLER_10_952 ();
 sg13g2_fill_1 FILLER_10_954 ();
 sg13g2_decap_4 FILLER_10_993 ();
 sg13g2_fill_1 FILLER_10_997 ();
 sg13g2_fill_2 FILLER_10_1030 ();
 sg13g2_fill_1 FILLER_10_1032 ();
 sg13g2_fill_1 FILLER_10_1044 ();
 sg13g2_fill_2 FILLER_10_1054 ();
 sg13g2_fill_1 FILLER_10_1056 ();
 sg13g2_fill_2 FILLER_10_1088 ();
 sg13g2_fill_2 FILLER_10_1103 ();
 sg13g2_fill_1 FILLER_10_1119 ();
 sg13g2_fill_2 FILLER_10_1125 ();
 sg13g2_fill_1 FILLER_10_1127 ();
 sg13g2_fill_2 FILLER_10_1134 ();
 sg13g2_fill_1 FILLER_10_1136 ();
 sg13g2_fill_2 FILLER_10_1150 ();
 sg13g2_fill_1 FILLER_10_1152 ();
 sg13g2_fill_2 FILLER_10_1180 ();
 sg13g2_fill_1 FILLER_10_1196 ();
 sg13g2_fill_2 FILLER_10_1231 ();
 sg13g2_fill_1 FILLER_10_1233 ();
 sg13g2_decap_8 FILLER_10_1300 ();
 sg13g2_decap_8 FILLER_10_1307 ();
 sg13g2_fill_1 FILLER_10_1314 ();
 sg13g2_fill_1 FILLER_11_0 ();
 sg13g2_fill_1 FILLER_11_36 ();
 sg13g2_fill_2 FILLER_11_74 ();
 sg13g2_fill_1 FILLER_11_76 ();
 sg13g2_fill_2 FILLER_11_90 ();
 sg13g2_fill_1 FILLER_11_92 ();
 sg13g2_decap_4 FILLER_11_157 ();
 sg13g2_decap_8 FILLER_11_170 ();
 sg13g2_decap_8 FILLER_11_177 ();
 sg13g2_decap_8 FILLER_11_184 ();
 sg13g2_fill_2 FILLER_11_270 ();
 sg13g2_fill_1 FILLER_11_272 ();
 sg13g2_decap_8 FILLER_11_277 ();
 sg13g2_fill_1 FILLER_11_284 ();
 sg13g2_decap_8 FILLER_11_319 ();
 sg13g2_fill_2 FILLER_11_363 ();
 sg13g2_fill_1 FILLER_11_365 ();
 sg13g2_fill_1 FILLER_11_412 ();
 sg13g2_fill_2 FILLER_11_417 ();
 sg13g2_fill_2 FILLER_11_427 ();
 sg13g2_fill_1 FILLER_11_429 ();
 sg13g2_decap_4 FILLER_11_434 ();
 sg13g2_fill_2 FILLER_11_438 ();
 sg13g2_fill_1 FILLER_11_453 ();
 sg13g2_fill_2 FILLER_11_495 ();
 sg13g2_fill_2 FILLER_11_506 ();
 sg13g2_fill_1 FILLER_11_508 ();
 sg13g2_fill_2 FILLER_11_513 ();
 sg13g2_fill_1 FILLER_11_515 ();
 sg13g2_fill_2 FILLER_11_535 ();
 sg13g2_fill_1 FILLER_11_537 ();
 sg13g2_decap_8 FILLER_11_547 ();
 sg13g2_decap_8 FILLER_11_615 ();
 sg13g2_decap_4 FILLER_11_622 ();
 sg13g2_fill_2 FILLER_11_626 ();
 sg13g2_fill_2 FILLER_11_651 ();
 sg13g2_fill_1 FILLER_11_653 ();
 sg13g2_decap_8 FILLER_11_663 ();
 sg13g2_decap_8 FILLER_11_670 ();
 sg13g2_decap_4 FILLER_11_677 ();
 sg13g2_fill_1 FILLER_11_681 ();
 sg13g2_decap_4 FILLER_11_703 ();
 sg13g2_fill_1 FILLER_11_707 ();
 sg13g2_fill_2 FILLER_11_720 ();
 sg13g2_decap_4 FILLER_11_765 ();
 sg13g2_fill_1 FILLER_11_769 ();
 sg13g2_decap_4 FILLER_11_774 ();
 sg13g2_fill_1 FILLER_11_778 ();
 sg13g2_decap_4 FILLER_11_783 ();
 sg13g2_fill_1 FILLER_11_824 ();
 sg13g2_fill_2 FILLER_11_846 ();
 sg13g2_fill_1 FILLER_11_848 ();
 sg13g2_fill_2 FILLER_11_871 ();
 sg13g2_fill_1 FILLER_11_873 ();
 sg13g2_fill_2 FILLER_11_903 ();
 sg13g2_fill_1 FILLER_11_905 ();
 sg13g2_fill_2 FILLER_11_932 ();
 sg13g2_fill_1 FILLER_11_934 ();
 sg13g2_fill_2 FILLER_11_940 ();
 sg13g2_fill_2 FILLER_11_948 ();
 sg13g2_fill_1 FILLER_11_950 ();
 sg13g2_fill_2 FILLER_11_960 ();
 sg13g2_decap_8 FILLER_11_989 ();
 sg13g2_fill_2 FILLER_11_996 ();
 sg13g2_fill_1 FILLER_11_1007 ();
 sg13g2_fill_1 FILLER_11_1054 ();
 sg13g2_fill_2 FILLER_11_1114 ();
 sg13g2_fill_1 FILLER_11_1116 ();
 sg13g2_fill_1 FILLER_11_1132 ();
 sg13g2_fill_1 FILLER_11_1146 ();
 sg13g2_fill_1 FILLER_11_1197 ();
 sg13g2_decap_8 FILLER_11_1240 ();
 sg13g2_decap_4 FILLER_11_1247 ();
 sg13g2_fill_1 FILLER_11_1251 ();
 sg13g2_fill_1 FILLER_11_1256 ();
 sg13g2_fill_2 FILLER_11_1275 ();
 sg13g2_fill_2 FILLER_11_1301 ();
 sg13g2_fill_1 FILLER_11_1303 ();
 sg13g2_fill_2 FILLER_11_1313 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_4 FILLER_12_50 ();
 sg13g2_fill_2 FILLER_12_54 ();
 sg13g2_fill_1 FILLER_12_174 ();
 sg13g2_fill_1 FILLER_12_179 ();
 sg13g2_decap_4 FILLER_12_194 ();
 sg13g2_fill_1 FILLER_12_198 ();
 sg13g2_fill_2 FILLER_12_226 ();
 sg13g2_fill_1 FILLER_12_228 ();
 sg13g2_decap_4 FILLER_12_261 ();
 sg13g2_decap_4 FILLER_12_270 ();
 sg13g2_decap_4 FILLER_12_278 ();
 sg13g2_decap_4 FILLER_12_292 ();
 sg13g2_fill_1 FILLER_12_296 ();
 sg13g2_decap_8 FILLER_12_301 ();
 sg13g2_decap_8 FILLER_12_308 ();
 sg13g2_fill_1 FILLER_12_315 ();
 sg13g2_fill_2 FILLER_12_326 ();
 sg13g2_fill_2 FILLER_12_341 ();
 sg13g2_decap_4 FILLER_12_361 ();
 sg13g2_fill_1 FILLER_12_420 ();
 sg13g2_fill_2 FILLER_12_438 ();
 sg13g2_fill_1 FILLER_12_440 ();
 sg13g2_fill_2 FILLER_12_454 ();
 sg13g2_fill_1 FILLER_12_456 ();
 sg13g2_decap_4 FILLER_12_484 ();
 sg13g2_fill_2 FILLER_12_488 ();
 sg13g2_decap_8 FILLER_12_504 ();
 sg13g2_fill_2 FILLER_12_511 ();
 sg13g2_fill_1 FILLER_12_513 ();
 sg13g2_fill_2 FILLER_12_573 ();
 sg13g2_decap_8 FILLER_12_620 ();
 sg13g2_decap_8 FILLER_12_663 ();
 sg13g2_decap_8 FILLER_12_691 ();
 sg13g2_fill_2 FILLER_12_698 ();
 sg13g2_fill_1 FILLER_12_700 ();
 sg13g2_fill_2 FILLER_12_706 ();
 sg13g2_fill_1 FILLER_12_708 ();
 sg13g2_decap_8 FILLER_12_742 ();
 sg13g2_decap_4 FILLER_12_749 ();
 sg13g2_decap_4 FILLER_12_801 ();
 sg13g2_decap_4 FILLER_12_814 ();
 sg13g2_decap_4 FILLER_12_823 ();
 sg13g2_fill_1 FILLER_12_827 ();
 sg13g2_fill_1 FILLER_12_926 ();
 sg13g2_fill_2 FILLER_12_979 ();
 sg13g2_decap_4 FILLER_12_990 ();
 sg13g2_fill_2 FILLER_12_1007 ();
 sg13g2_fill_1 FILLER_12_1009 ();
 sg13g2_fill_2 FILLER_12_1054 ();
 sg13g2_fill_1 FILLER_12_1056 ();
 sg13g2_fill_2 FILLER_12_1066 ();
 sg13g2_fill_2 FILLER_12_1167 ();
 sg13g2_fill_1 FILLER_12_1169 ();
 sg13g2_fill_1 FILLER_12_1184 ();
 sg13g2_fill_2 FILLER_12_1212 ();
 sg13g2_decap_8 FILLER_12_1247 ();
 sg13g2_decap_8 FILLER_12_1254 ();
 sg13g2_fill_2 FILLER_12_1261 ();
 sg13g2_fill_1 FILLER_12_1314 ();
 sg13g2_decap_4 FILLER_13_0 ();
 sg13g2_fill_1 FILLER_13_4 ();
 sg13g2_decap_8 FILLER_13_49 ();
 sg13g2_fill_2 FILLER_13_60 ();
 sg13g2_fill_1 FILLER_13_62 ();
 sg13g2_fill_1 FILLER_13_116 ();
 sg13g2_fill_2 FILLER_13_158 ();
 sg13g2_decap_4 FILLER_13_165 ();
 sg13g2_fill_1 FILLER_13_169 ();
 sg13g2_decap_4 FILLER_13_248 ();
 sg13g2_fill_2 FILLER_13_252 ();
 sg13g2_decap_8 FILLER_13_303 ();
 sg13g2_decap_8 FILLER_13_332 ();
 sg13g2_fill_1 FILLER_13_347 ();
 sg13g2_decap_4 FILLER_13_354 ();
 sg13g2_fill_1 FILLER_13_399 ();
 sg13g2_fill_2 FILLER_13_409 ();
 sg13g2_fill_2 FILLER_13_447 ();
 sg13g2_fill_2 FILLER_13_467 ();
 sg13g2_fill_1 FILLER_13_469 ();
 sg13g2_fill_1 FILLER_13_492 ();
 sg13g2_fill_2 FILLER_13_506 ();
 sg13g2_fill_2 FILLER_13_577 ();
 sg13g2_fill_2 FILLER_13_593 ();
 sg13g2_fill_1 FILLER_13_620 ();
 sg13g2_fill_1 FILLER_13_653 ();
 sg13g2_fill_2 FILLER_13_704 ();
 sg13g2_decap_4 FILLER_13_737 ();
 sg13g2_fill_2 FILLER_13_741 ();
 sg13g2_decap_8 FILLER_13_799 ();
 sg13g2_fill_1 FILLER_13_806 ();
 sg13g2_fill_2 FILLER_13_851 ();
 sg13g2_fill_2 FILLER_13_859 ();
 sg13g2_fill_1 FILLER_13_861 ();
 sg13g2_fill_2 FILLER_13_889 ();
 sg13g2_fill_1 FILLER_13_927 ();
 sg13g2_decap_8 FILLER_13_964 ();
 sg13g2_decap_8 FILLER_13_971 ();
 sg13g2_decap_8 FILLER_13_978 ();
 sg13g2_decap_4 FILLER_13_985 ();
 sg13g2_decap_4 FILLER_13_1026 ();
 sg13g2_fill_2 FILLER_13_1030 ();
 sg13g2_fill_2 FILLER_13_1063 ();
 sg13g2_fill_1 FILLER_13_1065 ();
 sg13g2_fill_2 FILLER_13_1071 ();
 sg13g2_fill_1 FILLER_13_1073 ();
 sg13g2_fill_1 FILLER_13_1102 ();
 sg13g2_fill_2 FILLER_13_1122 ();
 sg13g2_fill_2 FILLER_13_1137 ();
 sg13g2_fill_1 FILLER_13_1139 ();
 sg13g2_fill_2 FILLER_13_1162 ();
 sg13g2_fill_1 FILLER_13_1164 ();
 sg13g2_fill_1 FILLER_13_1210 ();
 sg13g2_decap_4 FILLER_13_1252 ();
 sg13g2_fill_2 FILLER_13_1256 ();
 sg13g2_fill_2 FILLER_13_1285 ();
 sg13g2_fill_1 FILLER_13_1314 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_fill_2 FILLER_14_49 ();
 sg13g2_fill_1 FILLER_14_106 ();
 sg13g2_fill_2 FILLER_14_168 ();
 sg13g2_fill_1 FILLER_14_170 ();
 sg13g2_fill_1 FILLER_14_204 ();
 sg13g2_fill_2 FILLER_14_210 ();
 sg13g2_fill_1 FILLER_14_212 ();
 sg13g2_fill_2 FILLER_14_222 ();
 sg13g2_fill_2 FILLER_14_246 ();
 sg13g2_fill_1 FILLER_14_248 ();
 sg13g2_fill_2 FILLER_14_341 ();
 sg13g2_fill_1 FILLER_14_343 ();
 sg13g2_fill_2 FILLER_14_395 ();
 sg13g2_fill_2 FILLER_14_403 ();
 sg13g2_fill_1 FILLER_14_405 ();
 sg13g2_fill_1 FILLER_14_444 ();
 sg13g2_fill_2 FILLER_14_449 ();
 sg13g2_fill_2 FILLER_14_511 ();
 sg13g2_fill_2 FILLER_14_539 ();
 sg13g2_fill_1 FILLER_14_541 ();
 sg13g2_decap_4 FILLER_14_569 ();
 sg13g2_fill_2 FILLER_14_573 ();
 sg13g2_decap_4 FILLER_14_579 ();
 sg13g2_fill_2 FILLER_14_583 ();
 sg13g2_fill_1 FILLER_14_616 ();
 sg13g2_decap_4 FILLER_14_621 ();
 sg13g2_fill_1 FILLER_14_625 ();
 sg13g2_fill_2 FILLER_14_635 ();
 sg13g2_fill_2 FILLER_14_717 ();
 sg13g2_fill_1 FILLER_14_719 ();
 sg13g2_fill_1 FILLER_14_740 ();
 sg13g2_fill_2 FILLER_14_809 ();
 sg13g2_fill_1 FILLER_14_811 ();
 sg13g2_fill_2 FILLER_14_853 ();
 sg13g2_fill_1 FILLER_14_855 ();
 sg13g2_fill_2 FILLER_14_880 ();
 sg13g2_fill_1 FILLER_14_882 ();
 sg13g2_fill_1 FILLER_14_892 ();
 sg13g2_fill_2 FILLER_14_902 ();
 sg13g2_fill_1 FILLER_14_904 ();
 sg13g2_decap_8 FILLER_14_914 ();
 sg13g2_decap_8 FILLER_14_921 ();
 sg13g2_decap_8 FILLER_14_928 ();
 sg13g2_fill_2 FILLER_14_935 ();
 sg13g2_decap_8 FILLER_14_1040 ();
 sg13g2_fill_2 FILLER_14_1047 ();
 sg13g2_decap_4 FILLER_14_1100 ();
 sg13g2_fill_1 FILLER_14_1104 ();
 sg13g2_fill_2 FILLER_14_1119 ();
 sg13g2_fill_1 FILLER_14_1121 ();
 sg13g2_decap_8 FILLER_14_1131 ();
 sg13g2_fill_2 FILLER_14_1203 ();
 sg13g2_fill_1 FILLER_14_1205 ();
 sg13g2_decap_4 FILLER_14_1258 ();
 sg13g2_fill_1 FILLER_14_1262 ();
 sg13g2_fill_2 FILLER_14_1303 ();
 sg13g2_fill_1 FILLER_14_1305 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_4 FILLER_15_7 ();
 sg13g2_fill_1 FILLER_15_11 ();
 sg13g2_fill_1 FILLER_15_16 ();
 sg13g2_decap_8 FILLER_15_45 ();
 sg13g2_fill_1 FILLER_15_52 ();
 sg13g2_fill_1 FILLER_15_111 ();
 sg13g2_fill_2 FILLER_15_174 ();
 sg13g2_fill_1 FILLER_15_176 ();
 sg13g2_fill_1 FILLER_15_203 ();
 sg13g2_fill_2 FILLER_15_221 ();
 sg13g2_fill_2 FILLER_15_268 ();
 sg13g2_fill_2 FILLER_15_349 ();
 sg13g2_fill_1 FILLER_15_351 ();
 sg13g2_fill_2 FILLER_15_394 ();
 sg13g2_fill_2 FILLER_15_423 ();
 sg13g2_fill_1 FILLER_15_425 ();
 sg13g2_fill_2 FILLER_15_435 ();
 sg13g2_fill_1 FILLER_15_437 ();
 sg13g2_decap_4 FILLER_15_477 ();
 sg13g2_fill_1 FILLER_15_481 ();
 sg13g2_fill_1 FILLER_15_514 ();
 sg13g2_fill_2 FILLER_15_555 ();
 sg13g2_decap_8 FILLER_15_572 ();
 sg13g2_decap_4 FILLER_15_612 ();
 sg13g2_fill_2 FILLER_15_616 ();
 sg13g2_decap_4 FILLER_15_637 ();
 sg13g2_fill_2 FILLER_15_641 ();
 sg13g2_decap_8 FILLER_15_648 ();
 sg13g2_decap_8 FILLER_15_655 ();
 sg13g2_fill_2 FILLER_15_662 ();
 sg13g2_decap_4 FILLER_15_741 ();
 sg13g2_fill_1 FILLER_15_745 ();
 sg13g2_fill_2 FILLER_15_751 ();
 sg13g2_fill_1 FILLER_15_753 ();
 sg13g2_fill_1 FILLER_15_771 ();
 sg13g2_fill_2 FILLER_15_804 ();
 sg13g2_fill_1 FILLER_15_806 ();
 sg13g2_decap_8 FILLER_15_869 ();
 sg13g2_fill_1 FILLER_15_876 ();
 sg13g2_decap_8 FILLER_15_881 ();
 sg13g2_decap_8 FILLER_15_888 ();
 sg13g2_decap_8 FILLER_15_895 ();
 sg13g2_decap_8 FILLER_15_910 ();
 sg13g2_decap_8 FILLER_15_917 ();
 sg13g2_fill_1 FILLER_15_924 ();
 sg13g2_fill_2 FILLER_15_929 ();
 sg13g2_fill_1 FILLER_15_945 ();
 sg13g2_fill_2 FILLER_15_952 ();
 sg13g2_fill_1 FILLER_15_954 ();
 sg13g2_fill_1 FILLER_15_1017 ();
 sg13g2_decap_8 FILLER_15_1027 ();
 sg13g2_decap_8 FILLER_15_1034 ();
 sg13g2_decap_8 FILLER_15_1041 ();
 sg13g2_decap_4 FILLER_15_1048 ();
 sg13g2_fill_2 FILLER_15_1052 ();
 sg13g2_decap_4 FILLER_15_1090 ();
 sg13g2_fill_1 FILLER_15_1094 ();
 sg13g2_decap_8 FILLER_15_1099 ();
 sg13g2_fill_2 FILLER_15_1106 ();
 sg13g2_fill_1 FILLER_15_1108 ();
 sg13g2_fill_2 FILLER_15_1141 ();
 sg13g2_decap_8 FILLER_15_1169 ();
 sg13g2_fill_2 FILLER_15_1217 ();
 sg13g2_decap_8 FILLER_15_1256 ();
 sg13g2_decap_8 FILLER_15_1263 ();
 sg13g2_fill_1 FILLER_15_1274 ();
 sg13g2_fill_1 FILLER_15_1293 ();
 sg13g2_decap_4 FILLER_15_1311 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_fill_1 FILLER_16_21 ();
 sg13g2_fill_2 FILLER_16_29 ();
 sg13g2_fill_1 FILLER_16_44 ();
 sg13g2_fill_1 FILLER_16_68 ();
 sg13g2_fill_1 FILLER_16_97 ();
 sg13g2_fill_2 FILLER_16_141 ();
 sg13g2_fill_1 FILLER_16_151 ();
 sg13g2_fill_1 FILLER_16_165 ();
 sg13g2_decap_8 FILLER_16_194 ();
 sg13g2_decap_4 FILLER_16_201 ();
 sg13g2_fill_2 FILLER_16_205 ();
 sg13g2_fill_2 FILLER_16_261 ();
 sg13g2_fill_1 FILLER_16_263 ();
 sg13g2_decap_8 FILLER_16_323 ();
 sg13g2_decap_4 FILLER_16_330 ();
 sg13g2_fill_1 FILLER_16_334 ();
 sg13g2_fill_1 FILLER_16_371 ();
 sg13g2_fill_2 FILLER_16_408 ();
 sg13g2_fill_1 FILLER_16_410 ();
 sg13g2_fill_2 FILLER_16_429 ();
 sg13g2_fill_1 FILLER_16_431 ();
 sg13g2_fill_2 FILLER_16_469 ();
 sg13g2_decap_8 FILLER_16_484 ();
 sg13g2_decap_8 FILLER_16_491 ();
 sg13g2_decap_4 FILLER_16_498 ();
 sg13g2_fill_1 FILLER_16_502 ();
 sg13g2_fill_2 FILLER_16_512 ();
 sg13g2_fill_2 FILLER_16_518 ();
 sg13g2_decap_8 FILLER_16_533 ();
 sg13g2_fill_2 FILLER_16_540 ();
 sg13g2_fill_2 FILLER_16_546 ();
 sg13g2_decap_4 FILLER_16_561 ();
 sg13g2_fill_1 FILLER_16_565 ();
 sg13g2_fill_2 FILLER_16_580 ();
 sg13g2_fill_2 FILLER_16_614 ();
 sg13g2_fill_1 FILLER_16_616 ();
 sg13g2_decap_8 FILLER_16_652 ();
 sg13g2_decap_8 FILLER_16_659 ();
 sg13g2_decap_4 FILLER_16_666 ();
 sg13g2_fill_1 FILLER_16_670 ();
 sg13g2_fill_2 FILLER_16_676 ();
 sg13g2_decap_8 FILLER_16_688 ();
 sg13g2_decap_8 FILLER_16_695 ();
 sg13g2_fill_2 FILLER_16_702 ();
 sg13g2_fill_1 FILLER_16_704 ();
 sg13g2_decap_8 FILLER_16_740 ();
 sg13g2_decap_8 FILLER_16_747 ();
 sg13g2_fill_1 FILLER_16_754 ();
 sg13g2_decap_4 FILLER_16_768 ();
 sg13g2_fill_1 FILLER_16_772 ();
 sg13g2_fill_1 FILLER_16_794 ();
 sg13g2_fill_2 FILLER_16_804 ();
 sg13g2_decap_4 FILLER_16_832 ();
 sg13g2_fill_1 FILLER_16_836 ();
 sg13g2_fill_1 FILLER_16_858 ();
 sg13g2_decap_8 FILLER_16_872 ();
 sg13g2_fill_1 FILLER_16_879 ();
 sg13g2_decap_4 FILLER_16_907 ();
 sg13g2_fill_2 FILLER_16_911 ();
 sg13g2_fill_2 FILLER_16_917 ();
 sg13g2_fill_1 FILLER_16_919 ();
 sg13g2_fill_1 FILLER_16_956 ();
 sg13g2_fill_2 FILLER_16_1001 ();
 sg13g2_fill_1 FILLER_16_1003 ();
 sg13g2_decap_8 FILLER_16_1017 ();
 sg13g2_fill_2 FILLER_16_1024 ();
 sg13g2_fill_1 FILLER_16_1026 ();
 sg13g2_decap_4 FILLER_16_1054 ();
 sg13g2_fill_2 FILLER_16_1084 ();
 sg13g2_fill_1 FILLER_16_1086 ();
 sg13g2_fill_1 FILLER_16_1150 ();
 sg13g2_decap_4 FILLER_16_1178 ();
 sg13g2_decap_8 FILLER_16_1257 ();
 sg13g2_decap_8 FILLER_16_1264 ();
 sg13g2_decap_8 FILLER_16_1302 ();
 sg13g2_decap_4 FILLER_16_1309 ();
 sg13g2_fill_2 FILLER_16_1313 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_fill_2 FILLER_17_14 ();
 sg13g2_fill_1 FILLER_17_16 ();
 sg13g2_fill_2 FILLER_17_27 ();
 sg13g2_decap_8 FILLER_17_38 ();
 sg13g2_fill_1 FILLER_17_45 ();
 sg13g2_decap_8 FILLER_17_68 ();
 sg13g2_fill_2 FILLER_17_75 ();
 sg13g2_fill_1 FILLER_17_87 ();
 sg13g2_fill_2 FILLER_17_93 ();
 sg13g2_fill_2 FILLER_17_123 ();
 sg13g2_decap_4 FILLER_17_166 ();
 sg13g2_fill_1 FILLER_17_170 ();
 sg13g2_decap_8 FILLER_17_179 ();
 sg13g2_fill_2 FILLER_17_186 ();
 sg13g2_fill_1 FILLER_17_188 ();
 sg13g2_fill_2 FILLER_17_216 ();
 sg13g2_fill_1 FILLER_17_218 ();
 sg13g2_decap_8 FILLER_17_266 ();
 sg13g2_decap_8 FILLER_17_322 ();
 sg13g2_fill_2 FILLER_17_329 ();
 sg13g2_fill_2 FILLER_17_372 ();
 sg13g2_fill_1 FILLER_17_374 ();
 sg13g2_fill_1 FILLER_17_388 ();
 sg13g2_fill_2 FILLER_17_412 ();
 sg13g2_fill_1 FILLER_17_414 ();
 sg13g2_fill_2 FILLER_17_474 ();
 sg13g2_decap_8 FILLER_17_481 ();
 sg13g2_fill_2 FILLER_17_488 ();
 sg13g2_fill_1 FILLER_17_490 ();
 sg13g2_fill_2 FILLER_17_597 ();
 sg13g2_fill_1 FILLER_17_599 ();
 sg13g2_fill_2 FILLER_17_659 ();
 sg13g2_fill_1 FILLER_17_665 ();
 sg13g2_fill_2 FILLER_17_670 ();
 sg13g2_fill_1 FILLER_17_672 ();
 sg13g2_decap_4 FILLER_17_683 ();
 sg13g2_fill_1 FILLER_17_687 ();
 sg13g2_decap_8 FILLER_17_697 ();
 sg13g2_decap_4 FILLER_17_740 ();
 sg13g2_decap_4 FILLER_17_771 ();
 sg13g2_fill_2 FILLER_17_775 ();
 sg13g2_fill_2 FILLER_17_799 ();
 sg13g2_fill_1 FILLER_17_801 ();
 sg13g2_decap_8 FILLER_17_820 ();
 sg13g2_decap_8 FILLER_17_827 ();
 sg13g2_fill_2 FILLER_17_834 ();
 sg13g2_fill_2 FILLER_17_927 ();
 sg13g2_fill_1 FILLER_17_929 ();
 sg13g2_fill_1 FILLER_17_971 ();
 sg13g2_fill_1 FILLER_17_976 ();
 sg13g2_fill_2 FILLER_17_981 ();
 sg13g2_fill_2 FILLER_17_991 ();
 sg13g2_decap_4 FILLER_17_1060 ();
 sg13g2_fill_2 FILLER_17_1064 ();
 sg13g2_fill_2 FILLER_17_1070 ();
 sg13g2_fill_1 FILLER_17_1076 ();
 sg13g2_fill_1 FILLER_17_1124 ();
 sg13g2_fill_2 FILLER_17_1145 ();
 sg13g2_fill_1 FILLER_17_1147 ();
 sg13g2_fill_1 FILLER_17_1190 ();
 sg13g2_fill_1 FILLER_17_1218 ();
 sg13g2_fill_2 FILLER_17_1232 ();
 sg13g2_fill_1 FILLER_17_1234 ();
 sg13g2_decap_8 FILLER_17_1243 ();
 sg13g2_decap_4 FILLER_17_1250 ();
 sg13g2_fill_2 FILLER_17_1254 ();
 sg13g2_decap_4 FILLER_17_1260 ();
 sg13g2_fill_1 FILLER_17_1314 ();
 sg13g2_decap_4 FILLER_18_0 ();
 sg13g2_fill_1 FILLER_18_4 ();
 sg13g2_fill_2 FILLER_18_41 ();
 sg13g2_fill_1 FILLER_18_43 ();
 sg13g2_decap_4 FILLER_18_71 ();
 sg13g2_fill_1 FILLER_18_115 ();
 sg13g2_fill_1 FILLER_18_126 ();
 sg13g2_fill_1 FILLER_18_154 ();
 sg13g2_fill_2 FILLER_18_165 ();
 sg13g2_fill_1 FILLER_18_167 ();
 sg13g2_decap_8 FILLER_18_172 ();
 sg13g2_decap_8 FILLER_18_179 ();
 sg13g2_decap_4 FILLER_18_186 ();
 sg13g2_fill_2 FILLER_18_190 ();
 sg13g2_decap_8 FILLER_18_260 ();
 sg13g2_decap_8 FILLER_18_267 ();
 sg13g2_fill_2 FILLER_18_274 ();
 sg13g2_decap_8 FILLER_18_324 ();
 sg13g2_fill_1 FILLER_18_331 ();
 sg13g2_fill_1 FILLER_18_358 ();
 sg13g2_decap_8 FILLER_18_368 ();
 sg13g2_decap_8 FILLER_18_375 ();
 sg13g2_fill_1 FILLER_18_382 ();
 sg13g2_fill_2 FILLER_18_441 ();
 sg13g2_decap_4 FILLER_18_534 ();
 sg13g2_fill_2 FILLER_18_587 ();
 sg13g2_fill_1 FILLER_18_589 ();
 sg13g2_decap_4 FILLER_18_697 ();
 sg13g2_fill_1 FILLER_18_701 ();
 sg13g2_fill_2 FILLER_18_732 ();
 sg13g2_fill_1 FILLER_18_774 ();
 sg13g2_fill_2 FILLER_18_811 ();
 sg13g2_fill_2 FILLER_18_849 ();
 sg13g2_fill_1 FILLER_18_851 ();
 sg13g2_fill_2 FILLER_18_879 ();
 sg13g2_fill_2 FILLER_18_944 ();
 sg13g2_fill_1 FILLER_18_951 ();
 sg13g2_fill_2 FILLER_18_969 ();
 sg13g2_fill_1 FILLER_18_971 ();
 sg13g2_fill_2 FILLER_18_1008 ();
 sg13g2_fill_2 FILLER_18_1045 ();
 sg13g2_fill_1 FILLER_18_1047 ();
 sg13g2_fill_1 FILLER_18_1075 ();
 sg13g2_fill_2 FILLER_18_1089 ();
 sg13g2_fill_1 FILLER_18_1091 ();
 sg13g2_fill_1 FILLER_18_1128 ();
 sg13g2_fill_2 FILLER_18_1138 ();
 sg13g2_fill_1 FILLER_18_1140 ();
 sg13g2_fill_2 FILLER_18_1154 ();
 sg13g2_fill_1 FILLER_18_1156 ();
 sg13g2_fill_1 FILLER_18_1170 ();
 sg13g2_fill_2 FILLER_18_1189 ();
 sg13g2_fill_1 FILLER_18_1191 ();
 sg13g2_fill_1 FILLER_18_1210 ();
 sg13g2_fill_1 FILLER_18_1215 ();
 sg13g2_fill_1 FILLER_18_1246 ();
 sg13g2_fill_1 FILLER_18_1314 ();
 sg13g2_fill_1 FILLER_19_0 ();
 sg13g2_fill_2 FILLER_19_53 ();
 sg13g2_fill_1 FILLER_19_111 ();
 sg13g2_fill_2 FILLER_19_127 ();
 sg13g2_fill_2 FILLER_19_138 ();
 sg13g2_fill_1 FILLER_19_140 ();
 sg13g2_decap_8 FILLER_19_191 ();
 sg13g2_fill_2 FILLER_19_198 ();
 sg13g2_fill_1 FILLER_19_200 ();
 sg13g2_fill_1 FILLER_19_232 ();
 sg13g2_decap_8 FILLER_19_268 ();
 sg13g2_decap_8 FILLER_19_275 ();
 sg13g2_fill_2 FILLER_19_282 ();
 sg13g2_fill_1 FILLER_19_326 ();
 sg13g2_fill_1 FILLER_19_371 ();
 sg13g2_fill_2 FILLER_19_399 ();
 sg13g2_fill_1 FILLER_19_401 ();
 sg13g2_fill_2 FILLER_19_457 ();
 sg13g2_fill_1 FILLER_19_459 ();
 sg13g2_fill_1 FILLER_19_497 ();
 sg13g2_fill_1 FILLER_19_539 ();
 sg13g2_decap_4 FILLER_19_609 ();
 sg13g2_fill_2 FILLER_19_618 ();
 sg13g2_fill_1 FILLER_19_620 ();
 sg13g2_fill_2 FILLER_19_729 ();
 sg13g2_fill_1 FILLER_19_743 ();
 sg13g2_fill_1 FILLER_19_757 ();
 sg13g2_fill_2 FILLER_19_794 ();
 sg13g2_fill_1 FILLER_19_850 ();
 sg13g2_decap_8 FILLER_19_873 ();
 sg13g2_fill_1 FILLER_19_880 ();
 sg13g2_fill_2 FILLER_19_894 ();
 sg13g2_fill_1 FILLER_19_937 ();
 sg13g2_fill_2 FILLER_19_948 ();
 sg13g2_fill_1 FILLER_19_950 ();
 sg13g2_decap_8 FILLER_19_982 ();
 sg13g2_decap_8 FILLER_19_989 ();
 sg13g2_decap_8 FILLER_19_996 ();
 sg13g2_decap_8 FILLER_19_1007 ();
 sg13g2_decap_4 FILLER_19_1014 ();
 sg13g2_fill_2 FILLER_19_1018 ();
 sg13g2_fill_1 FILLER_19_1033 ();
 sg13g2_fill_2 FILLER_19_1042 ();
 sg13g2_fill_2 FILLER_19_1048 ();
 sg13g2_fill_1 FILLER_19_1071 ();
 sg13g2_fill_2 FILLER_19_1085 ();
 sg13g2_decap_8 FILLER_19_1106 ();
 sg13g2_decap_8 FILLER_19_1113 ();
 sg13g2_fill_2 FILLER_19_1160 ();
 sg13g2_decap_8 FILLER_19_1166 ();
 sg13g2_fill_2 FILLER_19_1173 ();
 sg13g2_fill_1 FILLER_19_1175 ();
 sg13g2_decap_4 FILLER_19_1261 ();
 sg13g2_fill_1 FILLER_19_1265 ();
 sg13g2_fill_1 FILLER_19_1314 ();
 sg13g2_fill_2 FILLER_20_0 ();
 sg13g2_fill_1 FILLER_20_2 ();
 sg13g2_fill_2 FILLER_20_36 ();
 sg13g2_fill_1 FILLER_20_38 ();
 sg13g2_decap_8 FILLER_20_70 ();
 sg13g2_fill_2 FILLER_20_144 ();
 sg13g2_fill_1 FILLER_20_146 ();
 sg13g2_decap_8 FILLER_20_195 ();
 sg13g2_fill_2 FILLER_20_202 ();
 sg13g2_fill_1 FILLER_20_231 ();
 sg13g2_fill_2 FILLER_20_264 ();
 sg13g2_decap_4 FILLER_20_290 ();
 sg13g2_fill_1 FILLER_20_298 ();
 sg13g2_fill_2 FILLER_20_314 ();
 sg13g2_decap_4 FILLER_20_352 ();
 sg13g2_fill_2 FILLER_20_356 ();
 sg13g2_fill_1 FILLER_20_367 ();
 sg13g2_fill_2 FILLER_20_422 ();
 sg13g2_fill_1 FILLER_20_424 ();
 sg13g2_decap_8 FILLER_20_487 ();
 sg13g2_decap_8 FILLER_20_494 ();
 sg13g2_decap_8 FILLER_20_501 ();
 sg13g2_fill_2 FILLER_20_508 ();
 sg13g2_fill_1 FILLER_20_510 ();
 sg13g2_decap_8 FILLER_20_533 ();
 sg13g2_decap_8 FILLER_20_540 ();
 sg13g2_decap_8 FILLER_20_547 ();
 sg13g2_fill_1 FILLER_20_554 ();
 sg13g2_decap_4 FILLER_20_613 ();
 sg13g2_fill_2 FILLER_20_655 ();
 sg13g2_fill_1 FILLER_20_657 ();
 sg13g2_fill_2 FILLER_20_676 ();
 sg13g2_decap_4 FILLER_20_713 ();
 sg13g2_decap_8 FILLER_20_744 ();
 sg13g2_decap_4 FILLER_20_751 ();
 sg13g2_fill_2 FILLER_20_764 ();
 sg13g2_fill_1 FILLER_20_766 ();
 sg13g2_fill_2 FILLER_20_802 ();
 sg13g2_fill_2 FILLER_20_843 ();
 sg13g2_fill_1 FILLER_20_845 ();
 sg13g2_decap_8 FILLER_20_863 ();
 sg13g2_decap_8 FILLER_20_870 ();
 sg13g2_decap_8 FILLER_20_877 ();
 sg13g2_fill_2 FILLER_20_901 ();
 sg13g2_fill_1 FILLER_20_903 ();
 sg13g2_fill_2 FILLER_20_922 ();
 sg13g2_fill_1 FILLER_20_938 ();
 sg13g2_fill_2 FILLER_20_996 ();
 sg13g2_fill_1 FILLER_20_998 ();
 sg13g2_decap_8 FILLER_20_1003 ();
 sg13g2_fill_2 FILLER_20_1010 ();
 sg13g2_fill_1 FILLER_20_1012 ();
 sg13g2_fill_2 FILLER_20_1018 ();
 sg13g2_fill_1 FILLER_20_1020 ();
 sg13g2_fill_2 FILLER_20_1048 ();
 sg13g2_fill_1 FILLER_20_1050 ();
 sg13g2_decap_8 FILLER_20_1109 ();
 sg13g2_fill_1 FILLER_20_1129 ();
 sg13g2_fill_2 FILLER_20_1156 ();
 sg13g2_decap_8 FILLER_20_1266 ();
 sg13g2_fill_1 FILLER_20_1273 ();
 sg13g2_fill_1 FILLER_20_1278 ();
 sg13g2_fill_1 FILLER_20_1314 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_34 ();
 sg13g2_fill_1 FILLER_21_41 ();
 sg13g2_decap_4 FILLER_21_52 ();
 sg13g2_fill_2 FILLER_21_56 ();
 sg13g2_decap_8 FILLER_21_67 ();
 sg13g2_decap_4 FILLER_21_74 ();
 sg13g2_fill_2 FILLER_21_78 ();
 sg13g2_fill_1 FILLER_21_102 ();
 sg13g2_fill_2 FILLER_21_178 ();
 sg13g2_fill_1 FILLER_21_180 ();
 sg13g2_decap_8 FILLER_21_194 ();
 sg13g2_decap_8 FILLER_21_201 ();
 sg13g2_decap_4 FILLER_21_208 ();
 sg13g2_fill_1 FILLER_21_212 ();
 sg13g2_fill_1 FILLER_21_243 ();
 sg13g2_fill_2 FILLER_21_250 ();
 sg13g2_fill_1 FILLER_21_252 ();
 sg13g2_fill_1 FILLER_21_280 ();
 sg13g2_fill_2 FILLER_21_317 ();
 sg13g2_fill_1 FILLER_21_319 ();
 sg13g2_decap_8 FILLER_21_347 ();
 sg13g2_fill_2 FILLER_21_498 ();
 sg13g2_fill_1 FILLER_21_500 ();
 sg13g2_decap_8 FILLER_21_534 ();
 sg13g2_fill_2 FILLER_21_545 ();
 sg13g2_fill_1 FILLER_21_547 ();
 sg13g2_fill_2 FILLER_21_556 ();
 sg13g2_decap_4 FILLER_21_562 ();
 sg13g2_fill_1 FILLER_21_571 ();
 sg13g2_fill_1 FILLER_21_591 ();
 sg13g2_fill_2 FILLER_21_601 ();
 sg13g2_fill_1 FILLER_21_603 ();
 sg13g2_fill_1 FILLER_21_617 ();
 sg13g2_fill_1 FILLER_21_649 ();
 sg13g2_fill_1 FILLER_21_667 ();
 sg13g2_fill_2 FILLER_21_686 ();
 sg13g2_fill_2 FILLER_21_692 ();
 sg13g2_fill_1 FILLER_21_694 ();
 sg13g2_fill_1 FILLER_21_726 ();
 sg13g2_fill_2 FILLER_21_740 ();
 sg13g2_fill_1 FILLER_21_742 ();
 sg13g2_fill_1 FILLER_21_779 ();
 sg13g2_fill_2 FILLER_21_794 ();
 sg13g2_fill_1 FILLER_21_796 ();
 sg13g2_fill_2 FILLER_21_833 ();
 sg13g2_fill_2 FILLER_21_839 ();
 sg13g2_fill_1 FILLER_21_877 ();
 sg13g2_fill_2 FILLER_21_904 ();
 sg13g2_fill_1 FILLER_21_906 ();
 sg13g2_fill_2 FILLER_21_911 ();
 sg13g2_fill_1 FILLER_21_913 ();
 sg13g2_fill_1 FILLER_21_1032 ();
 sg13g2_decap_4 FILLER_21_1092 ();
 sg13g2_decap_8 FILLER_21_1140 ();
 sg13g2_decap_4 FILLER_21_1147 ();
 sg13g2_fill_2 FILLER_21_1151 ();
 sg13g2_fill_1 FILLER_21_1197 ();
 sg13g2_fill_2 FILLER_21_1211 ();
 sg13g2_fill_1 FILLER_21_1238 ();
 sg13g2_fill_1 FILLER_21_1261 ();
 sg13g2_fill_2 FILLER_21_1277 ();
 sg13g2_fill_2 FILLER_21_1312 ();
 sg13g2_fill_1 FILLER_21_1314 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_fill_1 FILLER_22_7 ();
 sg13g2_fill_1 FILLER_22_27 ();
 sg13g2_decap_4 FILLER_22_41 ();
 sg13g2_decap_4 FILLER_22_63 ();
 sg13g2_fill_1 FILLER_22_67 ();
 sg13g2_fill_1 FILLER_22_104 ();
 sg13g2_fill_1 FILLER_22_163 ();
 sg13g2_decap_8 FILLER_22_201 ();
 sg13g2_fill_2 FILLER_22_208 ();
 sg13g2_fill_1 FILLER_22_277 ();
 sg13g2_fill_2 FILLER_22_321 ();
 sg13g2_fill_2 FILLER_22_338 ();
 sg13g2_fill_1 FILLER_22_340 ();
 sg13g2_fill_2 FILLER_22_354 ();
 sg13g2_fill_2 FILLER_22_387 ();
 sg13g2_fill_2 FILLER_22_403 ();
 sg13g2_decap_8 FILLER_22_409 ();
 sg13g2_fill_1 FILLER_22_416 ();
 sg13g2_fill_2 FILLER_22_499 ();
 sg13g2_fill_1 FILLER_22_501 ();
 sg13g2_decap_8 FILLER_22_529 ();
 sg13g2_decap_4 FILLER_22_576 ();
 sg13g2_fill_1 FILLER_22_580 ();
 sg13g2_fill_2 FILLER_22_585 ();
 sg13g2_fill_1 FILLER_22_587 ();
 sg13g2_decap_4 FILLER_22_592 ();
 sg13g2_fill_2 FILLER_22_596 ();
 sg13g2_fill_2 FILLER_22_680 ();
 sg13g2_fill_2 FILLER_22_695 ();
 sg13g2_decap_4 FILLER_22_723 ();
 sg13g2_fill_1 FILLER_22_727 ();
 sg13g2_fill_2 FILLER_22_755 ();
 sg13g2_fill_2 FILLER_22_824 ();
 sg13g2_fill_2 FILLER_22_898 ();
 sg13g2_fill_1 FILLER_22_954 ();
 sg13g2_fill_1 FILLER_22_1009 ();
 sg13g2_fill_2 FILLER_22_1018 ();
 sg13g2_fill_2 FILLER_22_1044 ();
 sg13g2_fill_1 FILLER_22_1046 ();
 sg13g2_fill_1 FILLER_22_1137 ();
 sg13g2_decap_4 FILLER_22_1151 ();
 sg13g2_fill_1 FILLER_22_1155 ();
 sg13g2_decap_8 FILLER_22_1205 ();
 sg13g2_fill_2 FILLER_22_1212 ();
 sg13g2_fill_1 FILLER_22_1214 ();
 sg13g2_fill_1 FILLER_22_1314 ();
 sg13g2_decap_4 FILLER_23_0 ();
 sg13g2_decap_4 FILLER_23_58 ();
 sg13g2_fill_2 FILLER_23_62 ();
 sg13g2_fill_1 FILLER_23_142 ();
 sg13g2_decap_8 FILLER_23_197 ();
 sg13g2_decap_8 FILLER_23_204 ();
 sg13g2_fill_1 FILLER_23_260 ();
 sg13g2_fill_2 FILLER_23_274 ();
 sg13g2_fill_1 FILLER_23_276 ();
 sg13g2_fill_2 FILLER_23_286 ();
 sg13g2_decap_4 FILLER_23_292 ();
 sg13g2_decap_4 FILLER_23_300 ();
 sg13g2_fill_2 FILLER_23_313 ();
 sg13g2_fill_1 FILLER_23_320 ();
 sg13g2_decap_8 FILLER_23_365 ();
 sg13g2_fill_1 FILLER_23_372 ();
 sg13g2_fill_1 FILLER_23_399 ();
 sg13g2_fill_1 FILLER_23_404 ();
 sg13g2_fill_2 FILLER_23_431 ();
 sg13g2_fill_1 FILLER_23_433 ();
 sg13g2_fill_2 FILLER_23_459 ();
 sg13g2_fill_2 FILLER_23_506 ();
 sg13g2_fill_1 FILLER_23_508 ();
 sg13g2_fill_2 FILLER_23_568 ();
 sg13g2_fill_2 FILLER_23_588 ();
 sg13g2_decap_8 FILLER_23_677 ();
 sg13g2_fill_2 FILLER_23_684 ();
 sg13g2_fill_1 FILLER_23_686 ();
 sg13g2_fill_2 FILLER_23_696 ();
 sg13g2_fill_1 FILLER_23_711 ();
 sg13g2_fill_2 FILLER_23_792 ();
 sg13g2_fill_1 FILLER_23_794 ();
 sg13g2_fill_2 FILLER_23_818 ();
 sg13g2_fill_1 FILLER_23_820 ();
 sg13g2_fill_2 FILLER_23_835 ();
 sg13g2_fill_2 FILLER_23_886 ();
 sg13g2_fill_1 FILLER_23_888 ();
 sg13g2_decap_4 FILLER_23_953 ();
 sg13g2_fill_2 FILLER_23_974 ();
 sg13g2_fill_1 FILLER_23_976 ();
 sg13g2_fill_1 FILLER_23_1010 ();
 sg13g2_fill_2 FILLER_23_1046 ();
 sg13g2_decap_4 FILLER_23_1084 ();
 sg13g2_fill_1 FILLER_23_1088 ();
 sg13g2_fill_2 FILLER_23_1124 ();
 sg13g2_fill_2 FILLER_23_1164 ();
 sg13g2_fill_1 FILLER_23_1166 ();
 sg13g2_fill_2 FILLER_23_1173 ();
 sg13g2_decap_8 FILLER_23_1190 ();
 sg13g2_decap_8 FILLER_23_1197 ();
 sg13g2_decap_8 FILLER_23_1204 ();
 sg13g2_decap_8 FILLER_23_1211 ();
 sg13g2_fill_1 FILLER_23_1249 ();
 sg13g2_fill_1 FILLER_23_1314 ();
 sg13g2_fill_2 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_66 ();
 sg13g2_fill_2 FILLER_24_98 ();
 sg13g2_fill_1 FILLER_24_100 ();
 sg13g2_fill_2 FILLER_24_153 ();
 sg13g2_fill_1 FILLER_24_178 ();
 sg13g2_decap_8 FILLER_24_187 ();
 sg13g2_decap_8 FILLER_24_194 ();
 sg13g2_fill_2 FILLER_24_201 ();
 sg13g2_fill_2 FILLER_24_212 ();
 sg13g2_fill_1 FILLER_24_239 ();
 sg13g2_fill_2 FILLER_24_253 ();
 sg13g2_decap_4 FILLER_24_270 ();
 sg13g2_decap_4 FILLER_24_278 ();
 sg13g2_fill_2 FILLER_24_282 ();
 sg13g2_decap_8 FILLER_24_288 ();
 sg13g2_decap_8 FILLER_24_295 ();
 sg13g2_decap_8 FILLER_24_302 ();
 sg13g2_decap_8 FILLER_24_309 ();
 sg13g2_fill_2 FILLER_24_316 ();
 sg13g2_decap_8 FILLER_24_368 ();
 sg13g2_fill_2 FILLER_24_375 ();
 sg13g2_fill_2 FILLER_24_404 ();
 sg13g2_fill_1 FILLER_24_419 ();
 sg13g2_fill_2 FILLER_24_424 ();
 sg13g2_fill_1 FILLER_24_426 ();
 sg13g2_fill_1 FILLER_24_449 ();
 sg13g2_fill_1 FILLER_24_464 ();
 sg13g2_fill_2 FILLER_24_469 ();
 sg13g2_decap_4 FILLER_24_489 ();
 sg13g2_fill_2 FILLER_24_493 ();
 sg13g2_fill_1 FILLER_24_575 ();
 sg13g2_fill_1 FILLER_24_602 ();
 sg13g2_fill_2 FILLER_24_639 ();
 sg13g2_fill_1 FILLER_24_641 ();
 sg13g2_fill_1 FILLER_24_662 ();
 sg13g2_fill_2 FILLER_24_667 ();
 sg13g2_fill_1 FILLER_24_669 ();
 sg13g2_fill_2 FILLER_24_679 ();
 sg13g2_fill_2 FILLER_24_712 ();
 sg13g2_fill_2 FILLER_24_741 ();
 sg13g2_fill_1 FILLER_24_771 ();
 sg13g2_fill_2 FILLER_24_795 ();
 sg13g2_fill_1 FILLER_24_797 ();
 sg13g2_fill_2 FILLER_24_825 ();
 sg13g2_fill_2 FILLER_24_859 ();
 sg13g2_fill_1 FILLER_24_861 ();
 sg13g2_fill_2 FILLER_24_867 ();
 sg13g2_fill_1 FILLER_24_869 ();
 sg13g2_fill_1 FILLER_24_875 ();
 sg13g2_decap_8 FILLER_24_971 ();
 sg13g2_decap_8 FILLER_24_978 ();
 sg13g2_fill_1 FILLER_24_985 ();
 sg13g2_decap_8 FILLER_24_1003 ();
 sg13g2_fill_2 FILLER_24_1097 ();
 sg13g2_fill_1 FILLER_24_1099 ();
 sg13g2_fill_2 FILLER_24_1109 ();
 sg13g2_fill_2 FILLER_24_1149 ();
 sg13g2_fill_1 FILLER_24_1151 ();
 sg13g2_fill_2 FILLER_24_1158 ();
 sg13g2_fill_1 FILLER_24_1160 ();
 sg13g2_fill_2 FILLER_24_1174 ();
 sg13g2_fill_1 FILLER_24_1176 ();
 sg13g2_decap_4 FILLER_24_1215 ();
 sg13g2_fill_2 FILLER_24_1219 ();
 sg13g2_fill_2 FILLER_24_1230 ();
 sg13g2_fill_1 FILLER_24_1232 ();
 sg13g2_fill_1 FILLER_24_1241 ();
 sg13g2_fill_1 FILLER_24_1251 ();
 sg13g2_fill_2 FILLER_24_1266 ();
 sg13g2_fill_1 FILLER_24_1268 ();
 sg13g2_fill_1 FILLER_24_1286 ();
 sg13g2_fill_1 FILLER_24_1291 ();
 sg13g2_fill_1 FILLER_24_1314 ();
 sg13g2_fill_2 FILLER_25_0 ();
 sg13g2_fill_1 FILLER_25_2 ();
 sg13g2_fill_2 FILLER_25_33 ();
 sg13g2_fill_1 FILLER_25_35 ();
 sg13g2_fill_1 FILLER_25_62 ();
 sg13g2_fill_1 FILLER_25_71 ();
 sg13g2_fill_2 FILLER_25_85 ();
 sg13g2_fill_1 FILLER_25_105 ();
 sg13g2_fill_2 FILLER_25_112 ();
 sg13g2_fill_2 FILLER_25_127 ();
 sg13g2_fill_2 FILLER_25_152 ();
 sg13g2_fill_2 FILLER_25_171 ();
 sg13g2_fill_1 FILLER_25_173 ();
 sg13g2_decap_4 FILLER_25_178 ();
 sg13g2_fill_1 FILLER_25_187 ();
 sg13g2_decap_4 FILLER_25_208 ();
 sg13g2_fill_2 FILLER_25_212 ();
 sg13g2_fill_2 FILLER_25_223 ();
 sg13g2_fill_1 FILLER_25_225 ();
 sg13g2_fill_2 FILLER_25_236 ();
 sg13g2_decap_8 FILLER_25_260 ();
 sg13g2_fill_2 FILLER_25_267 ();
 sg13g2_fill_1 FILLER_25_329 ();
 sg13g2_fill_2 FILLER_25_378 ();
 sg13g2_fill_1 FILLER_25_422 ();
 sg13g2_decap_8 FILLER_25_477 ();
 sg13g2_fill_2 FILLER_25_484 ();
 sg13g2_fill_1 FILLER_25_486 ();
 sg13g2_fill_2 FILLER_25_500 ();
 sg13g2_decap_8 FILLER_25_515 ();
 sg13g2_fill_2 FILLER_25_522 ();
 sg13g2_fill_2 FILLER_25_529 ();
 sg13g2_fill_2 FILLER_25_618 ();
 sg13g2_fill_1 FILLER_25_620 ();
 sg13g2_fill_2 FILLER_25_667 ();
 sg13g2_fill_1 FILLER_25_669 ();
 sg13g2_fill_2 FILLER_25_701 ();
 sg13g2_fill_1 FILLER_25_726 ();
 sg13g2_fill_1 FILLER_25_740 ();
 sg13g2_fill_2 FILLER_25_754 ();
 sg13g2_fill_1 FILLER_25_756 ();
 sg13g2_fill_2 FILLER_25_775 ();
 sg13g2_fill_1 FILLER_25_777 ();
 sg13g2_fill_2 FILLER_25_824 ();
 sg13g2_fill_1 FILLER_25_856 ();
 sg13g2_fill_2 FILLER_25_872 ();
 sg13g2_fill_2 FILLER_25_902 ();
 sg13g2_fill_1 FILLER_25_915 ();
 sg13g2_fill_1 FILLER_25_925 ();
 sg13g2_decap_8 FILLER_25_939 ();
 sg13g2_decap_8 FILLER_25_946 ();
 sg13g2_decap_4 FILLER_25_953 ();
 sg13g2_fill_1 FILLER_25_957 ();
 sg13g2_decap_8 FILLER_25_969 ();
 sg13g2_decap_8 FILLER_25_1007 ();
 sg13g2_fill_2 FILLER_25_1027 ();
 sg13g2_fill_1 FILLER_25_1039 ();
 sg13g2_fill_1 FILLER_25_1067 ();
 sg13g2_fill_2 FILLER_25_1121 ();
 sg13g2_fill_1 FILLER_25_1123 ();
 sg13g2_fill_2 FILLER_25_1138 ();
 sg13g2_fill_2 FILLER_25_1226 ();
 sg13g2_fill_1 FILLER_25_1228 ();
 sg13g2_fill_2 FILLER_25_1238 ();
 sg13g2_fill_1 FILLER_25_1240 ();
 sg13g2_fill_1 FILLER_25_1273 ();
 sg13g2_fill_2 FILLER_25_1278 ();
 sg13g2_fill_1 FILLER_25_1280 ();
 sg13g2_fill_1 FILLER_25_1314 ();
 sg13g2_fill_2 FILLER_26_0 ();
 sg13g2_fill_1 FILLER_26_37 ();
 sg13g2_fill_2 FILLER_26_65 ();
 sg13g2_decap_4 FILLER_26_72 ();
 sg13g2_fill_2 FILLER_26_81 ();
 sg13g2_fill_2 FILLER_26_118 ();
 sg13g2_fill_1 FILLER_26_142 ();
 sg13g2_fill_1 FILLER_26_154 ();
 sg13g2_decap_4 FILLER_26_183 ();
 sg13g2_decap_4 FILLER_26_250 ();
 sg13g2_fill_1 FILLER_26_254 ();
 sg13g2_fill_2 FILLER_26_282 ();
 sg13g2_fill_1 FILLER_26_284 ();
 sg13g2_fill_1 FILLER_26_359 ();
 sg13g2_fill_2 FILLER_26_369 ();
 sg13g2_fill_1 FILLER_26_371 ();
 sg13g2_fill_1 FILLER_26_425 ();
 sg13g2_fill_2 FILLER_26_515 ();
 sg13g2_fill_1 FILLER_26_517 ();
 sg13g2_fill_1 FILLER_26_545 ();
 sg13g2_fill_1 FILLER_26_625 ();
 sg13g2_fill_2 FILLER_26_630 ();
 sg13g2_decap_8 FILLER_26_645 ();
 sg13g2_fill_2 FILLER_26_652 ();
 sg13g2_fill_1 FILLER_26_654 ();
 sg13g2_decap_8 FILLER_26_659 ();
 sg13g2_fill_1 FILLER_26_666 ();
 sg13g2_fill_1 FILLER_26_699 ();
 sg13g2_fill_2 FILLER_26_740 ();
 sg13g2_fill_2 FILLER_26_776 ();
 sg13g2_decap_4 FILLER_26_856 ();
 sg13g2_fill_1 FILLER_26_860 ();
 sg13g2_fill_2 FILLER_26_910 ();
 sg13g2_fill_2 FILLER_26_939 ();
 sg13g2_fill_2 FILLER_26_945 ();
 sg13g2_fill_1 FILLER_26_947 ();
 sg13g2_fill_2 FILLER_26_1011 ();
 sg13g2_fill_1 FILLER_26_1040 ();
 sg13g2_fill_2 FILLER_26_1068 ();
 sg13g2_fill_1 FILLER_26_1070 ();
 sg13g2_decap_4 FILLER_26_1125 ();
 sg13g2_fill_2 FILLER_26_1129 ();
 sg13g2_fill_2 FILLER_26_1161 ();
 sg13g2_fill_1 FILLER_26_1163 ();
 sg13g2_fill_2 FILLER_26_1191 ();
 sg13g2_fill_2 FILLER_26_1242 ();
 sg13g2_fill_2 FILLER_26_1284 ();
 sg13g2_fill_1 FILLER_26_1286 ();
 sg13g2_fill_1 FILLER_26_1314 ();
 sg13g2_decap_4 FILLER_27_0 ();
 sg13g2_fill_1 FILLER_27_4 ();
 sg13g2_fill_2 FILLER_27_38 ();
 sg13g2_fill_2 FILLER_27_58 ();
 sg13g2_fill_2 FILLER_27_87 ();
 sg13g2_fill_1 FILLER_27_162 ();
 sg13g2_decap_8 FILLER_27_214 ();
 sg13g2_decap_8 FILLER_27_221 ();
 sg13g2_fill_2 FILLER_27_228 ();
 sg13g2_fill_2 FILLER_27_257 ();
 sg13g2_fill_1 FILLER_27_259 ();
 sg13g2_fill_2 FILLER_27_264 ();
 sg13g2_fill_2 FILLER_27_306 ();
 sg13g2_fill_1 FILLER_27_308 ();
 sg13g2_decap_4 FILLER_27_313 ();
 sg13g2_fill_2 FILLER_27_367 ();
 sg13g2_fill_1 FILLER_27_369 ();
 sg13g2_fill_1 FILLER_27_387 ();
 sg13g2_fill_2 FILLER_27_405 ();
 sg13g2_fill_1 FILLER_27_440 ();
 sg13g2_fill_1 FILLER_27_447 ();
 sg13g2_fill_1 FILLER_27_525 ();
 sg13g2_decap_4 FILLER_27_656 ();
 sg13g2_fill_2 FILLER_27_709 ();
 sg13g2_fill_1 FILLER_27_711 ();
 sg13g2_fill_2 FILLER_27_748 ();
 sg13g2_fill_1 FILLER_27_750 ();
 sg13g2_decap_4 FILLER_27_778 ();
 sg13g2_fill_2 FILLER_27_813 ();
 sg13g2_decap_8 FILLER_27_855 ();
 sg13g2_fill_2 FILLER_27_862 ();
 sg13g2_fill_2 FILLER_27_900 ();
 sg13g2_fill_1 FILLER_27_902 ();
 sg13g2_decap_4 FILLER_27_930 ();
 sg13g2_fill_2 FILLER_27_934 ();
 sg13g2_fill_2 FILLER_27_963 ();
 sg13g2_fill_1 FILLER_27_970 ();
 sg13g2_fill_2 FILLER_27_1017 ();
 sg13g2_fill_1 FILLER_27_1019 ();
 sg13g2_fill_2 FILLER_27_1043 ();
 sg13g2_fill_2 FILLER_27_1058 ();
 sg13g2_fill_1 FILLER_27_1060 ();
 sg13g2_decap_8 FILLER_27_1129 ();
 sg13g2_decap_4 FILLER_27_1136 ();
 sg13g2_fill_2 FILLER_27_1140 ();
 sg13g2_fill_2 FILLER_27_1173 ();
 sg13g2_fill_1 FILLER_27_1175 ();
 sg13g2_fill_2 FILLER_27_1187 ();
 sg13g2_fill_2 FILLER_27_1224 ();
 sg13g2_fill_2 FILLER_27_1298 ();
 sg13g2_decap_4 FILLER_27_1309 ();
 sg13g2_fill_2 FILLER_27_1313 ();
 sg13g2_fill_2 FILLER_28_0 ();
 sg13g2_fill_2 FILLER_28_98 ();
 sg13g2_fill_2 FILLER_28_141 ();
 sg13g2_fill_1 FILLER_28_143 ();
 sg13g2_fill_2 FILLER_28_177 ();
 sg13g2_fill_1 FILLER_28_179 ();
 sg13g2_decap_8 FILLER_28_221 ();
 sg13g2_decap_8 FILLER_28_228 ();
 sg13g2_decap_8 FILLER_28_266 ();
 sg13g2_decap_4 FILLER_28_273 ();
 sg13g2_fill_2 FILLER_28_324 ();
 sg13g2_decap_4 FILLER_28_330 ();
 sg13g2_fill_2 FILLER_28_334 ();
 sg13g2_decap_4 FILLER_28_372 ();
 sg13g2_fill_2 FILLER_28_376 ();
 sg13g2_fill_2 FILLER_28_409 ();
 sg13g2_fill_2 FILLER_28_485 ();
 sg13g2_fill_2 FILLER_28_496 ();
 sg13g2_fill_1 FILLER_28_540 ();
 sg13g2_decap_4 FILLER_28_622 ();
 sg13g2_fill_2 FILLER_28_671 ();
 sg13g2_fill_1 FILLER_28_673 ();
 sg13g2_fill_1 FILLER_28_688 ();
 sg13g2_fill_2 FILLER_28_742 ();
 sg13g2_decap_4 FILLER_28_771 ();
 sg13g2_fill_2 FILLER_28_789 ();
 sg13g2_fill_1 FILLER_28_791 ();
 sg13g2_fill_1 FILLER_28_823 ();
 sg13g2_decap_4 FILLER_28_855 ();
 sg13g2_fill_1 FILLER_28_881 ();
 sg13g2_fill_2 FILLER_28_896 ();
 sg13g2_fill_1 FILLER_28_961 ();
 sg13g2_fill_1 FILLER_28_994 ();
 sg13g2_fill_2 FILLER_28_1022 ();
 sg13g2_fill_1 FILLER_28_1024 ();
 sg13g2_fill_2 FILLER_28_1034 ();
 sg13g2_fill_2 FILLER_28_1058 ();
 sg13g2_fill_1 FILLER_28_1060 ();
 sg13g2_decap_8 FILLER_28_1139 ();
 sg13g2_decap_8 FILLER_28_1146 ();
 sg13g2_decap_4 FILLER_28_1153 ();
 sg13g2_fill_2 FILLER_28_1157 ();
 sg13g2_fill_2 FILLER_28_1163 ();
 sg13g2_fill_1 FILLER_28_1178 ();
 sg13g2_fill_1 FILLER_28_1205 ();
 sg13g2_fill_2 FILLER_28_1250 ();
 sg13g2_fill_1 FILLER_28_1252 ();
 sg13g2_fill_1 FILLER_28_1284 ();
 sg13g2_fill_2 FILLER_28_1294 ();
 sg13g2_decap_8 FILLER_28_1300 ();
 sg13g2_decap_8 FILLER_28_1307 ();
 sg13g2_fill_1 FILLER_28_1314 ();
 sg13g2_fill_2 FILLER_29_0 ();
 sg13g2_fill_1 FILLER_29_2 ();
 sg13g2_fill_2 FILLER_29_39 ();
 sg13g2_fill_2 FILLER_29_46 ();
 sg13g2_fill_2 FILLER_29_92 ();
 sg13g2_fill_1 FILLER_29_94 ();
 sg13g2_fill_2 FILLER_29_108 ();
 sg13g2_fill_1 FILLER_29_110 ();
 sg13g2_fill_2 FILLER_29_159 ();
 sg13g2_fill_1 FILLER_29_161 ();
 sg13g2_decap_8 FILLER_29_230 ();
 sg13g2_decap_4 FILLER_29_237 ();
 sg13g2_fill_2 FILLER_29_241 ();
 sg13g2_fill_1 FILLER_29_252 ();
 sg13g2_fill_1 FILLER_29_281 ();
 sg13g2_decap_4 FILLER_29_322 ();
 sg13g2_decap_8 FILLER_29_332 ();
 sg13g2_fill_2 FILLER_29_339 ();
 sg13g2_fill_1 FILLER_29_341 ();
 sg13g2_fill_2 FILLER_29_423 ();
 sg13g2_fill_1 FILLER_29_425 ();
 sg13g2_fill_1 FILLER_29_471 ();
 sg13g2_fill_1 FILLER_29_476 ();
 sg13g2_decap_4 FILLER_29_498 ();
 sg13g2_fill_1 FILLER_29_502 ();
 sg13g2_fill_1 FILLER_29_584 ();
 sg13g2_decap_8 FILLER_29_612 ();
 sg13g2_decap_8 FILLER_29_619 ();
 sg13g2_fill_2 FILLER_29_626 ();
 sg13g2_fill_1 FILLER_29_660 ();
 sg13g2_fill_2 FILLER_29_714 ();
 sg13g2_fill_1 FILLER_29_716 ();
 sg13g2_fill_2 FILLER_29_726 ();
 sg13g2_fill_2 FILLER_29_780 ();
 sg13g2_fill_2 FILLER_29_801 ();
 sg13g2_fill_1 FILLER_29_803 ();
 sg13g2_fill_2 FILLER_29_823 ();
 sg13g2_fill_1 FILLER_29_825 ();
 sg13g2_decap_4 FILLER_29_844 ();
 sg13g2_fill_1 FILLER_29_848 ();
 sg13g2_fill_1 FILLER_29_858 ();
 sg13g2_fill_2 FILLER_29_863 ();
 sg13g2_fill_1 FILLER_29_865 ();
 sg13g2_fill_1 FILLER_29_893 ();
 sg13g2_fill_1 FILLER_29_917 ();
 sg13g2_decap_4 FILLER_29_950 ();
 sg13g2_fill_1 FILLER_29_954 ();
 sg13g2_decap_4 FILLER_29_1136 ();
 sg13g2_fill_2 FILLER_29_1157 ();
 sg13g2_fill_1 FILLER_29_1159 ();
 sg13g2_fill_1 FILLER_29_1173 ();
 sg13g2_fill_2 FILLER_29_1211 ();
 sg13g2_fill_1 FILLER_29_1265 ();
 sg13g2_fill_1 FILLER_29_1271 ();
 sg13g2_decap_8 FILLER_29_1291 ();
 sg13g2_decap_8 FILLER_29_1298 ();
 sg13g2_decap_8 FILLER_29_1305 ();
 sg13g2_fill_2 FILLER_29_1312 ();
 sg13g2_fill_1 FILLER_29_1314 ();
 sg13g2_fill_2 FILLER_30_0 ();
 sg13g2_fill_1 FILLER_30_2 ();
 sg13g2_fill_1 FILLER_30_44 ();
 sg13g2_fill_1 FILLER_30_76 ();
 sg13g2_fill_1 FILLER_30_141 ();
 sg13g2_fill_2 FILLER_30_170 ();
 sg13g2_fill_1 FILLER_30_212 ();
 sg13g2_fill_2 FILLER_30_240 ();
 sg13g2_fill_1 FILLER_30_272 ();
 sg13g2_fill_1 FILLER_30_286 ();
 sg13g2_fill_2 FILLER_30_295 ();
 sg13g2_fill_1 FILLER_30_297 ();
 sg13g2_decap_4 FILLER_30_334 ();
 sg13g2_fill_2 FILLER_30_343 ();
 sg13g2_fill_1 FILLER_30_345 ();
 sg13g2_fill_2 FILLER_30_387 ();
 sg13g2_fill_2 FILLER_30_404 ();
 sg13g2_fill_2 FILLER_30_425 ();
 sg13g2_fill_2 FILLER_30_490 ();
 sg13g2_fill_1 FILLER_30_492 ();
 sg13g2_fill_2 FILLER_30_497 ();
 sg13g2_fill_1 FILLER_30_499 ();
 sg13g2_decap_4 FILLER_30_504 ();
 sg13g2_fill_1 FILLER_30_518 ();
 sg13g2_fill_1 FILLER_30_542 ();
 sg13g2_fill_1 FILLER_30_551 ();
 sg13g2_fill_1 FILLER_30_581 ();
 sg13g2_fill_2 FILLER_30_609 ();
 sg13g2_fill_1 FILLER_30_611 ();
 sg13g2_decap_4 FILLER_30_616 ();
 sg13g2_fill_2 FILLER_30_620 ();
 sg13g2_decap_8 FILLER_30_656 ();
 sg13g2_decap_8 FILLER_30_663 ();
 sg13g2_decap_4 FILLER_30_670 ();
 sg13g2_fill_1 FILLER_30_674 ();
 sg13g2_decap_4 FILLER_30_679 ();
 sg13g2_fill_1 FILLER_30_683 ();
 sg13g2_fill_2 FILLER_30_692 ();
 sg13g2_fill_2 FILLER_30_726 ();
 sg13g2_fill_1 FILLER_30_728 ();
 sg13g2_fill_2 FILLER_30_751 ();
 sg13g2_fill_1 FILLER_30_753 ();
 sg13g2_fill_2 FILLER_30_775 ();
 sg13g2_fill_1 FILLER_30_777 ();
 sg13g2_decap_4 FILLER_30_822 ();
 sg13g2_fill_1 FILLER_30_839 ();
 sg13g2_fill_1 FILLER_30_883 ();
 sg13g2_fill_1 FILLER_30_926 ();
 sg13g2_decap_8 FILLER_30_944 ();
 sg13g2_fill_1 FILLER_30_983 ();
 sg13g2_decap_4 FILLER_30_997 ();
 sg13g2_fill_2 FILLER_30_1001 ();
 sg13g2_fill_2 FILLER_30_1035 ();
 sg13g2_fill_1 FILLER_30_1081 ();
 sg13g2_fill_2 FILLER_30_1119 ();
 sg13g2_fill_2 FILLER_30_1135 ();
 sg13g2_fill_1 FILLER_30_1137 ();
 sg13g2_decap_8 FILLER_30_1214 ();
 sg13g2_fill_2 FILLER_30_1240 ();
 sg13g2_fill_1 FILLER_30_1242 ();
 sg13g2_decap_4 FILLER_30_1256 ();
 sg13g2_fill_1 FILLER_30_1260 ();
 sg13g2_fill_2 FILLER_30_1278 ();
 sg13g2_fill_1 FILLER_30_1280 ();
 sg13g2_decap_8 FILLER_30_1308 ();
 sg13g2_decap_4 FILLER_31_0 ();
 sg13g2_fill_1 FILLER_31_4 ();
 sg13g2_fill_2 FILLER_31_16 ();
 sg13g2_fill_2 FILLER_31_51 ();
 sg13g2_fill_1 FILLER_31_53 ();
 sg13g2_fill_2 FILLER_31_69 ();
 sg13g2_fill_2 FILLER_31_86 ();
 sg13g2_decap_8 FILLER_31_158 ();
 sg13g2_fill_1 FILLER_31_195 ();
 sg13g2_fill_1 FILLER_31_202 ();
 sg13g2_fill_1 FILLER_31_223 ();
 sg13g2_decap_8 FILLER_31_277 ();
 sg13g2_fill_2 FILLER_31_284 ();
 sg13g2_fill_1 FILLER_31_286 ();
 sg13g2_fill_1 FILLER_31_360 ();
 sg13g2_fill_2 FILLER_31_370 ();
 sg13g2_fill_1 FILLER_31_372 ();
 sg13g2_fill_2 FILLER_31_386 ();
 sg13g2_fill_1 FILLER_31_388 ();
 sg13g2_fill_1 FILLER_31_394 ();
 sg13g2_fill_2 FILLER_31_437 ();
 sg13g2_fill_1 FILLER_31_439 ();
 sg13g2_fill_2 FILLER_31_446 ();
 sg13g2_fill_2 FILLER_31_501 ();
 sg13g2_fill_1 FILLER_31_503 ();
 sg13g2_decap_8 FILLER_31_573 ();
 sg13g2_fill_2 FILLER_31_580 ();
 sg13g2_fill_2 FILLER_31_608 ();
 sg13g2_fill_1 FILLER_31_610 ();
 sg13g2_fill_2 FILLER_31_630 ();
 sg13g2_fill_1 FILLER_31_632 ();
 sg13g2_decap_8 FILLER_31_666 ();
 sg13g2_decap_8 FILLER_31_673 ();
 sg13g2_decap_8 FILLER_31_680 ();
 sg13g2_fill_2 FILLER_31_687 ();
 sg13g2_fill_2 FILLER_31_725 ();
 sg13g2_fill_2 FILLER_31_831 ();
 sg13g2_fill_2 FILLER_31_843 ();
 sg13g2_fill_1 FILLER_31_872 ();
 sg13g2_fill_1 FILLER_31_913 ();
 sg13g2_fill_1 FILLER_31_940 ();
 sg13g2_decap_8 FILLER_31_945 ();
 sg13g2_decap_4 FILLER_31_952 ();
 sg13g2_fill_2 FILLER_31_960 ();
 sg13g2_fill_1 FILLER_31_970 ();
 sg13g2_decap_4 FILLER_31_997 ();
 sg13g2_fill_2 FILLER_31_1033 ();
 sg13g2_fill_1 FILLER_31_1035 ();
 sg13g2_fill_2 FILLER_31_1049 ();
 sg13g2_fill_1 FILLER_31_1051 ();
 sg13g2_fill_2 FILLER_31_1118 ();
 sg13g2_fill_1 FILLER_31_1120 ();
 sg13g2_fill_1 FILLER_31_1140 ();
 sg13g2_decap_4 FILLER_31_1147 ();
 sg13g2_fill_2 FILLER_31_1156 ();
 sg13g2_fill_1 FILLER_31_1158 ();
 sg13g2_fill_2 FILLER_31_1191 ();
 sg13g2_decap_4 FILLER_31_1208 ();
 sg13g2_fill_2 FILLER_31_1221 ();
 sg13g2_fill_1 FILLER_31_1223 ();
 sg13g2_decap_8 FILLER_31_1229 ();
 sg13g2_fill_2 FILLER_31_1236 ();
 sg13g2_fill_1 FILLER_31_1238 ();
 sg13g2_fill_2 FILLER_31_1279 ();
 sg13g2_fill_1 FILLER_31_1281 ();
 sg13g2_decap_4 FILLER_31_1309 ();
 sg13g2_fill_2 FILLER_31_1313 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_fill_2 FILLER_32_7 ();
 sg13g2_fill_1 FILLER_32_9 ();
 sg13g2_fill_2 FILLER_32_92 ();
 sg13g2_fill_1 FILLER_32_126 ();
 sg13g2_fill_1 FILLER_32_167 ();
 sg13g2_fill_1 FILLER_32_242 ();
 sg13g2_decap_8 FILLER_32_279 ();
 sg13g2_fill_1 FILLER_32_286 ();
 sg13g2_decap_4 FILLER_32_344 ();
 sg13g2_fill_1 FILLER_32_361 ();
 sg13g2_decap_4 FILLER_32_406 ();
 sg13g2_fill_1 FILLER_32_454 ();
 sg13g2_fill_2 FILLER_32_463 ();
 sg13g2_fill_1 FILLER_32_465 ();
 sg13g2_decap_8 FILLER_32_562 ();
 sg13g2_fill_2 FILLER_32_569 ();
 sg13g2_fill_1 FILLER_32_571 ();
 sg13g2_fill_2 FILLER_32_633 ();
 sg13g2_fill_1 FILLER_32_635 ();
 sg13g2_fill_2 FILLER_32_647 ();
 sg13g2_fill_1 FILLER_32_649 ();
 sg13g2_fill_2 FILLER_32_656 ();
 sg13g2_decap_4 FILLER_32_685 ();
 sg13g2_fill_2 FILLER_32_747 ();
 sg13g2_fill_1 FILLER_32_779 ();
 sg13g2_fill_2 FILLER_32_789 ();
 sg13g2_fill_1 FILLER_32_822 ();
 sg13g2_fill_2 FILLER_32_859 ();
 sg13g2_fill_2 FILLER_32_902 ();
 sg13g2_fill_2 FILLER_32_944 ();
 sg13g2_fill_2 FILLER_32_959 ();
 sg13g2_fill_1 FILLER_32_961 ();
 sg13g2_fill_2 FILLER_32_1019 ();
 sg13g2_fill_2 FILLER_32_1030 ();
 sg13g2_fill_2 FILLER_32_1041 ();
 sg13g2_fill_1 FILLER_32_1043 ();
 sg13g2_decap_4 FILLER_32_1077 ();
 sg13g2_fill_1 FILLER_32_1090 ();
 sg13g2_decap_8 FILLER_32_1136 ();
 sg13g2_decap_8 FILLER_32_1143 ();
 sg13g2_fill_1 FILLER_32_1150 ();
 sg13g2_fill_1 FILLER_32_1166 ();
 sg13g2_decap_4 FILLER_32_1171 ();
 sg13g2_fill_2 FILLER_32_1175 ();
 sg13g2_decap_8 FILLER_32_1198 ();
 sg13g2_fill_2 FILLER_32_1245 ();
 sg13g2_fill_1 FILLER_32_1247 ();
 sg13g2_fill_1 FILLER_32_1296 ();
 sg13g2_decap_8 FILLER_32_1306 ();
 sg13g2_fill_2 FILLER_32_1313 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_4 FILLER_33_7 ();
 sg13g2_fill_2 FILLER_33_11 ();
 sg13g2_fill_2 FILLER_33_93 ();
 sg13g2_fill_1 FILLER_33_95 ();
 sg13g2_fill_2 FILLER_33_132 ();
 sg13g2_fill_1 FILLER_33_238 ();
 sg13g2_decap_4 FILLER_33_249 ();
 sg13g2_fill_1 FILLER_33_318 ();
 sg13g2_decap_8 FILLER_33_346 ();
 sg13g2_decap_8 FILLER_33_407 ();
 sg13g2_decap_4 FILLER_33_414 ();
 sg13g2_decap_4 FILLER_33_466 ();
 sg13g2_fill_1 FILLER_33_470 ();
 sg13g2_decap_4 FILLER_33_528 ();
 sg13g2_fill_1 FILLER_33_532 ();
 sg13g2_fill_1 FILLER_33_546 ();
 sg13g2_fill_1 FILLER_33_551 ();
 sg13g2_fill_2 FILLER_33_565 ();
 sg13g2_fill_1 FILLER_33_567 ();
 sg13g2_fill_1 FILLER_33_631 ();
 sg13g2_fill_1 FILLER_33_668 ();
 sg13g2_decap_8 FILLER_33_678 ();
 sg13g2_fill_2 FILLER_33_685 ();
 sg13g2_fill_1 FILLER_33_687 ();
 sg13g2_fill_2 FILLER_33_706 ();
 sg13g2_fill_1 FILLER_33_708 ();
 sg13g2_fill_2 FILLER_33_724 ();
 sg13g2_fill_1 FILLER_33_731 ();
 sg13g2_fill_2 FILLER_33_785 ();
 sg13g2_fill_2 FILLER_33_800 ();
 sg13g2_fill_1 FILLER_33_802 ();
 sg13g2_decap_4 FILLER_33_872 ();
 sg13g2_fill_1 FILLER_33_876 ();
 sg13g2_fill_2 FILLER_33_971 ();
 sg13g2_fill_2 FILLER_33_1004 ();
 sg13g2_decap_8 FILLER_33_1019 ();
 sg13g2_decap_4 FILLER_33_1026 ();
 sg13g2_fill_1 FILLER_33_1030 ();
 sg13g2_decap_4 FILLER_33_1067 ();
 sg13g2_decap_8 FILLER_33_1080 ();
 sg13g2_decap_8 FILLER_33_1087 ();
 sg13g2_fill_1 FILLER_33_1098 ();
 sg13g2_decap_8 FILLER_33_1156 ();
 sg13g2_decap_8 FILLER_33_1163 ();
 sg13g2_decap_4 FILLER_33_1170 ();
 sg13g2_fill_1 FILLER_33_1174 ();
 sg13g2_fill_2 FILLER_33_1192 ();
 sg13g2_fill_1 FILLER_33_1194 ();
 sg13g2_fill_2 FILLER_33_1200 ();
 sg13g2_fill_1 FILLER_33_1202 ();
 sg13g2_fill_2 FILLER_33_1248 ();
 sg13g2_fill_1 FILLER_33_1250 ();
 sg13g2_decap_4 FILLER_33_1270 ();
 sg13g2_fill_2 FILLER_33_1274 ();
 sg13g2_decap_4 FILLER_33_1285 ();
 sg13g2_fill_2 FILLER_33_1289 ();
 sg13g2_decap_8 FILLER_33_1300 ();
 sg13g2_decap_8 FILLER_33_1307 ();
 sg13g2_fill_1 FILLER_33_1314 ();
 sg13g2_fill_2 FILLER_34_0 ();
 sg13g2_fill_1 FILLER_34_2 ();
 sg13g2_decap_4 FILLER_34_38 ();
 sg13g2_fill_2 FILLER_34_42 ();
 sg13g2_fill_1 FILLER_34_57 ();
 sg13g2_fill_1 FILLER_34_76 ();
 sg13g2_fill_2 FILLER_34_108 ();
 sg13g2_fill_1 FILLER_34_110 ();
 sg13g2_decap_4 FILLER_34_160 ();
 sg13g2_fill_1 FILLER_34_164 ();
 sg13g2_fill_1 FILLER_34_205 ();
 sg13g2_decap_4 FILLER_34_232 ();
 sg13g2_fill_2 FILLER_34_282 ();
 sg13g2_fill_1 FILLER_34_284 ();
 sg13g2_fill_1 FILLER_34_331 ();
 sg13g2_decap_8 FILLER_34_376 ();
 sg13g2_fill_2 FILLER_34_383 ();
 sg13g2_decap_4 FILLER_34_389 ();
 sg13g2_fill_2 FILLER_34_414 ();
 sg13g2_fill_1 FILLER_34_421 ();
 sg13g2_fill_2 FILLER_34_428 ();
 sg13g2_decap_8 FILLER_34_539 ();
 sg13g2_decap_8 FILLER_34_546 ();
 sg13g2_fill_1 FILLER_34_553 ();
 sg13g2_fill_2 FILLER_34_581 ();
 sg13g2_fill_1 FILLER_34_583 ();
 sg13g2_fill_2 FILLER_34_601 ();
 sg13g2_fill_1 FILLER_34_603 ();
 sg13g2_fill_2 FILLER_34_658 ();
 sg13g2_fill_1 FILLER_34_660 ();
 sg13g2_decap_8 FILLER_34_677 ();
 sg13g2_decap_4 FILLER_34_684 ();
 sg13g2_decap_8 FILLER_34_701 ();
 sg13g2_fill_2 FILLER_34_712 ();
 sg13g2_fill_1 FILLER_34_714 ();
 sg13g2_fill_2 FILLER_34_728 ();
 sg13g2_fill_1 FILLER_34_730 ();
 sg13g2_decap_4 FILLER_34_744 ();
 sg13g2_fill_1 FILLER_34_748 ();
 sg13g2_fill_2 FILLER_34_785 ();
 sg13g2_fill_2 FILLER_34_813 ();
 sg13g2_fill_1 FILLER_34_815 ();
 sg13g2_fill_2 FILLER_34_886 ();
 sg13g2_fill_1 FILLER_34_901 ();
 sg13g2_fill_2 FILLER_34_926 ();
 sg13g2_fill_2 FILLER_34_966 ();
 sg13g2_fill_1 FILLER_34_968 ();
 sg13g2_fill_2 FILLER_34_973 ();
 sg13g2_decap_8 FILLER_34_1019 ();
 sg13g2_decap_8 FILLER_34_1026 ();
 sg13g2_decap_8 FILLER_34_1078 ();
 sg13g2_decap_4 FILLER_34_1098 ();
 sg13g2_fill_1 FILLER_34_1102 ();
 sg13g2_fill_2 FILLER_34_1107 ();
 sg13g2_fill_2 FILLER_34_1132 ();
 sg13g2_fill_1 FILLER_34_1134 ();
 sg13g2_fill_1 FILLER_34_1195 ();
 sg13g2_fill_1 FILLER_34_1205 ();
 sg13g2_fill_2 FILLER_34_1232 ();
 sg13g2_fill_2 FILLER_34_1271 ();
 sg13g2_fill_1 FILLER_34_1273 ();
 sg13g2_decap_8 FILLER_34_1306 ();
 sg13g2_fill_2 FILLER_34_1313 ();
 sg13g2_fill_1 FILLER_35_0 ();
 sg13g2_fill_1 FILLER_35_49 ();
 sg13g2_fill_1 FILLER_35_55 ();
 sg13g2_decap_4 FILLER_35_74 ();
 sg13g2_fill_2 FILLER_35_82 ();
 sg13g2_fill_2 FILLER_35_126 ();
 sg13g2_decap_8 FILLER_35_161 ();
 sg13g2_decap_8 FILLER_35_168 ();
 sg13g2_decap_4 FILLER_35_181 ();
 sg13g2_fill_1 FILLER_35_185 ();
 sg13g2_fill_2 FILLER_35_198 ();
 sg13g2_fill_2 FILLER_35_226 ();
 sg13g2_fill_2 FILLER_35_305 ();
 sg13g2_fill_1 FILLER_35_307 ();
 sg13g2_decap_4 FILLER_35_313 ();
 sg13g2_fill_2 FILLER_35_317 ();
 sg13g2_fill_2 FILLER_35_336 ();
 sg13g2_fill_1 FILLER_35_338 ();
 sg13g2_fill_2 FILLER_35_348 ();
 sg13g2_fill_1 FILLER_35_350 ();
 sg13g2_fill_2 FILLER_35_364 ();
 sg13g2_fill_1 FILLER_35_366 ();
 sg13g2_fill_2 FILLER_35_398 ();
 sg13g2_fill_1 FILLER_35_400 ();
 sg13g2_fill_1 FILLER_35_426 ();
 sg13g2_decap_4 FILLER_35_495 ();
 sg13g2_fill_2 FILLER_35_530 ();
 sg13g2_fill_1 FILLER_35_532 ();
 sg13g2_fill_2 FILLER_35_546 ();
 sg13g2_decap_4 FILLER_35_554 ();
 sg13g2_fill_1 FILLER_35_558 ();
 sg13g2_fill_2 FILLER_35_601 ();
 sg13g2_fill_2 FILLER_35_617 ();
 sg13g2_fill_1 FILLER_35_619 ();
 sg13g2_fill_2 FILLER_35_633 ();
 sg13g2_fill_1 FILLER_35_635 ();
 sg13g2_decap_4 FILLER_35_674 ();
 sg13g2_decap_8 FILLER_35_732 ();
 sg13g2_fill_2 FILLER_35_739 ();
 sg13g2_fill_1 FILLER_35_746 ();
 sg13g2_decap_8 FILLER_35_809 ();
 sg13g2_decap_8 FILLER_35_816 ();
 sg13g2_fill_2 FILLER_35_823 ();
 sg13g2_fill_1 FILLER_35_825 ();
 sg13g2_fill_1 FILLER_35_895 ();
 sg13g2_fill_2 FILLER_35_922 ();
 sg13g2_decap_8 FILLER_35_978 ();
 sg13g2_fill_2 FILLER_35_985 ();
 sg13g2_fill_2 FILLER_35_991 ();
 sg13g2_fill_2 FILLER_35_1015 ();
 sg13g2_fill_1 FILLER_35_1017 ();
 sg13g2_fill_1 FILLER_35_1035 ();
 sg13g2_fill_2 FILLER_35_1050 ();
 sg13g2_fill_2 FILLER_35_1065 ();
 sg13g2_decap_8 FILLER_35_1107 ();
 sg13g2_decap_4 FILLER_35_1114 ();
 sg13g2_fill_2 FILLER_35_1172 ();
 sg13g2_fill_2 FILLER_35_1210 ();
 sg13g2_fill_1 FILLER_35_1212 ();
 sg13g2_fill_2 FILLER_35_1265 ();
 sg13g2_fill_1 FILLER_35_1267 ();
 sg13g2_fill_2 FILLER_35_1281 ();
 sg13g2_fill_1 FILLER_35_1283 ();
 sg13g2_decap_8 FILLER_35_1288 ();
 sg13g2_decap_8 FILLER_35_1295 ();
 sg13g2_decap_8 FILLER_35_1302 ();
 sg13g2_decap_4 FILLER_35_1309 ();
 sg13g2_fill_2 FILLER_35_1313 ();
 sg13g2_decap_4 FILLER_36_0 ();
 sg13g2_fill_2 FILLER_36_4 ();
 sg13g2_decap_4 FILLER_36_24 ();
 sg13g2_fill_1 FILLER_36_70 ();
 sg13g2_fill_2 FILLER_36_84 ();
 sg13g2_fill_1 FILLER_36_86 ();
 sg13g2_fill_1 FILLER_36_165 ();
 sg13g2_fill_2 FILLER_36_171 ();
 sg13g2_fill_1 FILLER_36_173 ();
 sg13g2_fill_2 FILLER_36_231 ();
 sg13g2_decap_4 FILLER_36_237 ();
 sg13g2_fill_1 FILLER_36_241 ();
 sg13g2_decap_8 FILLER_36_326 ();
 sg13g2_decap_4 FILLER_36_333 ();
 sg13g2_decap_8 FILLER_36_341 ();
 sg13g2_decap_8 FILLER_36_348 ();
 sg13g2_decap_8 FILLER_36_355 ();
 sg13g2_fill_2 FILLER_36_362 ();
 sg13g2_fill_2 FILLER_36_418 ();
 sg13g2_fill_1 FILLER_36_429 ();
 sg13g2_decap_8 FILLER_36_457 ();
 sg13g2_decap_8 FILLER_36_464 ();
 sg13g2_decap_8 FILLER_36_471 ();
 sg13g2_fill_2 FILLER_36_478 ();
 sg13g2_fill_2 FILLER_36_498 ();
 sg13g2_fill_1 FILLER_36_500 ();
 sg13g2_fill_1 FILLER_36_533 ();
 sg13g2_fill_1 FILLER_36_561 ();
 sg13g2_decap_8 FILLER_36_644 ();
 sg13g2_fill_2 FILLER_36_651 ();
 sg13g2_fill_1 FILLER_36_653 ();
 sg13g2_decap_4 FILLER_36_681 ();
 sg13g2_decap_8 FILLER_36_817 ();
 sg13g2_fill_2 FILLER_36_824 ();
 sg13g2_fill_1 FILLER_36_826 ();
 sg13g2_decap_4 FILLER_36_831 ();
 sg13g2_fill_2 FILLER_36_848 ();
 sg13g2_fill_1 FILLER_36_850 ();
 sg13g2_fill_2 FILLER_36_864 ();
 sg13g2_fill_2 FILLER_36_871 ();
 sg13g2_decap_4 FILLER_36_911 ();
 sg13g2_fill_1 FILLER_36_915 ();
 sg13g2_fill_2 FILLER_36_930 ();
 sg13g2_fill_1 FILLER_36_932 ();
 sg13g2_fill_1 FILLER_36_942 ();
 sg13g2_decap_4 FILLER_36_988 ();
 sg13g2_fill_2 FILLER_36_1033 ();
 sg13g2_fill_1 FILLER_36_1035 ();
 sg13g2_fill_1 FILLER_36_1101 ();
 sg13g2_fill_1 FILLER_36_1165 ();
 sg13g2_fill_2 FILLER_36_1215 ();
 sg13g2_fill_1 FILLER_36_1244 ();
 sg13g2_decap_8 FILLER_36_1281 ();
 sg13g2_decap_8 FILLER_36_1288 ();
 sg13g2_decap_8 FILLER_36_1295 ();
 sg13g2_decap_8 FILLER_36_1302 ();
 sg13g2_decap_4 FILLER_36_1309 ();
 sg13g2_fill_2 FILLER_36_1313 ();
 sg13g2_fill_2 FILLER_37_0 ();
 sg13g2_fill_1 FILLER_37_2 ();
 sg13g2_decap_8 FILLER_37_46 ();
 sg13g2_fill_1 FILLER_37_53 ();
 sg13g2_fill_1 FILLER_37_73 ();
 sg13g2_decap_4 FILLER_37_87 ();
 sg13g2_fill_2 FILLER_37_132 ();
 sg13g2_fill_1 FILLER_37_134 ();
 sg13g2_fill_1 FILLER_37_144 ();
 sg13g2_fill_1 FILLER_37_196 ();
 sg13g2_decap_8 FILLER_37_233 ();
 sg13g2_decap_8 FILLER_37_240 ();
 sg13g2_fill_2 FILLER_37_247 ();
 sg13g2_decap_4 FILLER_37_262 ();
 sg13g2_fill_1 FILLER_37_266 ();
 sg13g2_fill_1 FILLER_37_327 ();
 sg13g2_decap_8 FILLER_37_350 ();
 sg13g2_decap_8 FILLER_37_357 ();
 sg13g2_decap_4 FILLER_37_364 ();
 sg13g2_fill_1 FILLER_37_368 ();
 sg13g2_fill_1 FILLER_37_373 ();
 sg13g2_decap_8 FILLER_37_378 ();
 sg13g2_decap_4 FILLER_37_385 ();
 sg13g2_fill_1 FILLER_37_421 ();
 sg13g2_fill_2 FILLER_37_444 ();
 sg13g2_fill_1 FILLER_37_446 ();
 sg13g2_fill_1 FILLER_37_465 ();
 sg13g2_fill_2 FILLER_37_470 ();
 sg13g2_decap_4 FILLER_37_485 ();
 sg13g2_fill_2 FILLER_37_495 ();
 sg13g2_fill_1 FILLER_37_497 ();
 sg13g2_fill_2 FILLER_37_533 ();
 sg13g2_decap_4 FILLER_37_615 ();
 sg13g2_fill_2 FILLER_37_628 ();
 sg13g2_decap_8 FILLER_37_657 ();
 sg13g2_fill_2 FILLER_37_664 ();
 sg13g2_fill_2 FILLER_37_675 ();
 sg13g2_fill_1 FILLER_37_677 ();
 sg13g2_fill_2 FILLER_37_773 ();
 sg13g2_fill_2 FILLER_37_782 ();
 sg13g2_fill_1 FILLER_37_784 ();
 sg13g2_fill_1 FILLER_37_809 ();
 sg13g2_decap_8 FILLER_37_814 ();
 sg13g2_fill_1 FILLER_37_821 ();
 sg13g2_fill_2 FILLER_37_853 ();
 sg13g2_fill_2 FILLER_37_859 ();
 sg13g2_fill_1 FILLER_37_861 ();
 sg13g2_fill_2 FILLER_37_866 ();
 sg13g2_fill_2 FILLER_37_910 ();
 sg13g2_fill_1 FILLER_37_982 ();
 sg13g2_decap_4 FILLER_37_1000 ();
 sg13g2_fill_2 FILLER_37_1004 ();
 sg13g2_fill_2 FILLER_37_1067 ();
 sg13g2_fill_1 FILLER_37_1069 ();
 sg13g2_decap_4 FILLER_37_1079 ();
 sg13g2_fill_1 FILLER_37_1083 ();
 sg13g2_fill_2 FILLER_37_1128 ();
 sg13g2_decap_4 FILLER_37_1166 ();
 sg13g2_fill_1 FILLER_37_1170 ();
 sg13g2_decap_4 FILLER_37_1175 ();
 sg13g2_fill_1 FILLER_37_1179 ();
 sg13g2_fill_2 FILLER_37_1206 ();
 sg13g2_fill_2 FILLER_37_1229 ();
 sg13g2_fill_1 FILLER_37_1231 ();
 sg13g2_decap_8 FILLER_37_1264 ();
 sg13g2_decap_8 FILLER_37_1271 ();
 sg13g2_decap_8 FILLER_37_1278 ();
 sg13g2_decap_8 FILLER_37_1285 ();
 sg13g2_decap_8 FILLER_37_1292 ();
 sg13g2_decap_8 FILLER_37_1299 ();
 sg13g2_decap_8 FILLER_37_1306 ();
 sg13g2_fill_2 FILLER_37_1313 ();
 sg13g2_fill_2 FILLER_38_0 ();
 sg13g2_fill_1 FILLER_38_2 ();
 sg13g2_decap_8 FILLER_38_37 ();
 sg13g2_decap_8 FILLER_38_44 ();
 sg13g2_fill_1 FILLER_38_55 ();
 sg13g2_fill_1 FILLER_38_92 ();
 sg13g2_decap_4 FILLER_38_100 ();
 sg13g2_fill_2 FILLER_38_163 ();
 sg13g2_fill_1 FILLER_38_165 ();
 sg13g2_fill_2 FILLER_38_193 ();
 sg13g2_fill_1 FILLER_38_204 ();
 sg13g2_decap_4 FILLER_38_245 ();
 sg13g2_decap_8 FILLER_38_266 ();
 sg13g2_fill_1 FILLER_38_273 ();
 sg13g2_fill_1 FILLER_38_300 ();
 sg13g2_decap_4 FILLER_38_383 ();
 sg13g2_fill_2 FILLER_38_387 ();
 sg13g2_fill_2 FILLER_38_406 ();
 sg13g2_fill_2 FILLER_38_429 ();
 sg13g2_fill_2 FILLER_38_459 ();
 sg13g2_decap_8 FILLER_38_488 ();
 sg13g2_decap_8 FILLER_38_495 ();
 sg13g2_decap_4 FILLER_38_502 ();
 sg13g2_fill_1 FILLER_38_506 ();
 sg13g2_decap_8 FILLER_38_519 ();
 sg13g2_decap_4 FILLER_38_526 ();
 sg13g2_fill_2 FILLER_38_530 ();
 sg13g2_decap_8 FILLER_38_557 ();
 sg13g2_decap_8 FILLER_38_564 ();
 sg13g2_fill_2 FILLER_38_571 ();
 sg13g2_fill_1 FILLER_38_573 ();
 sg13g2_fill_1 FILLER_38_587 ();
 sg13g2_fill_2 FILLER_38_601 ();
 sg13g2_fill_1 FILLER_38_603 ();
 sg13g2_fill_2 FILLER_38_613 ();
 sg13g2_fill_1 FILLER_38_615 ();
 sg13g2_decap_8 FILLER_38_680 ();
 sg13g2_decap_8 FILLER_38_705 ();
 sg13g2_fill_2 FILLER_38_712 ();
 sg13g2_fill_2 FILLER_38_806 ();
 sg13g2_decap_8 FILLER_38_852 ();
 sg13g2_decap_4 FILLER_38_859 ();
 sg13g2_fill_2 FILLER_38_863 ();
 sg13g2_decap_8 FILLER_38_947 ();
 sg13g2_fill_2 FILLER_38_954 ();
 sg13g2_fill_2 FILLER_38_964 ();
 sg13g2_fill_1 FILLER_38_966 ();
 sg13g2_decap_8 FILLER_38_1008 ();
 sg13g2_decap_4 FILLER_38_1015 ();
 sg13g2_fill_2 FILLER_38_1051 ();
 sg13g2_fill_1 FILLER_38_1053 ();
 sg13g2_fill_2 FILLER_38_1073 ();
 sg13g2_fill_1 FILLER_38_1075 ();
 sg13g2_fill_2 FILLER_38_1095 ();
 sg13g2_fill_1 FILLER_38_1097 ();
 sg13g2_fill_2 FILLER_38_1116 ();
 sg13g2_fill_2 FILLER_38_1177 ();
 sg13g2_fill_1 FILLER_38_1205 ();
 sg13g2_fill_2 FILLER_38_1211 ();
 sg13g2_fill_1 FILLER_38_1213 ();
 sg13g2_fill_2 FILLER_38_1236 ();
 sg13g2_fill_1 FILLER_38_1238 ();
 sg13g2_decap_8 FILLER_38_1265 ();
 sg13g2_decap_8 FILLER_38_1272 ();
 sg13g2_decap_8 FILLER_38_1279 ();
 sg13g2_decap_8 FILLER_38_1286 ();
 sg13g2_decap_8 FILLER_38_1293 ();
 sg13g2_decap_8 FILLER_38_1300 ();
 sg13g2_decap_8 FILLER_38_1307 ();
 sg13g2_fill_1 FILLER_38_1314 ();
 sg13g2_fill_1 FILLER_39_0 ();
 sg13g2_fill_2 FILLER_39_42 ();
 sg13g2_fill_1 FILLER_39_44 ();
 sg13g2_fill_2 FILLER_39_72 ();
 sg13g2_fill_2 FILLER_39_97 ();
 sg13g2_fill_1 FILLER_39_99 ();
 sg13g2_fill_2 FILLER_39_217 ();
 sg13g2_fill_1 FILLER_39_219 ();
 sg13g2_fill_1 FILLER_39_254 ();
 sg13g2_decap_4 FILLER_39_279 ();
 sg13g2_fill_1 FILLER_39_283 ();
 sg13g2_fill_1 FILLER_39_337 ();
 sg13g2_fill_2 FILLER_39_401 ();
 sg13g2_fill_1 FILLER_39_403 ();
 sg13g2_fill_1 FILLER_39_452 ();
 sg13g2_fill_2 FILLER_39_464 ();
 sg13g2_fill_2 FILLER_39_479 ();
 sg13g2_fill_1 FILLER_39_481 ();
 sg13g2_fill_2 FILLER_39_509 ();
 sg13g2_decap_8 FILLER_39_515 ();
 sg13g2_fill_1 FILLER_39_522 ();
 sg13g2_decap_8 FILLER_39_532 ();
 sg13g2_fill_2 FILLER_39_539 ();
 sg13g2_fill_1 FILLER_39_541 ();
 sg13g2_decap_4 FILLER_39_546 ();
 sg13g2_decap_8 FILLER_39_554 ();
 sg13g2_fill_2 FILLER_39_561 ();
 sg13g2_fill_2 FILLER_39_589 ();
 sg13g2_decap_8 FILLER_39_604 ();
 sg13g2_decap_4 FILLER_39_611 ();
 sg13g2_fill_1 FILLER_39_615 ();
 sg13g2_fill_1 FILLER_39_633 ();
 sg13g2_fill_1 FILLER_39_709 ();
 sg13g2_decap_8 FILLER_39_714 ();
 sg13g2_fill_2 FILLER_39_721 ();
 sg13g2_fill_1 FILLER_39_723 ();
 sg13g2_fill_2 FILLER_39_770 ();
 sg13g2_fill_1 FILLER_39_797 ();
 sg13g2_decap_8 FILLER_39_868 ();
 sg13g2_fill_2 FILLER_39_875 ();
 sg13g2_fill_2 FILLER_39_885 ();
 sg13g2_fill_1 FILLER_39_887 ();
 sg13g2_fill_1 FILLER_39_932 ();
 sg13g2_decap_8 FILLER_39_946 ();
 sg13g2_decap_8 FILLER_39_953 ();
 sg13g2_fill_1 FILLER_39_960 ();
 sg13g2_decap_8 FILLER_39_997 ();
 sg13g2_decap_4 FILLER_39_1004 ();
 sg13g2_fill_1 FILLER_39_1008 ();
 sg13g2_decap_4 FILLER_39_1022 ();
 sg13g2_fill_2 FILLER_39_1026 ();
 sg13g2_fill_2 FILLER_39_1036 ();
 sg13g2_fill_1 FILLER_39_1038 ();
 sg13g2_fill_2 FILLER_39_1048 ();
 sg13g2_fill_2 FILLER_39_1122 ();
 sg13g2_fill_2 FILLER_39_1155 ();
 sg13g2_fill_1 FILLER_39_1157 ();
 sg13g2_decap_4 FILLER_39_1167 ();
 sg13g2_fill_2 FILLER_39_1198 ();
 sg13g2_decap_8 FILLER_39_1241 ();
 sg13g2_fill_2 FILLER_39_1248 ();
 sg13g2_decap_4 FILLER_39_1258 ();
 sg13g2_decap_8 FILLER_39_1271 ();
 sg13g2_decap_8 FILLER_39_1278 ();
 sg13g2_decap_8 FILLER_39_1285 ();
 sg13g2_decap_8 FILLER_39_1292 ();
 sg13g2_decap_8 FILLER_39_1299 ();
 sg13g2_decap_8 FILLER_39_1306 ();
 sg13g2_fill_2 FILLER_39_1313 ();
 sg13g2_decap_8 FILLER_40_0 ();
 sg13g2_fill_2 FILLER_40_7 ();
 sg13g2_fill_1 FILLER_40_9 ();
 sg13g2_decap_4 FILLER_40_14 ();
 sg13g2_fill_1 FILLER_40_18 ();
 sg13g2_fill_2 FILLER_40_41 ();
 sg13g2_fill_1 FILLER_40_47 ();
 sg13g2_fill_1 FILLER_40_74 ();
 sg13g2_fill_2 FILLER_40_88 ();
 sg13g2_fill_1 FILLER_40_90 ();
 sg13g2_fill_1 FILLER_40_95 ();
 sg13g2_fill_1 FILLER_40_136 ();
 sg13g2_decap_8 FILLER_40_150 ();
 sg13g2_fill_1 FILLER_40_196 ();
 sg13g2_fill_1 FILLER_40_214 ();
 sg13g2_fill_2 FILLER_40_247 ();
 sg13g2_fill_2 FILLER_40_258 ();
 sg13g2_decap_8 FILLER_40_269 ();
 sg13g2_decap_4 FILLER_40_276 ();
 sg13g2_fill_2 FILLER_40_280 ();
 sg13g2_decap_8 FILLER_40_286 ();
 sg13g2_fill_2 FILLER_40_293 ();
 sg13g2_fill_2 FILLER_40_351 ();
 sg13g2_fill_1 FILLER_40_380 ();
 sg13g2_fill_1 FILLER_40_408 ();
 sg13g2_fill_1 FILLER_40_445 ();
 sg13g2_fill_2 FILLER_40_478 ();
 sg13g2_fill_1 FILLER_40_480 ();
 sg13g2_fill_1 FILLER_40_499 ();
 sg13g2_fill_1 FILLER_40_532 ();
 sg13g2_fill_1 FILLER_40_540 ();
 sg13g2_fill_1 FILLER_40_707 ();
 sg13g2_decap_8 FILLER_40_725 ();
 sg13g2_fill_2 FILLER_40_740 ();
 sg13g2_fill_2 FILLER_40_774 ();
 sg13g2_fill_1 FILLER_40_776 ();
 sg13g2_fill_2 FILLER_40_807 ();
 sg13g2_decap_4 FILLER_40_848 ();
 sg13g2_fill_2 FILLER_40_883 ();
 sg13g2_decap_4 FILLER_40_889 ();
 sg13g2_fill_2 FILLER_40_893 ();
 sg13g2_decap_8 FILLER_40_908 ();
 sg13g2_decap_8 FILLER_40_928 ();
 sg13g2_decap_8 FILLER_40_935 ();
 sg13g2_decap_8 FILLER_40_942 ();
 sg13g2_decap_8 FILLER_40_949 ();
 sg13g2_decap_4 FILLER_40_956 ();
 sg13g2_fill_2 FILLER_40_960 ();
 sg13g2_decap_4 FILLER_40_970 ();
 sg13g2_decap_8 FILLER_40_991 ();
 sg13g2_decap_4 FILLER_40_998 ();
 sg13g2_fill_2 FILLER_40_1002 ();
 sg13g2_fill_2 FILLER_40_1017 ();
 sg13g2_fill_1 FILLER_40_1019 ();
 sg13g2_decap_8 FILLER_40_1029 ();
 sg13g2_decap_8 FILLER_40_1036 ();
 sg13g2_decap_8 FILLER_40_1043 ();
 sg13g2_decap_8 FILLER_40_1050 ();
 sg13g2_fill_1 FILLER_40_1111 ();
 sg13g2_fill_1 FILLER_40_1166 ();
 sg13g2_fill_2 FILLER_40_1194 ();
 sg13g2_fill_1 FILLER_40_1196 ();
 sg13g2_decap_8 FILLER_40_1232 ();
 sg13g2_fill_2 FILLER_40_1239 ();
 sg13g2_fill_1 FILLER_40_1241 ();
 sg13g2_decap_8 FILLER_40_1273 ();
 sg13g2_decap_8 FILLER_40_1280 ();
 sg13g2_decap_8 FILLER_40_1287 ();
 sg13g2_decap_8 FILLER_40_1294 ();
 sg13g2_decap_8 FILLER_40_1301 ();
 sg13g2_decap_8 FILLER_40_1308 ();
 sg13g2_decap_8 FILLER_41_0 ();
 sg13g2_decap_4 FILLER_41_7 ();
 sg13g2_fill_2 FILLER_41_21 ();
 sg13g2_fill_1 FILLER_41_23 ();
 sg13g2_decap_8 FILLER_41_28 ();
 sg13g2_fill_2 FILLER_41_35 ();
 sg13g2_fill_1 FILLER_41_37 ();
 sg13g2_fill_1 FILLER_41_85 ();
 sg13g2_decap_4 FILLER_41_127 ();
 sg13g2_fill_2 FILLER_41_141 ();
 sg13g2_fill_1 FILLER_41_143 ();
 sg13g2_decap_4 FILLER_41_148 ();
 sg13g2_fill_2 FILLER_41_152 ();
 sg13g2_decap_8 FILLER_41_161 ();
 sg13g2_fill_1 FILLER_41_203 ();
 sg13g2_fill_1 FILLER_41_240 ();
 sg13g2_decap_8 FILLER_41_269 ();
 sg13g2_fill_1 FILLER_41_276 ();
 sg13g2_fill_1 FILLER_41_357 ();
 sg13g2_decap_8 FILLER_41_381 ();
 sg13g2_fill_1 FILLER_41_430 ();
 sg13g2_fill_1 FILLER_41_457 ();
 sg13g2_fill_2 FILLER_41_498 ();
 sg13g2_fill_2 FILLER_41_564 ();
 sg13g2_fill_1 FILLER_41_566 ();
 sg13g2_fill_2 FILLER_41_633 ();
 sg13g2_fill_1 FILLER_41_635 ();
 sg13g2_fill_2 FILLER_41_653 ();
 sg13g2_fill_1 FILLER_41_655 ();
 sg13g2_fill_2 FILLER_41_669 ();
 sg13g2_fill_1 FILLER_41_684 ();
 sg13g2_decap_4 FILLER_41_740 ();
 sg13g2_fill_1 FILLER_41_744 ();
 sg13g2_fill_2 FILLER_41_773 ();
 sg13g2_fill_2 FILLER_41_806 ();
 sg13g2_fill_1 FILLER_41_808 ();
 sg13g2_fill_2 FILLER_41_854 ();
 sg13g2_decap_4 FILLER_41_892 ();
 sg13g2_fill_1 FILLER_41_896 ();
 sg13g2_decap_4 FILLER_41_937 ();
 sg13g2_decap_4 FILLER_41_1027 ();
 sg13g2_fill_1 FILLER_41_1058 ();
 sg13g2_fill_1 FILLER_41_1077 ();
 sg13g2_fill_1 FILLER_41_1088 ();
 sg13g2_fill_2 FILLER_41_1167 ();
 sg13g2_fill_1 FILLER_41_1182 ();
 sg13g2_decap_8 FILLER_41_1192 ();
 sg13g2_fill_2 FILLER_41_1199 ();
 sg13g2_decap_8 FILLER_41_1269 ();
 sg13g2_decap_8 FILLER_41_1276 ();
 sg13g2_decap_8 FILLER_41_1283 ();
 sg13g2_decap_8 FILLER_41_1290 ();
 sg13g2_decap_8 FILLER_41_1297 ();
 sg13g2_decap_8 FILLER_41_1304 ();
 sg13g2_decap_4 FILLER_41_1311 ();
 sg13g2_fill_2 FILLER_42_0 ();
 sg13g2_fill_1 FILLER_42_2 ();
 sg13g2_fill_1 FILLER_42_31 ();
 sg13g2_fill_1 FILLER_42_133 ();
 sg13g2_decap_8 FILLER_42_167 ();
 sg13g2_decap_8 FILLER_42_174 ();
 sg13g2_decap_4 FILLER_42_181 ();
 sg13g2_decap_4 FILLER_42_260 ();
 sg13g2_fill_1 FILLER_42_264 ();
 sg13g2_decap_8 FILLER_42_279 ();
 sg13g2_decap_8 FILLER_42_286 ();
 sg13g2_decap_8 FILLER_42_293 ();
 sg13g2_decap_4 FILLER_42_300 ();
 sg13g2_fill_1 FILLER_42_304 ();
 sg13g2_decap_8 FILLER_42_309 ();
 sg13g2_fill_2 FILLER_42_316 ();
 sg13g2_decap_4 FILLER_42_327 ();
 sg13g2_fill_2 FILLER_42_344 ();
 sg13g2_decap_8 FILLER_42_359 ();
 sg13g2_fill_2 FILLER_42_376 ();
 sg13g2_fill_1 FILLER_42_378 ();
 sg13g2_fill_1 FILLER_42_392 ();
 sg13g2_fill_1 FILLER_42_401 ();
 sg13g2_fill_2 FILLER_42_430 ();
 sg13g2_fill_2 FILLER_42_459 ();
 sg13g2_fill_1 FILLER_42_461 ();
 sg13g2_fill_2 FILLER_42_472 ();
 sg13g2_fill_1 FILLER_42_474 ();
 sg13g2_decap_4 FILLER_42_533 ();
 sg13g2_fill_1 FILLER_42_537 ();
 sg13g2_decap_4 FILLER_42_590 ();
 sg13g2_fill_1 FILLER_42_594 ();
 sg13g2_decap_8 FILLER_42_603 ();
 sg13g2_decap_4 FILLER_42_610 ();
 sg13g2_decap_4 FILLER_42_664 ();
 sg13g2_fill_2 FILLER_42_668 ();
 sg13g2_fill_2 FILLER_42_741 ();
 sg13g2_fill_1 FILLER_42_743 ();
 sg13g2_decap_8 FILLER_42_791 ();
 sg13g2_decap_8 FILLER_42_798 ();
 sg13g2_fill_1 FILLER_42_805 ();
 sg13g2_decap_4 FILLER_42_832 ();
 sg13g2_fill_2 FILLER_42_911 ();
 sg13g2_fill_1 FILLER_42_913 ();
 sg13g2_fill_2 FILLER_42_964 ();
 sg13g2_fill_1 FILLER_42_966 ();
 sg13g2_fill_2 FILLER_42_999 ();
 sg13g2_fill_1 FILLER_42_1033 ();
 sg13g2_decap_8 FILLER_42_1051 ();
 sg13g2_fill_2 FILLER_42_1066 ();
 sg13g2_fill_2 FILLER_42_1082 ();
 sg13g2_fill_1 FILLER_42_1084 ();
 sg13g2_fill_2 FILLER_42_1094 ();
 sg13g2_fill_2 FILLER_42_1150 ();
 sg13g2_fill_1 FILLER_42_1152 ();
 sg13g2_fill_2 FILLER_42_1168 ();
 sg13g2_fill_1 FILLER_42_1174 ();
 sg13g2_fill_2 FILLER_42_1180 ();
 sg13g2_decap_8 FILLER_42_1188 ();
 sg13g2_decap_8 FILLER_42_1195 ();
 sg13g2_fill_2 FILLER_42_1206 ();
 sg13g2_fill_1 FILLER_42_1208 ();
 sg13g2_decap_8 FILLER_42_1231 ();
 sg13g2_decap_4 FILLER_42_1238 ();
 sg13g2_fill_1 FILLER_42_1242 ();
 sg13g2_fill_2 FILLER_42_1254 ();
 sg13g2_fill_1 FILLER_42_1256 ();
 sg13g2_decap_8 FILLER_42_1274 ();
 sg13g2_decap_8 FILLER_42_1281 ();
 sg13g2_decap_8 FILLER_42_1288 ();
 sg13g2_decap_8 FILLER_42_1295 ();
 sg13g2_decap_8 FILLER_42_1302 ();
 sg13g2_decap_4 FILLER_42_1309 ();
 sg13g2_fill_2 FILLER_42_1313 ();
 sg13g2_decap_8 FILLER_43_0 ();
 sg13g2_fill_1 FILLER_43_7 ();
 sg13g2_decap_8 FILLER_43_12 ();
 sg13g2_decap_8 FILLER_43_19 ();
 sg13g2_fill_2 FILLER_43_26 ();
 sg13g2_fill_1 FILLER_43_33 ();
 sg13g2_fill_2 FILLER_43_39 ();
 sg13g2_fill_2 FILLER_43_54 ();
 sg13g2_fill_1 FILLER_43_71 ();
 sg13g2_fill_1 FILLER_43_100 ();
 sg13g2_fill_2 FILLER_43_115 ();
 sg13g2_fill_1 FILLER_43_117 ();
 sg13g2_fill_2 FILLER_43_149 ();
 sg13g2_decap_8 FILLER_43_179 ();
 sg13g2_fill_1 FILLER_43_198 ();
 sg13g2_fill_1 FILLER_43_262 ();
 sg13g2_fill_2 FILLER_43_291 ();
 sg13g2_fill_1 FILLER_43_293 ();
 sg13g2_decap_8 FILLER_43_298 ();
 sg13g2_decap_4 FILLER_43_305 ();
 sg13g2_fill_1 FILLER_43_309 ();
 sg13g2_decap_8 FILLER_43_316 ();
 sg13g2_decap_8 FILLER_43_323 ();
 sg13g2_fill_1 FILLER_43_330 ();
 sg13g2_decap_8 FILLER_43_340 ();
 sg13g2_decap_8 FILLER_43_347 ();
 sg13g2_fill_2 FILLER_43_376 ();
 sg13g2_fill_2 FILLER_43_392 ();
 sg13g2_decap_4 FILLER_43_409 ();
 sg13g2_fill_2 FILLER_43_413 ();
 sg13g2_fill_2 FILLER_43_492 ();
 sg13g2_fill_1 FILLER_43_494 ();
 sg13g2_fill_2 FILLER_43_518 ();
 sg13g2_fill_1 FILLER_43_520 ();
 sg13g2_decap_4 FILLER_43_552 ();
 sg13g2_fill_1 FILLER_43_556 ();
 sg13g2_fill_1 FILLER_43_566 ();
 sg13g2_decap_8 FILLER_43_580 ();
 sg13g2_fill_2 FILLER_43_587 ();
 sg13g2_fill_1 FILLER_43_589 ();
 sg13g2_fill_2 FILLER_43_598 ();
 sg13g2_fill_2 FILLER_43_609 ();
 sg13g2_fill_1 FILLER_43_611 ();
 sg13g2_fill_1 FILLER_43_685 ();
 sg13g2_fill_2 FILLER_43_724 ();
 sg13g2_decap_8 FILLER_43_739 ();
 sg13g2_fill_1 FILLER_43_746 ();
 sg13g2_fill_1 FILLER_43_786 ();
 sg13g2_decap_8 FILLER_43_800 ();
 sg13g2_fill_2 FILLER_43_807 ();
 sg13g2_fill_1 FILLER_43_818 ();
 sg13g2_decap_8 FILLER_43_823 ();
 sg13g2_decap_8 FILLER_43_830 ();
 sg13g2_decap_4 FILLER_43_837 ();
 sg13g2_fill_2 FILLER_43_872 ();
 sg13g2_fill_2 FILLER_43_884 ();
 sg13g2_fill_1 FILLER_43_886 ();
 sg13g2_decap_4 FILLER_43_896 ();
 sg13g2_fill_2 FILLER_43_900 ();
 sg13g2_decap_8 FILLER_43_906 ();
 sg13g2_decap_4 FILLER_43_932 ();
 sg13g2_fill_1 FILLER_43_962 ();
 sg13g2_fill_1 FILLER_43_987 ();
 sg13g2_decap_8 FILLER_43_1050 ();
 sg13g2_decap_4 FILLER_43_1057 ();
 sg13g2_fill_2 FILLER_43_1061 ();
 sg13g2_decap_4 FILLER_43_1109 ();
 sg13g2_fill_2 FILLER_43_1113 ();
 sg13g2_fill_2 FILLER_43_1125 ();
 sg13g2_fill_1 FILLER_43_1127 ();
 sg13g2_fill_1 FILLER_43_1137 ();
 sg13g2_decap_4 FILLER_43_1159 ();
 sg13g2_fill_1 FILLER_43_1163 ();
 sg13g2_decap_8 FILLER_43_1181 ();
 sg13g2_fill_1 FILLER_43_1188 ();
 sg13g2_decap_8 FILLER_43_1233 ();
 sg13g2_fill_1 FILLER_43_1240 ();
 sg13g2_fill_2 FILLER_43_1246 ();
 sg13g2_decap_8 FILLER_43_1280 ();
 sg13g2_decap_8 FILLER_43_1287 ();
 sg13g2_decap_8 FILLER_43_1294 ();
 sg13g2_decap_8 FILLER_43_1301 ();
 sg13g2_decap_8 FILLER_43_1308 ();
 sg13g2_decap_4 FILLER_44_0 ();
 sg13g2_fill_2 FILLER_44_44 ();
 sg13g2_fill_1 FILLER_44_46 ();
 sg13g2_fill_2 FILLER_44_72 ();
 sg13g2_fill_1 FILLER_44_74 ();
 sg13g2_fill_1 FILLER_44_97 ();
 sg13g2_fill_1 FILLER_44_107 ();
 sg13g2_fill_1 FILLER_44_155 ();
 sg13g2_fill_1 FILLER_44_160 ();
 sg13g2_decap_4 FILLER_44_165 ();
 sg13g2_fill_2 FILLER_44_195 ();
 sg13g2_fill_1 FILLER_44_197 ();
 sg13g2_fill_2 FILLER_44_220 ();
 sg13g2_decap_4 FILLER_44_258 ();
 sg13g2_fill_1 FILLER_44_262 ();
 sg13g2_fill_1 FILLER_44_276 ();
 sg13g2_decap_8 FILLER_44_322 ();
 sg13g2_decap_4 FILLER_44_329 ();
 sg13g2_fill_1 FILLER_44_333 ();
 sg13g2_fill_1 FILLER_44_338 ();
 sg13g2_fill_1 FILLER_44_344 ();
 sg13g2_fill_1 FILLER_44_349 ();
 sg13g2_decap_8 FILLER_44_409 ();
 sg13g2_decap_8 FILLER_44_416 ();
 sg13g2_decap_4 FILLER_44_423 ();
 sg13g2_fill_1 FILLER_44_427 ();
 sg13g2_fill_2 FILLER_44_454 ();
 sg13g2_fill_1 FILLER_44_456 ();
 sg13g2_decap_8 FILLER_44_487 ();
 sg13g2_decap_4 FILLER_44_525 ();
 sg13g2_fill_1 FILLER_44_546 ();
 sg13g2_fill_2 FILLER_44_606 ();
 sg13g2_fill_1 FILLER_44_608 ();
 sg13g2_fill_2 FILLER_44_622 ();
 sg13g2_fill_1 FILLER_44_624 ();
 sg13g2_fill_2 FILLER_44_634 ();
 sg13g2_fill_1 FILLER_44_645 ();
 sg13g2_decap_8 FILLER_44_659 ();
 sg13g2_fill_2 FILLER_44_666 ();
 sg13g2_decap_8 FILLER_44_681 ();
 sg13g2_decap_4 FILLER_44_688 ();
 sg13g2_fill_2 FILLER_44_696 ();
 sg13g2_fill_2 FILLER_44_711 ();
 sg13g2_fill_1 FILLER_44_713 ();
 sg13g2_fill_1 FILLER_44_731 ();
 sg13g2_decap_8 FILLER_44_764 ();
 sg13g2_fill_1 FILLER_44_886 ();
 sg13g2_decap_8 FILLER_44_923 ();
 sg13g2_decap_8 FILLER_44_930 ();
 sg13g2_decap_4 FILLER_44_937 ();
 sg13g2_fill_1 FILLER_44_941 ();
 sg13g2_fill_2 FILLER_44_951 ();
 sg13g2_fill_1 FILLER_44_953 ();
 sg13g2_fill_2 FILLER_44_960 ();
 sg13g2_decap_4 FILLER_44_996 ();
 sg13g2_fill_2 FILLER_44_1000 ();
 sg13g2_fill_2 FILLER_44_1014 ();
 sg13g2_fill_2 FILLER_44_1042 ();
 sg13g2_fill_1 FILLER_44_1044 ();
 sg13g2_decap_4 FILLER_44_1049 ();
 sg13g2_fill_2 FILLER_44_1053 ();
 sg13g2_fill_2 FILLER_44_1126 ();
 sg13g2_fill_1 FILLER_44_1128 ();
 sg13g2_decap_4 FILLER_44_1156 ();
 sg13g2_decap_8 FILLER_44_1225 ();
 sg13g2_fill_2 FILLER_44_1232 ();
 sg13g2_fill_1 FILLER_44_1234 ();
 sg13g2_decap_8 FILLER_44_1267 ();
 sg13g2_decap_8 FILLER_44_1274 ();
 sg13g2_decap_8 FILLER_44_1281 ();
 sg13g2_decap_8 FILLER_44_1288 ();
 sg13g2_decap_8 FILLER_44_1295 ();
 sg13g2_decap_8 FILLER_44_1302 ();
 sg13g2_decap_4 FILLER_44_1309 ();
 sg13g2_fill_2 FILLER_44_1313 ();
 sg13g2_decap_8 FILLER_45_0 ();
 sg13g2_fill_2 FILLER_45_7 ();
 sg13g2_fill_2 FILLER_45_13 ();
 sg13g2_fill_2 FILLER_45_56 ();
 sg13g2_fill_1 FILLER_45_58 ();
 sg13g2_fill_2 FILLER_45_100 ();
 sg13g2_fill_1 FILLER_45_102 ();
 sg13g2_fill_1 FILLER_45_131 ();
 sg13g2_decap_4 FILLER_45_187 ();
 sg13g2_fill_2 FILLER_45_205 ();
 sg13g2_fill_1 FILLER_45_207 ();
 sg13g2_fill_2 FILLER_45_265 ();
 sg13g2_fill_1 FILLER_45_267 ();
 sg13g2_fill_2 FILLER_45_272 ();
 sg13g2_fill_2 FILLER_45_323 ();
 sg13g2_decap_4 FILLER_45_401 ();
 sg13g2_fill_1 FILLER_45_426 ();
 sg13g2_fill_1 FILLER_45_436 ();
 sg13g2_fill_1 FILLER_45_441 ();
 sg13g2_decap_8 FILLER_45_447 ();
 sg13g2_decap_4 FILLER_45_458 ();
 sg13g2_decap_8 FILLER_45_471 ();
 sg13g2_decap_8 FILLER_45_478 ();
 sg13g2_decap_4 FILLER_45_485 ();
 sg13g2_decap_8 FILLER_45_506 ();
 sg13g2_fill_2 FILLER_45_513 ();
 sg13g2_fill_1 FILLER_45_515 ();
 sg13g2_fill_1 FILLER_45_529 ();
 sg13g2_fill_1 FILLER_45_645 ();
 sg13g2_decap_8 FILLER_45_673 ();
 sg13g2_fill_1 FILLER_45_680 ();
 sg13g2_fill_1 FILLER_45_698 ();
 sg13g2_decap_4 FILLER_45_734 ();
 sg13g2_fill_1 FILLER_45_738 ();
 sg13g2_fill_1 FILLER_45_766 ();
 sg13g2_fill_2 FILLER_45_795 ();
 sg13g2_decap_4 FILLER_45_828 ();
 sg13g2_fill_2 FILLER_45_917 ();
 sg13g2_fill_2 FILLER_45_969 ();
 sg13g2_decap_8 FILLER_45_989 ();
 sg13g2_decap_8 FILLER_45_996 ();
 sg13g2_fill_2 FILLER_45_1003 ();
 sg13g2_decap_4 FILLER_45_1036 ();
 sg13g2_fill_2 FILLER_45_1094 ();
 sg13g2_fill_2 FILLER_45_1115 ();
 sg13g2_fill_1 FILLER_45_1117 ();
 sg13g2_fill_1 FILLER_45_1150 ();
 sg13g2_fill_1 FILLER_45_1196 ();
 sg13g2_decap_8 FILLER_45_1225 ();
 sg13g2_decap_8 FILLER_45_1232 ();
 sg13g2_fill_1 FILLER_45_1271 ();
 sg13g2_decap_8 FILLER_45_1281 ();
 sg13g2_decap_8 FILLER_45_1288 ();
 sg13g2_decap_8 FILLER_45_1295 ();
 sg13g2_decap_8 FILLER_45_1302 ();
 sg13g2_decap_4 FILLER_45_1309 ();
 sg13g2_fill_2 FILLER_45_1313 ();
 sg13g2_decap_4 FILLER_46_0 ();
 sg13g2_fill_2 FILLER_46_55 ();
 sg13g2_fill_1 FILLER_46_75 ();
 sg13g2_decap_8 FILLER_46_103 ();
 sg13g2_fill_2 FILLER_46_110 ();
 sg13g2_decap_8 FILLER_46_122 ();
 sg13g2_fill_2 FILLER_46_129 ();
 sg13g2_decap_8 FILLER_46_135 ();
 sg13g2_decap_8 FILLER_46_142 ();
 sg13g2_decap_8 FILLER_46_149 ();
 sg13g2_fill_1 FILLER_46_165 ();
 sg13g2_fill_1 FILLER_46_184 ();
 sg13g2_fill_1 FILLER_46_191 ();
 sg13g2_decap_8 FILLER_46_257 ();
 sg13g2_fill_1 FILLER_46_264 ();
 sg13g2_fill_1 FILLER_46_278 ();
 sg13g2_fill_2 FILLER_46_283 ();
 sg13g2_fill_1 FILLER_46_285 ();
 sg13g2_fill_1 FILLER_46_355 ();
 sg13g2_fill_1 FILLER_46_365 ();
 sg13g2_fill_2 FILLER_46_404 ();
 sg13g2_fill_2 FILLER_46_433 ();
 sg13g2_fill_1 FILLER_46_448 ();
 sg13g2_decap_4 FILLER_46_508 ();
 sg13g2_fill_1 FILLER_46_525 ();
 sg13g2_fill_2 FILLER_46_562 ();
 sg13g2_fill_1 FILLER_46_564 ();
 sg13g2_decap_4 FILLER_46_641 ();
 sg13g2_fill_1 FILLER_46_645 ();
 sg13g2_fill_2 FILLER_46_655 ();
 sg13g2_fill_1 FILLER_46_657 ();
 sg13g2_decap_4 FILLER_46_662 ();
 sg13g2_fill_2 FILLER_46_666 ();
 sg13g2_decap_8 FILLER_46_681 ();
 sg13g2_fill_1 FILLER_46_688 ();
 sg13g2_decap_8 FILLER_46_729 ();
 sg13g2_decap_4 FILLER_46_736 ();
 sg13g2_fill_2 FILLER_46_748 ();
 sg13g2_fill_2 FILLER_46_782 ();
 sg13g2_fill_1 FILLER_46_810 ();
 sg13g2_decap_8 FILLER_46_826 ();
 sg13g2_decap_8 FILLER_46_833 ();
 sg13g2_fill_2 FILLER_46_840 ();
 sg13g2_fill_1 FILLER_46_842 ();
 sg13g2_fill_2 FILLER_46_853 ();
 sg13g2_fill_1 FILLER_46_861 ();
 sg13g2_fill_1 FILLER_46_875 ();
 sg13g2_fill_2 FILLER_46_981 ();
 sg13g2_fill_1 FILLER_46_1000 ();
 sg13g2_decap_8 FILLER_46_1037 ();
 sg13g2_decap_4 FILLER_46_1044 ();
 sg13g2_fill_2 FILLER_46_1048 ();
 sg13g2_fill_1 FILLER_46_1097 ();
 sg13g2_decap_8 FILLER_46_1111 ();
 sg13g2_decap_4 FILLER_46_1118 ();
 sg13g2_fill_1 FILLER_46_1122 ();
 sg13g2_fill_1 FILLER_46_1162 ();
 sg13g2_decap_4 FILLER_46_1177 ();
 sg13g2_fill_1 FILLER_46_1186 ();
 sg13g2_fill_1 FILLER_46_1205 ();
 sg13g2_fill_1 FILLER_46_1242 ();
 sg13g2_fill_2 FILLER_46_1260 ();
 sg13g2_decap_8 FILLER_46_1270 ();
 sg13g2_decap_8 FILLER_46_1277 ();
 sg13g2_decap_8 FILLER_46_1284 ();
 sg13g2_decap_8 FILLER_46_1291 ();
 sg13g2_decap_8 FILLER_46_1298 ();
 sg13g2_decap_8 FILLER_46_1305 ();
 sg13g2_fill_2 FILLER_46_1312 ();
 sg13g2_fill_1 FILLER_46_1314 ();
 sg13g2_decap_4 FILLER_47_0 ();
 sg13g2_fill_2 FILLER_47_36 ();
 sg13g2_fill_2 FILLER_47_71 ();
 sg13g2_fill_2 FILLER_47_112 ();
 sg13g2_fill_1 FILLER_47_114 ();
 sg13g2_decap_8 FILLER_47_131 ();
 sg13g2_decap_8 FILLER_47_138 ();
 sg13g2_decap_4 FILLER_47_145 ();
 sg13g2_fill_2 FILLER_47_149 ();
 sg13g2_decap_8 FILLER_47_155 ();
 sg13g2_fill_1 FILLER_47_162 ();
 sg13g2_fill_2 FILLER_47_196 ();
 sg13g2_fill_1 FILLER_47_198 ();
 sg13g2_fill_1 FILLER_47_204 ();
 sg13g2_fill_1 FILLER_47_234 ();
 sg13g2_decap_4 FILLER_47_257 ();
 sg13g2_fill_1 FILLER_47_261 ();
 sg13g2_fill_1 FILLER_47_386 ();
 sg13g2_decap_4 FILLER_47_396 ();
 sg13g2_fill_1 FILLER_47_446 ();
 sg13g2_decap_4 FILLER_47_489 ();
 sg13g2_fill_1 FILLER_47_573 ();
 sg13g2_fill_1 FILLER_47_587 ();
 sg13g2_fill_2 FILLER_47_606 ();
 sg13g2_fill_1 FILLER_47_608 ();
 sg13g2_fill_2 FILLER_47_688 ();
 sg13g2_fill_1 FILLER_47_690 ();
 sg13g2_fill_2 FILLER_47_732 ();
 sg13g2_fill_1 FILLER_47_734 ();
 sg13g2_fill_1 FILLER_47_789 ();
 sg13g2_fill_2 FILLER_47_803 ();
 sg13g2_fill_1 FILLER_47_823 ();
 sg13g2_decap_8 FILLER_47_833 ();
 sg13g2_decap_8 FILLER_47_840 ();
 sg13g2_fill_1 FILLER_47_847 ();
 sg13g2_fill_1 FILLER_47_889 ();
 sg13g2_fill_2 FILLER_47_900 ();
 sg13g2_decap_8 FILLER_47_915 ();
 sg13g2_fill_2 FILLER_47_926 ();
 sg13g2_fill_1 FILLER_47_928 ();
 sg13g2_fill_2 FILLER_47_955 ();
 sg13g2_fill_1 FILLER_47_985 ();
 sg13g2_fill_2 FILLER_47_1018 ();
 sg13g2_fill_1 FILLER_47_1020 ();
 sg13g2_fill_1 FILLER_47_1043 ();
 sg13g2_fill_1 FILLER_47_1084 ();
 sg13g2_fill_2 FILLER_47_1094 ();
 sg13g2_fill_1 FILLER_47_1096 ();
 sg13g2_fill_1 FILLER_47_1116 ();
 sg13g2_fill_2 FILLER_47_1138 ();
 sg13g2_fill_1 FILLER_47_1140 ();
 sg13g2_fill_1 FILLER_47_1213 ();
 sg13g2_decap_8 FILLER_47_1245 ();
 sg13g2_fill_1 FILLER_47_1252 ();
 sg13g2_decap_8 FILLER_47_1280 ();
 sg13g2_decap_8 FILLER_47_1287 ();
 sg13g2_decap_8 FILLER_47_1294 ();
 sg13g2_decap_8 FILLER_47_1301 ();
 sg13g2_decap_8 FILLER_47_1308 ();
 sg13g2_decap_4 FILLER_48_0 ();
 sg13g2_fill_2 FILLER_48_4 ();
 sg13g2_fill_2 FILLER_48_34 ();
 sg13g2_fill_2 FILLER_48_58 ();
 sg13g2_fill_1 FILLER_48_60 ();
 sg13g2_fill_2 FILLER_48_75 ();
 sg13g2_fill_2 FILLER_48_91 ();
 sg13g2_fill_1 FILLER_48_93 ();
 sg13g2_fill_1 FILLER_48_115 ();
 sg13g2_fill_1 FILLER_48_122 ();
 sg13g2_fill_1 FILLER_48_132 ();
 sg13g2_fill_1 FILLER_48_173 ();
 sg13g2_fill_2 FILLER_48_188 ();
 sg13g2_decap_8 FILLER_48_228 ();
 sg13g2_decap_8 FILLER_48_235 ();
 sg13g2_decap_8 FILLER_48_242 ();
 sg13g2_fill_2 FILLER_48_249 ();
 sg13g2_fill_2 FILLER_48_287 ();
 sg13g2_fill_1 FILLER_48_289 ();
 sg13g2_fill_1 FILLER_48_296 ();
 sg13g2_fill_2 FILLER_48_332 ();
 sg13g2_fill_1 FILLER_48_334 ();
 sg13g2_decap_4 FILLER_48_348 ();
 sg13g2_fill_2 FILLER_48_379 ();
 sg13g2_fill_1 FILLER_48_381 ();
 sg13g2_decap_4 FILLER_48_386 ();
 sg13g2_fill_2 FILLER_48_401 ();
 sg13g2_fill_2 FILLER_48_450 ();
 sg13g2_fill_1 FILLER_48_452 ();
 sg13g2_fill_1 FILLER_48_458 ();
 sg13g2_fill_1 FILLER_48_467 ();
 sg13g2_decap_4 FILLER_48_477 ();
 sg13g2_fill_1 FILLER_48_481 ();
 sg13g2_decap_4 FILLER_48_524 ();
 sg13g2_fill_2 FILLER_48_528 ();
 sg13g2_fill_2 FILLER_48_535 ();
 sg13g2_fill_2 FILLER_48_547 ();
 sg13g2_fill_1 FILLER_48_549 ();
 sg13g2_fill_2 FILLER_48_606 ();
 sg13g2_fill_1 FILLER_48_608 ();
 sg13g2_decap_8 FILLER_48_654 ();
 sg13g2_fill_2 FILLER_48_661 ();
 sg13g2_fill_1 FILLER_48_663 ();
 sg13g2_fill_2 FILLER_48_677 ();
 sg13g2_decap_8 FILLER_48_692 ();
 sg13g2_decap_8 FILLER_48_699 ();
 sg13g2_fill_1 FILLER_48_706 ();
 sg13g2_fill_2 FILLER_48_724 ();
 sg13g2_fill_2 FILLER_48_781 ();
 sg13g2_fill_1 FILLER_48_783 ();
 sg13g2_fill_2 FILLER_48_855 ();
 sg13g2_decap_8 FILLER_48_865 ();
 sg13g2_fill_2 FILLER_48_890 ();
 sg13g2_decap_8 FILLER_48_905 ();
 sg13g2_decap_8 FILLER_48_912 ();
 sg13g2_decap_4 FILLER_48_919 ();
 sg13g2_fill_1 FILLER_48_932 ();
 sg13g2_fill_2 FILLER_48_937 ();
 sg13g2_fill_1 FILLER_48_983 ();
 sg13g2_fill_1 FILLER_48_1011 ();
 sg13g2_decap_4 FILLER_48_1036 ();
 sg13g2_decap_4 FILLER_48_1049 ();
 sg13g2_fill_2 FILLER_48_1053 ();
 sg13g2_fill_2 FILLER_48_1072 ();
 sg13g2_decap_8 FILLER_48_1085 ();
 sg13g2_fill_2 FILLER_48_1133 ();
 sg13g2_decap_8 FILLER_48_1176 ();
 sg13g2_fill_2 FILLER_48_1183 ();
 sg13g2_fill_1 FILLER_48_1185 ();
 sg13g2_fill_1 FILLER_48_1194 ();
 sg13g2_decap_8 FILLER_48_1272 ();
 sg13g2_decap_8 FILLER_48_1279 ();
 sg13g2_decap_8 FILLER_48_1286 ();
 sg13g2_decap_8 FILLER_48_1293 ();
 sg13g2_decap_8 FILLER_48_1300 ();
 sg13g2_decap_8 FILLER_48_1307 ();
 sg13g2_fill_1 FILLER_48_1314 ();
 sg13g2_decap_8 FILLER_49_0 ();
 sg13g2_decap_4 FILLER_49_7 ();
 sg13g2_fill_1 FILLER_49_15 ();
 sg13g2_fill_1 FILLER_49_40 ();
 sg13g2_fill_2 FILLER_49_50 ();
 sg13g2_fill_1 FILLER_49_68 ();
 sg13g2_fill_2 FILLER_49_83 ();
 sg13g2_fill_1 FILLER_49_149 ();
 sg13g2_fill_1 FILLER_49_190 ();
 sg13g2_decap_8 FILLER_49_232 ();
 sg13g2_decap_8 FILLER_49_239 ();
 sg13g2_fill_2 FILLER_49_246 ();
 sg13g2_fill_1 FILLER_49_248 ();
 sg13g2_fill_2 FILLER_49_254 ();
 sg13g2_fill_2 FILLER_49_292 ();
 sg13g2_fill_2 FILLER_49_304 ();
 sg13g2_fill_2 FILLER_49_311 ();
 sg13g2_fill_1 FILLER_49_313 ();
 sg13g2_fill_2 FILLER_49_327 ();
 sg13g2_fill_1 FILLER_49_329 ();
 sg13g2_fill_2 FILLER_49_335 ();
 sg13g2_fill_2 FILLER_49_341 ();
 sg13g2_fill_1 FILLER_49_384 ();
 sg13g2_decap_8 FILLER_49_412 ();
 sg13g2_decap_8 FILLER_49_451 ();
 sg13g2_decap_8 FILLER_49_458 ();
 sg13g2_decap_4 FILLER_49_465 ();
 sg13g2_fill_2 FILLER_49_469 ();
 sg13g2_fill_1 FILLER_49_480 ();
 sg13g2_fill_1 FILLER_49_486 ();
 sg13g2_fill_2 FILLER_49_509 ();
 sg13g2_fill_2 FILLER_49_543 ();
 sg13g2_fill_1 FILLER_49_549 ();
 sg13g2_fill_1 FILLER_49_555 ();
 sg13g2_fill_1 FILLER_49_560 ();
 sg13g2_fill_2 FILLER_49_593 ();
 sg13g2_fill_1 FILLER_49_595 ();
 sg13g2_fill_2 FILLER_49_622 ();
 sg13g2_fill_1 FILLER_49_624 ();
 sg13g2_fill_2 FILLER_49_630 ();
 sg13g2_fill_1 FILLER_49_637 ();
 sg13g2_fill_1 FILLER_49_644 ();
 sg13g2_decap_4 FILLER_49_654 ();
 sg13g2_fill_2 FILLER_49_658 ();
 sg13g2_decap_8 FILLER_49_700 ();
 sg13g2_decap_8 FILLER_49_707 ();
 sg13g2_decap_8 FILLER_49_714 ();
 sg13g2_fill_2 FILLER_49_721 ();
 sg13g2_fill_1 FILLER_49_723 ();
 sg13g2_fill_2 FILLER_49_754 ();
 sg13g2_fill_1 FILLER_49_756 ();
 sg13g2_fill_1 FILLER_49_854 ();
 sg13g2_fill_2 FILLER_49_868 ();
 sg13g2_fill_1 FILLER_49_870 ();
 sg13g2_fill_2 FILLER_49_987 ();
 sg13g2_fill_1 FILLER_49_989 ();
 sg13g2_fill_1 FILLER_49_1000 ();
 sg13g2_fill_1 FILLER_49_1016 ();
 sg13g2_fill_1 FILLER_49_1049 ();
 sg13g2_decap_4 FILLER_49_1056 ();
 sg13g2_fill_1 FILLER_49_1060 ();
 sg13g2_decap_8 FILLER_49_1074 ();
 sg13g2_fill_2 FILLER_49_1137 ();
 sg13g2_fill_1 FILLER_49_1139 ();
 sg13g2_decap_8 FILLER_49_1171 ();
 sg13g2_decap_8 FILLER_49_1178 ();
 sg13g2_fill_1 FILLER_49_1185 ();
 sg13g2_fill_2 FILLER_49_1226 ();
 sg13g2_fill_2 FILLER_49_1242 ();
 sg13g2_fill_1 FILLER_49_1272 ();
 sg13g2_decap_8 FILLER_49_1282 ();
 sg13g2_decap_8 FILLER_49_1289 ();
 sg13g2_decap_8 FILLER_49_1296 ();
 sg13g2_decap_8 FILLER_49_1303 ();
 sg13g2_decap_4 FILLER_49_1310 ();
 sg13g2_fill_1 FILLER_49_1314 ();
 sg13g2_decap_8 FILLER_50_0 ();
 sg13g2_fill_1 FILLER_50_53 ();
 sg13g2_fill_1 FILLER_50_136 ();
 sg13g2_decap_8 FILLER_50_158 ();
 sg13g2_fill_1 FILLER_50_165 ();
 sg13g2_fill_1 FILLER_50_186 ();
 sg13g2_decap_8 FILLER_50_192 ();
 sg13g2_decap_4 FILLER_50_199 ();
 sg13g2_decap_4 FILLER_50_219 ();
 sg13g2_decap_8 FILLER_50_241 ();
 sg13g2_decap_8 FILLER_50_248 ();
 sg13g2_fill_2 FILLER_50_255 ();
 sg13g2_fill_1 FILLER_50_257 ();
 sg13g2_fill_2 FILLER_50_306 ();
 sg13g2_fill_1 FILLER_50_308 ();
 sg13g2_decap_8 FILLER_50_314 ();
 sg13g2_fill_2 FILLER_50_321 ();
 sg13g2_fill_1 FILLER_50_323 ();
 sg13g2_fill_2 FILLER_50_351 ();
 sg13g2_fill_2 FILLER_50_370 ();
 sg13g2_fill_1 FILLER_50_372 ();
 sg13g2_decap_4 FILLER_50_434 ();
 sg13g2_fill_1 FILLER_50_455 ();
 sg13g2_decap_4 FILLER_50_461 ();
 sg13g2_fill_1 FILLER_50_465 ();
 sg13g2_fill_1 FILLER_50_470 ();
 sg13g2_fill_1 FILLER_50_512 ();
 sg13g2_fill_2 FILLER_50_549 ();
 sg13g2_fill_1 FILLER_50_587 ();
 sg13g2_fill_2 FILLER_50_628 ();
 sg13g2_fill_1 FILLER_50_630 ();
 sg13g2_fill_2 FILLER_50_667 ();
 sg13g2_fill_2 FILLER_50_696 ();
 sg13g2_fill_1 FILLER_50_698 ();
 sg13g2_decap_4 FILLER_50_703 ();
 sg13g2_fill_2 FILLER_50_707 ();
 sg13g2_fill_2 FILLER_50_722 ();
 sg13g2_fill_2 FILLER_50_751 ();
 sg13g2_fill_1 FILLER_50_781 ();
 sg13g2_fill_2 FILLER_50_787 ();
 sg13g2_fill_1 FILLER_50_789 ();
 sg13g2_fill_1 FILLER_50_846 ();
 sg13g2_fill_2 FILLER_50_853 ();
 sg13g2_fill_1 FILLER_50_855 ();
 sg13g2_fill_1 FILLER_50_869 ();
 sg13g2_fill_1 FILLER_50_897 ();
 sg13g2_fill_2 FILLER_50_911 ();
 sg13g2_decap_8 FILLER_50_992 ();
 sg13g2_fill_1 FILLER_50_999 ();
 sg13g2_fill_2 FILLER_50_1004 ();
 sg13g2_fill_2 FILLER_50_1092 ();
 sg13g2_fill_1 FILLER_50_1094 ();
 sg13g2_fill_2 FILLER_50_1163 ();
 sg13g2_fill_1 FILLER_50_1192 ();
 sg13g2_fill_1 FILLER_50_1232 ();
 sg13g2_fill_2 FILLER_50_1264 ();
 sg13g2_fill_1 FILLER_50_1266 ();
 sg13g2_fill_1 FILLER_50_1271 ();
 sg13g2_decap_8 FILLER_50_1276 ();
 sg13g2_decap_8 FILLER_50_1283 ();
 sg13g2_decap_8 FILLER_50_1290 ();
 sg13g2_decap_8 FILLER_50_1297 ();
 sg13g2_decap_8 FILLER_50_1304 ();
 sg13g2_decap_4 FILLER_50_1311 ();
 sg13g2_decap_4 FILLER_51_0 ();
 sg13g2_decap_4 FILLER_51_40 ();
 sg13g2_fill_2 FILLER_51_57 ();
 sg13g2_fill_1 FILLER_51_59 ();
 sg13g2_fill_2 FILLER_51_73 ();
 sg13g2_fill_2 FILLER_51_83 ();
 sg13g2_fill_2 FILLER_51_110 ();
 sg13g2_fill_2 FILLER_51_117 ();
 sg13g2_decap_4 FILLER_51_137 ();
 sg13g2_fill_1 FILLER_51_141 ();
 sg13g2_fill_2 FILLER_51_155 ();
 sg13g2_fill_1 FILLER_51_171 ();
 sg13g2_decap_8 FILLER_51_192 ();
 sg13g2_fill_2 FILLER_51_199 ();
 sg13g2_decap_8 FILLER_51_221 ();
 sg13g2_decap_4 FILLER_51_228 ();
 sg13g2_decap_4 FILLER_51_244 ();
 sg13g2_decap_4 FILLER_51_261 ();
 sg13g2_fill_2 FILLER_51_292 ();
 sg13g2_decap_8 FILLER_51_307 ();
 sg13g2_fill_2 FILLER_51_318 ();
 sg13g2_fill_1 FILLER_51_320 ();
 sg13g2_fill_2 FILLER_51_368 ();
 sg13g2_fill_1 FILLER_51_370 ();
 sg13g2_fill_1 FILLER_51_386 ();
 sg13g2_fill_1 FILLER_51_392 ();
 sg13g2_fill_2 FILLER_51_399 ();
 sg13g2_fill_1 FILLER_51_401 ();
 sg13g2_decap_8 FILLER_51_442 ();
 sg13g2_fill_1 FILLER_51_449 ();
 sg13g2_fill_1 FILLER_51_523 ();
 sg13g2_fill_2 FILLER_51_538 ();
 sg13g2_fill_1 FILLER_51_549 ();
 sg13g2_fill_2 FILLER_51_603 ();
 sg13g2_fill_2 FILLER_51_631 ();
 sg13g2_fill_2 FILLER_51_666 ();
 sg13g2_fill_1 FILLER_51_668 ();
 sg13g2_decap_4 FILLER_51_690 ();
 sg13g2_decap_4 FILLER_51_722 ();
 sg13g2_fill_1 FILLER_51_726 ();
 sg13g2_fill_2 FILLER_51_732 ();
 sg13g2_fill_2 FILLER_51_806 ();
 sg13g2_fill_1 FILLER_51_808 ();
 sg13g2_fill_2 FILLER_51_818 ();
 sg13g2_fill_1 FILLER_51_820 ();
 sg13g2_fill_1 FILLER_51_868 ();
 sg13g2_fill_2 FILLER_51_897 ();
 sg13g2_fill_1 FILLER_51_899 ();
 sg13g2_decap_8 FILLER_51_995 ();
 sg13g2_decap_8 FILLER_51_1002 ();
 sg13g2_decap_4 FILLER_51_1009 ();
 sg13g2_decap_8 FILLER_51_1075 ();
 sg13g2_decap_8 FILLER_51_1082 ();
 sg13g2_decap_8 FILLER_51_1089 ();
 sg13g2_fill_1 FILLER_51_1096 ();
 sg13g2_fill_2 FILLER_51_1106 ();
 sg13g2_fill_1 FILLER_51_1153 ();
 sg13g2_fill_1 FILLER_51_1187 ();
 sg13g2_fill_2 FILLER_51_1199 ();
 sg13g2_fill_1 FILLER_51_1201 ();
 sg13g2_fill_2 FILLER_51_1233 ();
 sg13g2_fill_2 FILLER_51_1245 ();
 sg13g2_decap_8 FILLER_51_1294 ();
 sg13g2_decap_8 FILLER_51_1301 ();
 sg13g2_decap_8 FILLER_51_1308 ();
 sg13g2_decap_4 FILLER_52_0 ();
 sg13g2_fill_2 FILLER_52_4 ();
 sg13g2_fill_2 FILLER_52_46 ();
 sg13g2_fill_2 FILLER_52_75 ();
 sg13g2_fill_1 FILLER_52_77 ();
 sg13g2_fill_2 FILLER_52_87 ();
 sg13g2_fill_1 FILLER_52_125 ();
 sg13g2_decap_8 FILLER_52_130 ();
 sg13g2_fill_2 FILLER_52_137 ();
 sg13g2_fill_2 FILLER_52_166 ();
 sg13g2_fill_2 FILLER_52_179 ();
 sg13g2_fill_2 FILLER_52_191 ();
 sg13g2_decap_8 FILLER_52_198 ();
 sg13g2_fill_2 FILLER_52_205 ();
 sg13g2_decap_4 FILLER_52_223 ();
 sg13g2_fill_2 FILLER_52_227 ();
 sg13g2_fill_2 FILLER_52_314 ();
 sg13g2_fill_2 FILLER_52_326 ();
 sg13g2_fill_1 FILLER_52_328 ();
 sg13g2_fill_2 FILLER_52_338 ();
 sg13g2_fill_2 FILLER_52_357 ();
 sg13g2_fill_1 FILLER_52_407 ();
 sg13g2_fill_2 FILLER_52_507 ();
 sg13g2_fill_1 FILLER_52_522 ();
 sg13g2_decap_4 FILLER_52_550 ();
 sg13g2_fill_1 FILLER_52_554 ();
 sg13g2_fill_2 FILLER_52_563 ();
 sg13g2_decap_8 FILLER_52_606 ();
 sg13g2_fill_2 FILLER_52_613 ();
 sg13g2_fill_1 FILLER_52_615 ();
 sg13g2_fill_1 FILLER_52_657 ();
 sg13g2_fill_2 FILLER_52_667 ();
 sg13g2_fill_1 FILLER_52_669 ();
 sg13g2_decap_8 FILLER_52_688 ();
 sg13g2_decap_8 FILLER_52_708 ();
 sg13g2_fill_1 FILLER_52_782 ();
 sg13g2_fill_2 FILLER_52_821 ();
 sg13g2_fill_1 FILLER_52_823 ();
 sg13g2_decap_8 FILLER_52_857 ();
 sg13g2_fill_2 FILLER_52_864 ();
 sg13g2_fill_2 FILLER_52_883 ();
 sg13g2_fill_1 FILLER_52_885 ();
 sg13g2_fill_2 FILLER_52_904 ();
 sg13g2_fill_1 FILLER_52_906 ();
 sg13g2_fill_2 FILLER_52_940 ();
 sg13g2_fill_1 FILLER_52_942 ();
 sg13g2_decap_4 FILLER_52_973 ();
 sg13g2_fill_2 FILLER_52_1018 ();
 sg13g2_fill_1 FILLER_52_1028 ();
 sg13g2_fill_2 FILLER_52_1056 ();
 sg13g2_fill_2 FILLER_52_1099 ();
 sg13g2_fill_1 FILLER_52_1101 ();
 sg13g2_decap_8 FILLER_52_1106 ();
 sg13g2_fill_1 FILLER_52_1117 ();
 sg13g2_fill_1 FILLER_52_1158 ();
 sg13g2_fill_2 FILLER_52_1206 ();
 sg13g2_fill_1 FILLER_52_1208 ();
 sg13g2_fill_2 FILLER_52_1236 ();
 sg13g2_fill_1 FILLER_52_1262 ();
 sg13g2_decap_4 FILLER_52_1275 ();
 sg13g2_fill_1 FILLER_52_1279 ();
 sg13g2_decap_8 FILLER_52_1289 ();
 sg13g2_decap_8 FILLER_52_1296 ();
 sg13g2_decap_8 FILLER_52_1303 ();
 sg13g2_decap_4 FILLER_52_1310 ();
 sg13g2_fill_1 FILLER_52_1314 ();
 sg13g2_decap_8 FILLER_53_0 ();
 sg13g2_decap_4 FILLER_53_7 ();
 sg13g2_fill_1 FILLER_53_11 ();
 sg13g2_decap_4 FILLER_53_48 ();
 sg13g2_fill_2 FILLER_53_79 ();
 sg13g2_decap_4 FILLER_53_114 ();
 sg13g2_fill_1 FILLER_53_118 ();
 sg13g2_decap_4 FILLER_53_132 ();
 sg13g2_fill_1 FILLER_53_136 ();
 sg13g2_fill_1 FILLER_53_155 ();
 sg13g2_fill_2 FILLER_53_165 ();
 sg13g2_fill_1 FILLER_53_167 ();
 sg13g2_decap_4 FILLER_53_192 ();
 sg13g2_fill_2 FILLER_53_239 ();
 sg13g2_fill_1 FILLER_53_241 ();
 sg13g2_decap_8 FILLER_53_245 ();
 sg13g2_decap_4 FILLER_53_252 ();
 sg13g2_fill_1 FILLER_53_256 ();
 sg13g2_fill_1 FILLER_53_333 ();
 sg13g2_fill_2 FILLER_53_348 ();
 sg13g2_fill_2 FILLER_53_423 ();
 sg13g2_fill_1 FILLER_53_434 ();
 sg13g2_fill_1 FILLER_53_467 ();
 sg13g2_fill_2 FILLER_53_495 ();
 sg13g2_fill_1 FILLER_53_497 ();
 sg13g2_decap_8 FILLER_53_527 ();
 sg13g2_fill_2 FILLER_53_534 ();
 sg13g2_decap_4 FILLER_53_540 ();
 sg13g2_fill_1 FILLER_53_544 ();
 sg13g2_fill_2 FILLER_53_590 ();
 sg13g2_fill_1 FILLER_53_592 ();
 sg13g2_decap_8 FILLER_53_597 ();
 sg13g2_decap_4 FILLER_53_617 ();
 sg13g2_fill_2 FILLER_53_625 ();
 sg13g2_fill_1 FILLER_53_627 ();
 sg13g2_decap_8 FILLER_53_684 ();
 sg13g2_decap_8 FILLER_53_691 ();
 sg13g2_fill_2 FILLER_53_707 ();
 sg13g2_fill_1 FILLER_53_709 ();
 sg13g2_fill_2 FILLER_53_737 ();
 sg13g2_fill_1 FILLER_53_739 ();
 sg13g2_fill_2 FILLER_53_772 ();
 sg13g2_fill_2 FILLER_53_801 ();
 sg13g2_fill_1 FILLER_53_803 ();
 sg13g2_fill_2 FILLER_53_817 ();
 sg13g2_fill_2 FILLER_53_824 ();
 sg13g2_fill_1 FILLER_53_826 ();
 sg13g2_fill_2 FILLER_53_836 ();
 sg13g2_fill_1 FILLER_53_838 ();
 sg13g2_fill_1 FILLER_53_866 ();
 sg13g2_fill_2 FILLER_53_930 ();
 sg13g2_fill_1 FILLER_53_932 ();
 sg13g2_fill_1 FILLER_53_946 ();
 sg13g2_decap_8 FILLER_53_959 ();
 sg13g2_decap_4 FILLER_53_966 ();
 sg13g2_decap_4 FILLER_53_1024 ();
 sg13g2_fill_2 FILLER_53_1036 ();
 sg13g2_fill_1 FILLER_53_1060 ();
 sg13g2_fill_2 FILLER_53_1070 ();
 sg13g2_fill_1 FILLER_53_1077 ();
 sg13g2_fill_2 FILLER_53_1104 ();
 sg13g2_decap_8 FILLER_53_1110 ();
 sg13g2_decap_4 FILLER_53_1117 ();
 sg13g2_fill_2 FILLER_53_1121 ();
 sg13g2_fill_1 FILLER_53_1131 ();
 sg13g2_fill_2 FILLER_53_1159 ();
 sg13g2_fill_2 FILLER_53_1175 ();
 sg13g2_fill_1 FILLER_53_1177 ();
 sg13g2_fill_2 FILLER_53_1187 ();
 sg13g2_fill_1 FILLER_53_1198 ();
 sg13g2_fill_2 FILLER_53_1212 ();
 sg13g2_decap_8 FILLER_53_1291 ();
 sg13g2_decap_8 FILLER_53_1298 ();
 sg13g2_decap_8 FILLER_53_1305 ();
 sg13g2_fill_2 FILLER_53_1312 ();
 sg13g2_fill_1 FILLER_53_1314 ();
 sg13g2_decap_4 FILLER_54_0 ();
 sg13g2_fill_2 FILLER_54_4 ();
 sg13g2_fill_2 FILLER_54_46 ();
 sg13g2_fill_2 FILLER_54_61 ();
 sg13g2_fill_1 FILLER_54_67 ();
 sg13g2_fill_2 FILLER_54_78 ();
 sg13g2_fill_1 FILLER_54_80 ();
 sg13g2_decap_4 FILLER_54_108 ();
 sg13g2_fill_2 FILLER_54_112 ();
 sg13g2_fill_1 FILLER_54_118 ();
 sg13g2_fill_1 FILLER_54_124 ();
 sg13g2_decap_4 FILLER_54_135 ();
 sg13g2_fill_1 FILLER_54_139 ();
 sg13g2_fill_1 FILLER_54_147 ();
 sg13g2_fill_1 FILLER_54_181 ();
 sg13g2_decap_4 FILLER_54_189 ();
 sg13g2_fill_1 FILLER_54_229 ();
 sg13g2_decap_4 FILLER_54_253 ();
 sg13g2_fill_1 FILLER_54_257 ();
 sg13g2_fill_1 FILLER_54_266 ();
 sg13g2_fill_1 FILLER_54_277 ();
 sg13g2_fill_1 FILLER_54_297 ();
 sg13g2_fill_2 FILLER_54_327 ();
 sg13g2_fill_2 FILLER_54_383 ();
 sg13g2_fill_2 FILLER_54_421 ();
 sg13g2_fill_1 FILLER_54_460 ();
 sg13g2_fill_2 FILLER_54_519 ();
 sg13g2_fill_1 FILLER_54_521 ();
 sg13g2_decap_4 FILLER_54_567 ();
 sg13g2_fill_1 FILLER_54_571 ();
 sg13g2_fill_1 FILLER_54_589 ();
 sg13g2_decap_8 FILLER_54_599 ();
 sg13g2_decap_8 FILLER_54_606 ();
 sg13g2_fill_2 FILLER_54_617 ();
 sg13g2_fill_2 FILLER_54_637 ();
 sg13g2_fill_1 FILLER_54_639 ();
 sg13g2_fill_2 FILLER_54_653 ();
 sg13g2_fill_1 FILLER_54_655 ();
 sg13g2_decap_4 FILLER_54_692 ();
 sg13g2_fill_2 FILLER_54_696 ();
 sg13g2_fill_2 FILLER_54_711 ();
 sg13g2_fill_1 FILLER_54_713 ();
 sg13g2_fill_2 FILLER_54_732 ();
 sg13g2_fill_1 FILLER_54_734 ();
 sg13g2_fill_1 FILLER_54_754 ();
 sg13g2_decap_8 FILLER_54_761 ();
 sg13g2_decap_8 FILLER_54_768 ();
 sg13g2_fill_2 FILLER_54_829 ();
 sg13g2_fill_1 FILLER_54_831 ();
 sg13g2_fill_1 FILLER_54_836 ();
 sg13g2_decap_4 FILLER_54_845 ();
 sg13g2_fill_2 FILLER_54_952 ();
 sg13g2_fill_1 FILLER_54_954 ();
 sg13g2_fill_2 FILLER_54_968 ();
 sg13g2_fill_1 FILLER_54_970 ();
 sg13g2_fill_1 FILLER_54_1071 ();
 sg13g2_fill_2 FILLER_54_1099 ();
 sg13g2_fill_2 FILLER_54_1141 ();
 sg13g2_fill_2 FILLER_54_1156 ();
 sg13g2_fill_1 FILLER_54_1158 ();
 sg13g2_fill_1 FILLER_54_1192 ();
 sg13g2_fill_2 FILLER_54_1212 ();
 sg13g2_fill_1 FILLER_54_1214 ();
 sg13g2_fill_2 FILLER_54_1244 ();
 sg13g2_fill_1 FILLER_54_1246 ();
 sg13g2_fill_2 FILLER_54_1253 ();
 sg13g2_fill_1 FILLER_54_1255 ();
 sg13g2_fill_1 FILLER_54_1265 ();
 sg13g2_decap_4 FILLER_54_1270 ();
 sg13g2_fill_1 FILLER_54_1274 ();
 sg13g2_decap_8 FILLER_54_1284 ();
 sg13g2_decap_8 FILLER_54_1291 ();
 sg13g2_decap_8 FILLER_54_1298 ();
 sg13g2_decap_8 FILLER_54_1305 ();
 sg13g2_fill_2 FILLER_54_1312 ();
 sg13g2_fill_1 FILLER_54_1314 ();
 sg13g2_fill_2 FILLER_55_0 ();
 sg13g2_fill_1 FILLER_55_36 ();
 sg13g2_decap_4 FILLER_55_103 ();
 sg13g2_fill_2 FILLER_55_107 ();
 sg13g2_decap_8 FILLER_55_154 ();
 sg13g2_fill_1 FILLER_55_165 ();
 sg13g2_fill_2 FILLER_55_176 ();
 sg13g2_fill_2 FILLER_55_185 ();
 sg13g2_fill_1 FILLER_55_187 ();
 sg13g2_fill_1 FILLER_55_206 ();
 sg13g2_decap_8 FILLER_55_259 ();
 sg13g2_decap_8 FILLER_55_266 ();
 sg13g2_fill_1 FILLER_55_296 ();
 sg13g2_fill_2 FILLER_55_306 ();
 sg13g2_fill_2 FILLER_55_313 ();
 sg13g2_fill_1 FILLER_55_315 ();
 sg13g2_fill_2 FILLER_55_322 ();
 sg13g2_fill_1 FILLER_55_333 ();
 sg13g2_fill_1 FILLER_55_394 ();
 sg13g2_fill_2 FILLER_55_431 ();
 sg13g2_fill_1 FILLER_55_433 ();
 sg13g2_decap_8 FILLER_55_463 ();
 sg13g2_fill_1 FILLER_55_470 ();
 sg13g2_decap_8 FILLER_55_507 ();
 sg13g2_decap_4 FILLER_55_514 ();
 sg13g2_fill_2 FILLER_55_518 ();
 sg13g2_decap_4 FILLER_55_560 ();
 sg13g2_fill_1 FILLER_55_564 ();
 sg13g2_decap_4 FILLER_55_576 ();
 sg13g2_fill_1 FILLER_55_580 ();
 sg13g2_fill_2 FILLER_55_621 ();
 sg13g2_fill_1 FILLER_55_629 ();
 sg13g2_fill_1 FILLER_55_663 ();
 sg13g2_fill_1 FILLER_55_699 ();
 sg13g2_fill_2 FILLER_55_748 ();
 sg13g2_fill_1 FILLER_55_750 ();
 sg13g2_fill_1 FILLER_55_759 ();
 sg13g2_decap_8 FILLER_55_773 ();
 sg13g2_fill_1 FILLER_55_780 ();
 sg13g2_fill_1 FILLER_55_816 ();
 sg13g2_decap_4 FILLER_55_821 ();
 sg13g2_fill_2 FILLER_55_825 ();
 sg13g2_decap_8 FILLER_55_835 ();
 sg13g2_decap_8 FILLER_55_842 ();
 sg13g2_decap_4 FILLER_55_849 ();
 sg13g2_decap_8 FILLER_55_863 ();
 sg13g2_fill_2 FILLER_55_870 ();
 sg13g2_fill_1 FILLER_55_872 ();
 sg13g2_fill_2 FILLER_55_912 ();
 sg13g2_fill_1 FILLER_55_919 ();
 sg13g2_fill_2 FILLER_55_956 ();
 sg13g2_fill_2 FILLER_55_997 ();
 sg13g2_fill_2 FILLER_55_1068 ();
 sg13g2_fill_1 FILLER_55_1070 ();
 sg13g2_fill_2 FILLER_55_1113 ();
 sg13g2_fill_1 FILLER_55_1120 ();
 sg13g2_fill_2 FILLER_55_1173 ();
 sg13g2_fill_1 FILLER_55_1175 ();
 sg13g2_decap_8 FILLER_55_1288 ();
 sg13g2_decap_8 FILLER_55_1295 ();
 sg13g2_decap_8 FILLER_55_1302 ();
 sg13g2_decap_4 FILLER_55_1309 ();
 sg13g2_fill_2 FILLER_55_1313 ();
 sg13g2_decap_8 FILLER_56_0 ();
 sg13g2_fill_2 FILLER_56_7 ();
 sg13g2_fill_1 FILLER_56_45 ();
 sg13g2_fill_1 FILLER_56_74 ();
 sg13g2_decap_4 FILLER_56_126 ();
 sg13g2_fill_2 FILLER_56_146 ();
 sg13g2_fill_2 FILLER_56_197 ();
 sg13g2_decap_8 FILLER_56_255 ();
 sg13g2_decap_8 FILLER_56_262 ();
 sg13g2_fill_2 FILLER_56_274 ();
 sg13g2_fill_2 FILLER_56_280 ();
 sg13g2_fill_1 FILLER_56_380 ();
 sg13g2_fill_1 FILLER_56_416 ();
 sg13g2_decap_8 FILLER_56_470 ();
 sg13g2_decap_4 FILLER_56_514 ();
 sg13g2_fill_1 FILLER_56_518 ();
 sg13g2_fill_2 FILLER_56_537 ();
 sg13g2_fill_1 FILLER_56_545 ();
 sg13g2_decap_4 FILLER_56_566 ();
 sg13g2_fill_2 FILLER_56_646 ();
 sg13g2_fill_1 FILLER_56_648 ();
 sg13g2_fill_1 FILLER_56_662 ();
 sg13g2_fill_2 FILLER_56_717 ();
 sg13g2_fill_1 FILLER_56_732 ();
 sg13g2_decap_4 FILLER_56_750 ();
 sg13g2_fill_2 FILLER_56_754 ();
 sg13g2_fill_1 FILLER_56_774 ();
 sg13g2_fill_1 FILLER_56_780 ();
 sg13g2_fill_2 FILLER_56_810 ();
 sg13g2_decap_4 FILLER_56_821 ();
 sg13g2_fill_2 FILLER_56_830 ();
 sg13g2_fill_1 FILLER_56_859 ();
 sg13g2_fill_2 FILLER_56_878 ();
 sg13g2_fill_1 FILLER_56_880 ();
 sg13g2_fill_2 FILLER_56_894 ();
 sg13g2_fill_1 FILLER_56_896 ();
 sg13g2_fill_2 FILLER_56_927 ();
 sg13g2_fill_2 FILLER_56_969 ();
 sg13g2_fill_1 FILLER_56_971 ();
 sg13g2_fill_1 FILLER_56_1049 ();
 sg13g2_fill_2 FILLER_56_1099 ();
 sg13g2_decap_8 FILLER_56_1138 ();
 sg13g2_fill_2 FILLER_56_1145 ();
 sg13g2_fill_1 FILLER_56_1192 ();
 sg13g2_fill_2 FILLER_56_1233 ();
 sg13g2_fill_1 FILLER_56_1235 ();
 sg13g2_decap_4 FILLER_56_1248 ();
 sg13g2_fill_1 FILLER_56_1261 ();
 sg13g2_fill_1 FILLER_56_1275 ();
 sg13g2_decap_8 FILLER_56_1285 ();
 sg13g2_decap_8 FILLER_56_1292 ();
 sg13g2_decap_8 FILLER_56_1299 ();
 sg13g2_decap_8 FILLER_56_1306 ();
 sg13g2_fill_2 FILLER_56_1313 ();
 sg13g2_decap_8 FILLER_57_0 ();
 sg13g2_decap_4 FILLER_57_7 ();
 sg13g2_fill_2 FILLER_57_59 ();
 sg13g2_fill_1 FILLER_57_74 ();
 sg13g2_fill_1 FILLER_57_89 ();
 sg13g2_fill_1 FILLER_57_155 ();
 sg13g2_fill_2 FILLER_57_181 ();
 sg13g2_decap_4 FILLER_57_210 ();
 sg13g2_decap_8 FILLER_57_241 ();
 sg13g2_decap_8 FILLER_57_248 ();
 sg13g2_decap_4 FILLER_57_255 ();
 sg13g2_fill_1 FILLER_57_259 ();
 sg13g2_fill_2 FILLER_57_300 ();
 sg13g2_fill_1 FILLER_57_302 ();
 sg13g2_fill_1 FILLER_57_308 ();
 sg13g2_decap_8 FILLER_57_317 ();
 sg13g2_decap_8 FILLER_57_324 ();
 sg13g2_fill_2 FILLER_57_331 ();
 sg13g2_fill_1 FILLER_57_333 ();
 sg13g2_fill_2 FILLER_57_343 ();
 sg13g2_fill_2 FILLER_57_371 ();
 sg13g2_fill_2 FILLER_57_382 ();
 sg13g2_fill_1 FILLER_57_384 ();
 sg13g2_decap_8 FILLER_57_467 ();
 sg13g2_decap_8 FILLER_57_524 ();
 sg13g2_fill_1 FILLER_57_531 ();
 sg13g2_fill_1 FILLER_57_599 ();
 sg13g2_decap_8 FILLER_57_649 ();
 sg13g2_decap_4 FILLER_57_656 ();
 sg13g2_fill_2 FILLER_57_660 ();
 sg13g2_fill_1 FILLER_57_667 ();
 sg13g2_fill_2 FILLER_57_672 ();
 sg13g2_fill_1 FILLER_57_712 ();
 sg13g2_fill_1 FILLER_57_726 ();
 sg13g2_fill_2 FILLER_57_787 ();
 sg13g2_fill_2 FILLER_57_794 ();
 sg13g2_fill_2 FILLER_57_814 ();
 sg13g2_fill_2 FILLER_57_852 ();
 sg13g2_fill_1 FILLER_57_854 ();
 sg13g2_decap_8 FILLER_57_890 ();
 sg13g2_decap_8 FILLER_57_897 ();
 sg13g2_decap_4 FILLER_57_904 ();
 sg13g2_fill_1 FILLER_57_950 ();
 sg13g2_fill_1 FILLER_57_970 ();
 sg13g2_decap_4 FILLER_57_976 ();
 sg13g2_fill_2 FILLER_57_1030 ();
 sg13g2_fill_1 FILLER_57_1032 ();
 sg13g2_fill_2 FILLER_57_1047 ();
 sg13g2_fill_2 FILLER_57_1095 ();
 sg13g2_fill_1 FILLER_57_1097 ();
 sg13g2_fill_2 FILLER_57_1107 ();
 sg13g2_fill_1 FILLER_57_1109 ();
 sg13g2_decap_8 FILLER_57_1123 ();
 sg13g2_decap_8 FILLER_57_1130 ();
 sg13g2_decap_4 FILLER_57_1137 ();
 sg13g2_fill_1 FILLER_57_1141 ();
 sg13g2_decap_8 FILLER_57_1229 ();
 sg13g2_decap_8 FILLER_57_1236 ();
 sg13g2_fill_2 FILLER_57_1243 ();
 sg13g2_fill_1 FILLER_57_1254 ();
 sg13g2_decap_8 FILLER_57_1282 ();
 sg13g2_decap_8 FILLER_57_1289 ();
 sg13g2_decap_8 FILLER_57_1296 ();
 sg13g2_decap_8 FILLER_57_1303 ();
 sg13g2_decap_4 FILLER_57_1310 ();
 sg13g2_fill_1 FILLER_57_1314 ();
 sg13g2_decap_8 FILLER_58_0 ();
 sg13g2_fill_2 FILLER_58_7 ();
 sg13g2_fill_1 FILLER_58_9 ();
 sg13g2_fill_1 FILLER_58_17 ();
 sg13g2_fill_2 FILLER_58_42 ();
 sg13g2_fill_1 FILLER_58_44 ();
 sg13g2_fill_2 FILLER_58_62 ();
 sg13g2_decap_4 FILLER_58_101 ();
 sg13g2_fill_2 FILLER_58_105 ();
 sg13g2_fill_2 FILLER_58_124 ();
 sg13g2_fill_1 FILLER_58_126 ();
 sg13g2_fill_1 FILLER_58_169 ();
 sg13g2_decap_4 FILLER_58_198 ();
 sg13g2_fill_2 FILLER_58_206 ();
 sg13g2_fill_1 FILLER_58_208 ();
 sg13g2_decap_8 FILLER_58_222 ();
 sg13g2_fill_1 FILLER_58_229 ();
 sg13g2_fill_1 FILLER_58_251 ();
 sg13g2_decap_8 FILLER_58_332 ();
 sg13g2_fill_2 FILLER_58_339 ();
 sg13g2_fill_1 FILLER_58_341 ();
 sg13g2_decap_4 FILLER_58_350 ();
 sg13g2_fill_2 FILLER_58_354 ();
 sg13g2_decap_8 FILLER_58_369 ();
 sg13g2_decap_4 FILLER_58_376 ();
 sg13g2_fill_1 FILLER_58_380 ();
 sg13g2_decap_4 FILLER_58_389 ();
 sg13g2_fill_1 FILLER_58_410 ();
 sg13g2_fill_1 FILLER_58_424 ();
 sg13g2_decap_8 FILLER_58_474 ();
 sg13g2_decap_4 FILLER_58_520 ();
 sg13g2_fill_2 FILLER_58_524 ();
 sg13g2_fill_2 FILLER_58_567 ();
 sg13g2_fill_2 FILLER_58_581 ();
 sg13g2_fill_1 FILLER_58_588 ();
 sg13g2_fill_2 FILLER_58_621 ();
 sg13g2_fill_1 FILLER_58_643 ();
 sg13g2_fill_2 FILLER_58_653 ();
 sg13g2_fill_2 FILLER_58_663 ();
 sg13g2_decap_8 FILLER_58_724 ();
 sg13g2_decap_8 FILLER_58_731 ();
 sg13g2_decap_4 FILLER_58_738 ();
 sg13g2_fill_2 FILLER_58_742 ();
 sg13g2_fill_2 FILLER_58_775 ();
 sg13g2_fill_2 FILLER_58_813 ();
 sg13g2_fill_1 FILLER_58_842 ();
 sg13g2_fill_2 FILLER_58_853 ();
 sg13g2_fill_1 FILLER_58_855 ();
 sg13g2_fill_1 FILLER_58_887 ();
 sg13g2_fill_1 FILLER_58_901 ();
 sg13g2_fill_2 FILLER_58_911 ();
 sg13g2_fill_1 FILLER_58_927 ();
 sg13g2_fill_1 FILLER_58_996 ();
 sg13g2_fill_2 FILLER_58_1012 ();
 sg13g2_fill_1 FILLER_58_1037 ();
 sg13g2_fill_2 FILLER_58_1051 ();
 sg13g2_fill_1 FILLER_58_1053 ();
 sg13g2_fill_1 FILLER_58_1067 ();
 sg13g2_decap_8 FILLER_58_1112 ();
 sg13g2_decap_8 FILLER_58_1119 ();
 sg13g2_fill_2 FILLER_58_1139 ();
 sg13g2_fill_2 FILLER_58_1204 ();
 sg13g2_fill_1 FILLER_58_1206 ();
 sg13g2_fill_2 FILLER_58_1216 ();
 sg13g2_fill_1 FILLER_58_1218 ();
 sg13g2_fill_2 FILLER_58_1224 ();
 sg13g2_fill_1 FILLER_58_1226 ();
 sg13g2_decap_8 FILLER_58_1281 ();
 sg13g2_decap_8 FILLER_58_1288 ();
 sg13g2_decap_8 FILLER_58_1295 ();
 sg13g2_decap_8 FILLER_58_1302 ();
 sg13g2_decap_4 FILLER_58_1309 ();
 sg13g2_fill_2 FILLER_58_1313 ();
 sg13g2_decap_8 FILLER_59_0 ();
 sg13g2_fill_1 FILLER_59_7 ();
 sg13g2_fill_1 FILLER_59_35 ();
 sg13g2_decap_8 FILLER_59_66 ();
 sg13g2_fill_1 FILLER_59_86 ();
 sg13g2_decap_4 FILLER_59_99 ();
 sg13g2_decap_8 FILLER_59_107 ();
 sg13g2_decap_4 FILLER_59_114 ();
 sg13g2_fill_1 FILLER_59_118 ();
 sg13g2_fill_2 FILLER_59_149 ();
 sg13g2_fill_1 FILLER_59_151 ();
 sg13g2_decap_4 FILLER_59_162 ();
 sg13g2_fill_1 FILLER_59_166 ();
 sg13g2_fill_2 FILLER_59_178 ();
 sg13g2_fill_2 FILLER_59_203 ();
 sg13g2_fill_1 FILLER_59_205 ();
 sg13g2_fill_1 FILLER_59_271 ();
 sg13g2_fill_2 FILLER_59_308 ();
 sg13g2_fill_1 FILLER_59_310 ();
 sg13g2_decap_4 FILLER_59_342 ();
 sg13g2_fill_1 FILLER_59_351 ();
 sg13g2_decap_4 FILLER_59_356 ();
 sg13g2_fill_1 FILLER_59_360 ();
 sg13g2_fill_1 FILLER_59_366 ();
 sg13g2_fill_2 FILLER_59_412 ();
 sg13g2_fill_1 FILLER_59_414 ();
 sg13g2_fill_2 FILLER_59_424 ();
 sg13g2_fill_1 FILLER_59_426 ();
 sg13g2_decap_4 FILLER_59_458 ();
 sg13g2_fill_1 FILLER_59_462 ();
 sg13g2_fill_2 FILLER_59_490 ();
 sg13g2_fill_1 FILLER_59_492 ();
 sg13g2_fill_2 FILLER_59_507 ();
 sg13g2_decap_8 FILLER_59_513 ();
 sg13g2_decap_8 FILLER_59_520 ();
 sg13g2_fill_1 FILLER_59_531 ();
 sg13g2_fill_1 FILLER_59_572 ();
 sg13g2_fill_2 FILLER_59_615 ();
 sg13g2_fill_2 FILLER_59_626 ();
 sg13g2_decap_8 FILLER_59_632 ();
 sg13g2_decap_8 FILLER_59_639 ();
 sg13g2_decap_8 FILLER_59_646 ();
 sg13g2_decap_4 FILLER_59_712 ();
 sg13g2_fill_1 FILLER_59_716 ();
 sg13g2_decap_8 FILLER_59_726 ();
 sg13g2_decap_8 FILLER_59_733 ();
 sg13g2_fill_2 FILLER_59_740 ();
 sg13g2_fill_1 FILLER_59_742 ();
 sg13g2_fill_2 FILLER_59_765 ();
 sg13g2_fill_1 FILLER_59_767 ();
 sg13g2_fill_2 FILLER_59_783 ();
 sg13g2_fill_2 FILLER_59_830 ();
 sg13g2_fill_2 FILLER_59_860 ();
 sg13g2_fill_2 FILLER_59_919 ();
 sg13g2_fill_2 FILLER_59_964 ();
 sg13g2_fill_1 FILLER_59_966 ();
 sg13g2_fill_2 FILLER_59_999 ();
 sg13g2_fill_2 FILLER_59_1032 ();
 sg13g2_fill_1 FILLER_59_1034 ();
 sg13g2_fill_2 FILLER_59_1095 ();
 sg13g2_fill_2 FILLER_59_1124 ();
 sg13g2_fill_1 FILLER_59_1153 ();
 sg13g2_fill_2 FILLER_59_1159 ();
 sg13g2_fill_1 FILLER_59_1161 ();
 sg13g2_fill_1 FILLER_59_1172 ();
 sg13g2_fill_1 FILLER_59_1187 ();
 sg13g2_fill_2 FILLER_59_1211 ();
 sg13g2_fill_1 FILLER_59_1213 ();
 sg13g2_fill_2 FILLER_59_1263 ();
 sg13g2_decap_8 FILLER_59_1287 ();
 sg13g2_decap_8 FILLER_59_1294 ();
 sg13g2_decap_8 FILLER_59_1301 ();
 sg13g2_decap_8 FILLER_59_1308 ();
 sg13g2_fill_2 FILLER_60_0 ();
 sg13g2_fill_1 FILLER_60_2 ();
 sg13g2_fill_2 FILLER_60_43 ();
 sg13g2_decap_8 FILLER_60_72 ();
 sg13g2_fill_1 FILLER_60_79 ();
 sg13g2_fill_1 FILLER_60_98 ();
 sg13g2_fill_2 FILLER_60_104 ();
 sg13g2_fill_1 FILLER_60_106 ();
 sg13g2_fill_1 FILLER_60_126 ();
 sg13g2_fill_2 FILLER_60_141 ();
 sg13g2_fill_2 FILLER_60_209 ();
 sg13g2_decap_8 FILLER_60_224 ();
 sg13g2_decap_8 FILLER_60_231 ();
 sg13g2_decap_8 FILLER_60_238 ();
 sg13g2_fill_2 FILLER_60_245 ();
 sg13g2_decap_4 FILLER_60_252 ();
 sg13g2_fill_2 FILLER_60_269 ();
 sg13g2_fill_1 FILLER_60_271 ();
 sg13g2_fill_2 FILLER_60_299 ();
 sg13g2_decap_8 FILLER_60_323 ();
 sg13g2_fill_2 FILLER_60_330 ();
 sg13g2_fill_1 FILLER_60_332 ();
 sg13g2_fill_2 FILLER_60_369 ();
 sg13g2_fill_2 FILLER_60_398 ();
 sg13g2_fill_1 FILLER_60_400 ();
 sg13g2_fill_1 FILLER_60_410 ();
 sg13g2_decap_4 FILLER_60_420 ();
 sg13g2_fill_2 FILLER_60_456 ();
 sg13g2_fill_1 FILLER_60_458 ();
 sg13g2_decap_8 FILLER_60_476 ();
 sg13g2_decap_8 FILLER_60_483 ();
 sg13g2_decap_4 FILLER_60_490 ();
 sg13g2_fill_2 FILLER_60_494 ();
 sg13g2_fill_1 FILLER_60_532 ();
 sg13g2_fill_2 FILLER_60_555 ();
 sg13g2_fill_1 FILLER_60_557 ();
 sg13g2_decap_8 FILLER_60_567 ();
 sg13g2_decap_4 FILLER_60_574 ();
 sg13g2_fill_2 FILLER_60_578 ();
 sg13g2_decap_8 FILLER_60_611 ();
 sg13g2_fill_1 FILLER_60_618 ();
 sg13g2_fill_1 FILLER_60_624 ();
 sg13g2_fill_2 FILLER_60_665 ();
 sg13g2_fill_2 FILLER_60_699 ();
 sg13g2_fill_1 FILLER_60_701 ();
 sg13g2_decap_4 FILLER_60_706 ();
 sg13g2_fill_2 FILLER_60_710 ();
 sg13g2_fill_2 FILLER_60_720 ();
 sg13g2_fill_1 FILLER_60_722 ();
 sg13g2_fill_1 FILLER_60_750 ();
 sg13g2_decap_8 FILLER_60_799 ();
 sg13g2_decap_8 FILLER_60_806 ();
 sg13g2_decap_8 FILLER_60_813 ();
 sg13g2_fill_1 FILLER_60_820 ();
 sg13g2_decap_8 FILLER_60_825 ();
 sg13g2_decap_4 FILLER_60_832 ();
 sg13g2_fill_1 FILLER_60_836 ();
 sg13g2_fill_2 FILLER_60_899 ();
 sg13g2_fill_1 FILLER_60_901 ();
 sg13g2_fill_2 FILLER_60_928 ();
 sg13g2_fill_1 FILLER_60_939 ();
 sg13g2_fill_2 FILLER_60_944 ();
 sg13g2_fill_1 FILLER_60_946 ();
 sg13g2_decap_8 FILLER_60_956 ();
 sg13g2_decap_8 FILLER_60_963 ();
 sg13g2_fill_2 FILLER_60_970 ();
 sg13g2_decap_8 FILLER_60_976 ();
 sg13g2_decap_8 FILLER_60_983 ();
 sg13g2_fill_2 FILLER_60_1027 ();
 sg13g2_fill_2 FILLER_60_1093 ();
 sg13g2_decap_8 FILLER_60_1108 ();
 sg13g2_fill_2 FILLER_60_1151 ();
 sg13g2_fill_1 FILLER_60_1153 ();
 sg13g2_fill_2 FILLER_60_1182 ();
 sg13g2_fill_2 FILLER_60_1210 ();
 sg13g2_fill_1 FILLER_60_1212 ();
 sg13g2_fill_2 FILLER_60_1251 ();
 sg13g2_fill_1 FILLER_60_1258 ();
 sg13g2_fill_1 FILLER_60_1267 ();
 sg13g2_decap_8 FILLER_60_1295 ();
 sg13g2_decap_8 FILLER_60_1302 ();
 sg13g2_decap_4 FILLER_60_1309 ();
 sg13g2_fill_2 FILLER_60_1313 ();
 sg13g2_fill_1 FILLER_61_23 ();
 sg13g2_decap_4 FILLER_61_70 ();
 sg13g2_fill_1 FILLER_61_74 ();
 sg13g2_fill_1 FILLER_61_112 ();
 sg13g2_fill_2 FILLER_61_146 ();
 sg13g2_fill_1 FILLER_61_148 ();
 sg13g2_decap_8 FILLER_61_162 ();
 sg13g2_fill_2 FILLER_61_169 ();
 sg13g2_fill_1 FILLER_61_171 ();
 sg13g2_decap_8 FILLER_61_203 ();
 sg13g2_decap_4 FILLER_61_210 ();
 sg13g2_fill_2 FILLER_61_214 ();
 sg13g2_decap_8 FILLER_61_220 ();
 sg13g2_decap_8 FILLER_61_227 ();
 sg13g2_decap_8 FILLER_61_234 ();
 sg13g2_fill_1 FILLER_61_241 ();
 sg13g2_fill_1 FILLER_61_292 ();
 sg13g2_fill_1 FILLER_61_337 ();
 sg13g2_fill_1 FILLER_61_365 ();
 sg13g2_fill_2 FILLER_61_371 ();
 sg13g2_fill_2 FILLER_61_459 ();
 sg13g2_fill_1 FILLER_61_461 ();
 sg13g2_fill_2 FILLER_61_489 ();
 sg13g2_fill_1 FILLER_61_500 ();
 sg13g2_fill_2 FILLER_61_505 ();
 sg13g2_fill_1 FILLER_61_507 ();
 sg13g2_fill_2 FILLER_61_513 ();
 sg13g2_decap_8 FILLER_61_560 ();
 sg13g2_decap_8 FILLER_61_567 ();
 sg13g2_decap_4 FILLER_61_574 ();
 sg13g2_fill_1 FILLER_61_578 ();
 sg13g2_fill_2 FILLER_61_601 ();
 sg13g2_fill_1 FILLER_61_603 ();
 sg13g2_fill_2 FILLER_61_617 ();
 sg13g2_fill_1 FILLER_61_619 ();
 sg13g2_fill_2 FILLER_61_670 ();
 sg13g2_fill_1 FILLER_61_676 ();
 sg13g2_fill_1 FILLER_61_681 ();
 sg13g2_decap_8 FILLER_61_695 ();
 sg13g2_decap_8 FILLER_61_702 ();
 sg13g2_decap_8 FILLER_61_709 ();
 sg13g2_fill_2 FILLER_61_716 ();
 sg13g2_fill_1 FILLER_61_718 ();
 sg13g2_fill_1 FILLER_61_760 ();
 sg13g2_decap_8 FILLER_61_788 ();
 sg13g2_decap_8 FILLER_61_795 ();
 sg13g2_decap_4 FILLER_61_802 ();
 sg13g2_decap_8 FILLER_61_814 ();
 sg13g2_decap_4 FILLER_61_821 ();
 sg13g2_fill_1 FILLER_61_825 ();
 sg13g2_decap_8 FILLER_61_831 ();
 sg13g2_fill_1 FILLER_61_838 ();
 sg13g2_fill_2 FILLER_61_875 ();
 sg13g2_fill_1 FILLER_61_877 ();
 sg13g2_decap_4 FILLER_61_927 ();
 sg13g2_fill_1 FILLER_61_931 ();
 sg13g2_fill_2 FILLER_61_941 ();
 sg13g2_decap_4 FILLER_61_987 ();
 sg13g2_fill_1 FILLER_61_1012 ();
 sg13g2_fill_2 FILLER_61_1035 ();
 sg13g2_fill_2 FILLER_61_1042 ();
 sg13g2_fill_1 FILLER_61_1071 ();
 sg13g2_fill_2 FILLER_61_1087 ();
 sg13g2_fill_1 FILLER_61_1089 ();
 sg13g2_fill_2 FILLER_61_1099 ();
 sg13g2_fill_1 FILLER_61_1101 ();
 sg13g2_decap_8 FILLER_61_1115 ();
 sg13g2_fill_2 FILLER_61_1122 ();
 sg13g2_fill_1 FILLER_61_1146 ();
 sg13g2_fill_1 FILLER_61_1172 ();
 sg13g2_decap_4 FILLER_61_1210 ();
 sg13g2_fill_2 FILLER_61_1214 ();
 sg13g2_fill_2 FILLER_61_1255 ();
 sg13g2_fill_1 FILLER_61_1257 ();
 sg13g2_decap_8 FILLER_61_1262 ();
 sg13g2_decap_8 FILLER_61_1269 ();
 sg13g2_fill_2 FILLER_61_1276 ();
 sg13g2_decap_8 FILLER_61_1287 ();
 sg13g2_decap_8 FILLER_61_1294 ();
 sg13g2_decap_8 FILLER_61_1301 ();
 sg13g2_decap_8 FILLER_61_1308 ();
 sg13g2_decap_4 FILLER_62_0 ();
 sg13g2_fill_2 FILLER_62_48 ();
 sg13g2_fill_2 FILLER_62_73 ();
 sg13g2_fill_1 FILLER_62_130 ();
 sg13g2_fill_2 FILLER_62_140 ();
 sg13g2_fill_1 FILLER_62_142 ();
 sg13g2_decap_8 FILLER_62_157 ();
 sg13g2_decap_4 FILLER_62_164 ();
 sg13g2_fill_2 FILLER_62_168 ();
 sg13g2_decap_4 FILLER_62_174 ();
 sg13g2_fill_2 FILLER_62_178 ();
 sg13g2_fill_2 FILLER_62_184 ();
 sg13g2_decap_8 FILLER_62_202 ();
 sg13g2_fill_1 FILLER_62_209 ();
 sg13g2_fill_1 FILLER_62_238 ();
 sg13g2_decap_4 FILLER_62_257 ();
 sg13g2_fill_2 FILLER_62_261 ();
 sg13g2_fill_2 FILLER_62_290 ();
 sg13g2_fill_1 FILLER_62_292 ();
 sg13g2_fill_2 FILLER_62_320 ();
 sg13g2_fill_1 FILLER_62_322 ();
 sg13g2_fill_1 FILLER_62_386 ();
 sg13g2_fill_2 FILLER_62_409 ();
 sg13g2_fill_1 FILLER_62_411 ();
 sg13g2_fill_1 FILLER_62_438 ();
 sg13g2_decap_4 FILLER_62_458 ();
 sg13g2_fill_2 FILLER_62_475 ();
 sg13g2_fill_1 FILLER_62_477 ();
 sg13g2_fill_1 FILLER_62_536 ();
 sg13g2_fill_2 FILLER_62_541 ();
 sg13g2_fill_1 FILLER_62_543 ();
 sg13g2_fill_1 FILLER_62_576 ();
 sg13g2_decap_4 FILLER_62_581 ();
 sg13g2_fill_1 FILLER_62_585 ();
 sg13g2_fill_1 FILLER_62_612 ();
 sg13g2_fill_2 FILLER_62_640 ();
 sg13g2_decap_8 FILLER_62_670 ();
 sg13g2_decap_8 FILLER_62_677 ();
 sg13g2_decap_8 FILLER_62_684 ();
 sg13g2_decap_8 FILLER_62_691 ();
 sg13g2_decap_8 FILLER_62_698 ();
 sg13g2_decap_8 FILLER_62_705 ();
 sg13g2_decap_8 FILLER_62_712 ();
 sg13g2_fill_2 FILLER_62_719 ();
 sg13g2_fill_2 FILLER_62_743 ();
 sg13g2_fill_1 FILLER_62_745 ();
 sg13g2_fill_1 FILLER_62_755 ();
 sg13g2_fill_1 FILLER_62_761 ();
 sg13g2_fill_2 FILLER_62_848 ();
 sg13g2_fill_1 FILLER_62_850 ();
 sg13g2_decap_4 FILLER_62_870 ();
 sg13g2_fill_1 FILLER_62_878 ();
 sg13g2_fill_1 FILLER_62_896 ();
 sg13g2_fill_2 FILLER_62_946 ();
 sg13g2_fill_2 FILLER_62_980 ();
 sg13g2_decap_8 FILLER_62_991 ();
 sg13g2_decap_8 FILLER_62_998 ();
 sg13g2_fill_2 FILLER_62_1009 ();
 sg13g2_decap_8 FILLER_62_1015 ();
 sg13g2_decap_8 FILLER_62_1022 ();
 sg13g2_decap_4 FILLER_62_1029 ();
 sg13g2_decap_4 FILLER_62_1037 ();
 sg13g2_fill_1 FILLER_62_1041 ();
 sg13g2_decap_8 FILLER_62_1054 ();
 sg13g2_fill_1 FILLER_62_1069 ();
 sg13g2_decap_8 FILLER_62_1090 ();
 sg13g2_fill_2 FILLER_62_1097 ();
 sg13g2_fill_1 FILLER_62_1099 ();
 sg13g2_decap_4 FILLER_62_1144 ();
 sg13g2_fill_2 FILLER_62_1161 ();
 sg13g2_fill_1 FILLER_62_1163 ();
 sg13g2_fill_2 FILLER_62_1204 ();
 sg13g2_decap_8 FILLER_62_1219 ();
 sg13g2_fill_1 FILLER_62_1238 ();
 sg13g2_decap_8 FILLER_62_1258 ();
 sg13g2_decap_8 FILLER_62_1265 ();
 sg13g2_decap_8 FILLER_62_1272 ();
 sg13g2_decap_8 FILLER_62_1279 ();
 sg13g2_decap_8 FILLER_62_1286 ();
 sg13g2_decap_8 FILLER_62_1293 ();
 sg13g2_decap_8 FILLER_62_1300 ();
 sg13g2_decap_8 FILLER_62_1307 ();
 sg13g2_fill_1 FILLER_62_1314 ();
 sg13g2_fill_2 FILLER_63_39 ();
 sg13g2_fill_2 FILLER_63_55 ();
 sg13g2_fill_1 FILLER_63_57 ();
 sg13g2_fill_1 FILLER_63_71 ();
 sg13g2_fill_1 FILLER_63_99 ();
 sg13g2_fill_1 FILLER_63_147 ();
 sg13g2_decap_8 FILLER_63_162 ();
 sg13g2_decap_8 FILLER_63_173 ();
 sg13g2_decap_4 FILLER_63_180 ();
 sg13g2_fill_1 FILLER_63_184 ();
 sg13g2_fill_2 FILLER_63_198 ();
 sg13g2_fill_1 FILLER_63_200 ();
 sg13g2_fill_2 FILLER_63_214 ();
 sg13g2_decap_8 FILLER_63_249 ();
 sg13g2_decap_8 FILLER_63_256 ();
 sg13g2_fill_1 FILLER_63_263 ();
 sg13g2_fill_1 FILLER_63_272 ();
 sg13g2_fill_1 FILLER_63_283 ();
 sg13g2_fill_2 FILLER_63_303 ();
 sg13g2_fill_1 FILLER_63_305 ();
 sg13g2_fill_1 FILLER_63_356 ();
 sg13g2_fill_2 FILLER_63_366 ();
 sg13g2_decap_4 FILLER_63_423 ();
 sg13g2_fill_2 FILLER_63_427 ();
 sg13g2_decap_8 FILLER_63_442 ();
 sg13g2_decap_8 FILLER_63_449 ();
 sg13g2_fill_2 FILLER_63_499 ();
 sg13g2_fill_1 FILLER_63_501 ();
 sg13g2_fill_2 FILLER_63_520 ();
 sg13g2_fill_1 FILLER_63_522 ();
 sg13g2_decap_8 FILLER_63_537 ();
 sg13g2_decap_4 FILLER_63_544 ();
 sg13g2_fill_1 FILLER_63_611 ();
 sg13g2_fill_2 FILLER_63_652 ();
 sg13g2_fill_1 FILLER_63_654 ();
 sg13g2_fill_2 FILLER_63_667 ();
 sg13g2_fill_1 FILLER_63_669 ();
 sg13g2_fill_2 FILLER_63_675 ();
 sg13g2_decap_8 FILLER_63_704 ();
 sg13g2_decap_8 FILLER_63_715 ();
 sg13g2_decap_4 FILLER_63_722 ();
 sg13g2_fill_2 FILLER_63_726 ();
 sg13g2_decap_4 FILLER_63_732 ();
 sg13g2_fill_1 FILLER_63_736 ();
 sg13g2_fill_1 FILLER_63_754 ();
 sg13g2_fill_2 FILLER_63_787 ();
 sg13g2_fill_1 FILLER_63_789 ();
 sg13g2_fill_2 FILLER_63_867 ();
 sg13g2_fill_1 FILLER_63_869 ();
 sg13g2_fill_2 FILLER_63_919 ();
 sg13g2_fill_1 FILLER_63_921 ();
 sg13g2_fill_2 FILLER_63_949 ();
 sg13g2_fill_1 FILLER_63_951 ();
 sg13g2_fill_1 FILLER_63_974 ();
 sg13g2_fill_2 FILLER_63_993 ();
 sg13g2_decap_4 FILLER_63_1008 ();
 sg13g2_decap_4 FILLER_63_1017 ();
 sg13g2_fill_1 FILLER_63_1021 ();
 sg13g2_decap_8 FILLER_63_1026 ();
 sg13g2_fill_1 FILLER_63_1033 ();
 sg13g2_decap_8 FILLER_63_1039 ();
 sg13g2_decap_8 FILLER_63_1046 ();
 sg13g2_decap_4 FILLER_63_1053 ();
 sg13g2_decap_8 FILLER_63_1066 ();
 sg13g2_decap_8 FILLER_63_1077 ();
 sg13g2_fill_2 FILLER_63_1084 ();
 sg13g2_fill_1 FILLER_63_1086 ();
 sg13g2_decap_4 FILLER_63_1149 ();
 sg13g2_fill_1 FILLER_63_1170 ();
 sg13g2_fill_2 FILLER_63_1184 ();
 sg13g2_fill_1 FILLER_63_1186 ();
 sg13g2_fill_1 FILLER_63_1232 ();
 sg13g2_decap_8 FILLER_63_1274 ();
 sg13g2_decap_8 FILLER_63_1281 ();
 sg13g2_decap_8 FILLER_63_1288 ();
 sg13g2_decap_8 FILLER_63_1295 ();
 sg13g2_decap_8 FILLER_63_1302 ();
 sg13g2_decap_4 FILLER_63_1309 ();
 sg13g2_fill_2 FILLER_63_1313 ();
 sg13g2_fill_2 FILLER_64_0 ();
 sg13g2_fill_1 FILLER_64_2 ();
 sg13g2_fill_1 FILLER_64_36 ();
 sg13g2_fill_2 FILLER_64_52 ();
 sg13g2_decap_8 FILLER_64_67 ();
 sg13g2_fill_2 FILLER_64_120 ();
 sg13g2_fill_1 FILLER_64_122 ();
 sg13g2_fill_1 FILLER_64_129 ();
 sg13g2_fill_2 FILLER_64_163 ();
 sg13g2_decap_8 FILLER_64_178 ();
 sg13g2_decap_4 FILLER_64_185 ();
 sg13g2_fill_1 FILLER_64_189 ();
 sg13g2_decap_8 FILLER_64_259 ();
 sg13g2_decap_8 FILLER_64_266 ();
 sg13g2_decap_8 FILLER_64_273 ();
 sg13g2_decap_4 FILLER_64_280 ();
 sg13g2_fill_1 FILLER_64_306 ();
 sg13g2_decap_8 FILLER_64_317 ();
 sg13g2_fill_1 FILLER_64_324 ();
 sg13g2_fill_1 FILLER_64_329 ();
 sg13g2_fill_1 FILLER_64_334 ();
 sg13g2_fill_2 FILLER_64_340 ();
 sg13g2_fill_2 FILLER_64_378 ();
 sg13g2_fill_2 FILLER_64_385 ();
 sg13g2_fill_1 FILLER_64_387 ();
 sg13g2_decap_4 FILLER_64_392 ();
 sg13g2_decap_4 FILLER_64_424 ();
 sg13g2_decap_4 FILLER_64_436 ();
 sg13g2_decap_8 FILLER_64_459 ();
 sg13g2_fill_1 FILLER_64_466 ();
 sg13g2_fill_2 FILLER_64_483 ();
 sg13g2_decap_8 FILLER_64_489 ();
 sg13g2_fill_2 FILLER_64_505 ();
 sg13g2_decap_4 FILLER_64_542 ();
 sg13g2_fill_1 FILLER_64_546 ();
 sg13g2_decap_4 FILLER_64_569 ();
 sg13g2_fill_2 FILLER_64_605 ();
 sg13g2_fill_1 FILLER_64_607 ();
 sg13g2_fill_1 FILLER_64_645 ();
 sg13g2_decap_8 FILLER_64_652 ();
 sg13g2_decap_4 FILLER_64_659 ();
 sg13g2_fill_1 FILLER_64_668 ();
 sg13g2_decap_4 FILLER_64_700 ();
 sg13g2_fill_2 FILLER_64_704 ();
 sg13g2_fill_2 FILLER_64_734 ();
 sg13g2_fill_1 FILLER_64_736 ();
 sg13g2_fill_1 FILLER_64_750 ();
 sg13g2_fill_1 FILLER_64_755 ();
 sg13g2_fill_2 FILLER_64_783 ();
 sg13g2_fill_2 FILLER_64_808 ();
 sg13g2_fill_2 FILLER_64_837 ();
 sg13g2_fill_1 FILLER_64_890 ();
 sg13g2_fill_2 FILLER_64_915 ();
 sg13g2_fill_1 FILLER_64_954 ();
 sg13g2_decap_4 FILLER_64_1077 ();
 sg13g2_fill_1 FILLER_64_1081 ();
 sg13g2_decap_8 FILLER_64_1168 ();
 sg13g2_decap_4 FILLER_64_1188 ();
 sg13g2_fill_2 FILLER_64_1228 ();
 sg13g2_fill_1 FILLER_64_1230 ();
 sg13g2_decap_8 FILLER_64_1290 ();
 sg13g2_decap_8 FILLER_64_1297 ();
 sg13g2_decap_8 FILLER_64_1304 ();
 sg13g2_decap_4 FILLER_64_1311 ();
 sg13g2_fill_2 FILLER_65_0 ();
 sg13g2_fill_2 FILLER_65_45 ();
 sg13g2_fill_1 FILLER_65_47 ();
 sg13g2_decap_4 FILLER_65_62 ();
 sg13g2_fill_1 FILLER_65_128 ();
 sg13g2_fill_1 FILLER_65_172 ();
 sg13g2_fill_1 FILLER_65_237 ();
 sg13g2_decap_4 FILLER_65_263 ();
 sg13g2_fill_2 FILLER_65_271 ();
 sg13g2_fill_1 FILLER_65_273 ();
 sg13g2_fill_2 FILLER_65_279 ();
 sg13g2_decap_4 FILLER_65_285 ();
 sg13g2_decap_4 FILLER_65_293 ();
 sg13g2_fill_1 FILLER_65_297 ();
 sg13g2_fill_1 FILLER_65_302 ();
 sg13g2_decap_8 FILLER_65_320 ();
 sg13g2_decap_8 FILLER_65_327 ();
 sg13g2_decap_8 FILLER_65_334 ();
 sg13g2_fill_2 FILLER_65_367 ();
 sg13g2_fill_1 FILLER_65_373 ();
 sg13g2_decap_8 FILLER_65_410 ();
 sg13g2_decap_4 FILLER_65_417 ();
 sg13g2_fill_1 FILLER_65_421 ();
 sg13g2_fill_1 FILLER_65_459 ();
 sg13g2_decap_8 FILLER_65_469 ();
 sg13g2_fill_2 FILLER_65_516 ();
 sg13g2_fill_1 FILLER_65_518 ();
 sg13g2_fill_2 FILLER_65_528 ();
 sg13g2_fill_1 FILLER_65_530 ();
 sg13g2_decap_4 FILLER_65_558 ();
 sg13g2_fill_2 FILLER_65_562 ();
 sg13g2_decap_8 FILLER_65_604 ();
 sg13g2_fill_2 FILLER_65_611 ();
 sg13g2_decap_8 FILLER_65_656 ();
 sg13g2_fill_2 FILLER_65_663 ();
 sg13g2_fill_1 FILLER_65_665 ();
 sg13g2_decap_8 FILLER_65_710 ();
 sg13g2_decap_8 FILLER_65_717 ();
 sg13g2_decap_8 FILLER_65_724 ();
 sg13g2_decap_8 FILLER_65_731 ();
 sg13g2_decap_8 FILLER_65_738 ();
 sg13g2_fill_2 FILLER_65_757 ();
 sg13g2_fill_1 FILLER_65_759 ();
 sg13g2_fill_1 FILLER_65_779 ();
 sg13g2_fill_1 FILLER_65_793 ();
 sg13g2_fill_1 FILLER_65_806 ();
 sg13g2_fill_2 FILLER_65_939 ();
 sg13g2_fill_1 FILLER_65_941 ();
 sg13g2_fill_1 FILLER_65_964 ();
 sg13g2_fill_2 FILLER_65_1125 ();
 sg13g2_fill_2 FILLER_65_1167 ();
 sg13g2_fill_1 FILLER_65_1169 ();
 sg13g2_fill_2 FILLER_65_1197 ();
 sg13g2_fill_1 FILLER_65_1199 ();
 sg13g2_decap_8 FILLER_65_1224 ();
 sg13g2_fill_2 FILLER_65_1231 ();
 sg13g2_fill_1 FILLER_65_1233 ();
 sg13g2_fill_1 FILLER_65_1243 ();
 sg13g2_fill_2 FILLER_65_1250 ();
 sg13g2_fill_2 FILLER_65_1276 ();
 sg13g2_fill_1 FILLER_65_1278 ();
 sg13g2_decap_8 FILLER_65_1288 ();
 sg13g2_decap_8 FILLER_65_1295 ();
 sg13g2_decap_8 FILLER_65_1302 ();
 sg13g2_decap_4 FILLER_65_1309 ();
 sg13g2_fill_2 FILLER_65_1313 ();
 sg13g2_decap_8 FILLER_66_0 ();
 sg13g2_fill_1 FILLER_66_7 ();
 sg13g2_fill_1 FILLER_66_124 ();
 sg13g2_fill_1 FILLER_66_161 ();
 sg13g2_fill_2 FILLER_66_176 ();
 sg13g2_decap_4 FILLER_66_258 ();
 sg13g2_fill_2 FILLER_66_307 ();
 sg13g2_fill_1 FILLER_66_309 ();
 sg13g2_fill_2 FILLER_66_315 ();
 sg13g2_fill_1 FILLER_66_323 ();
 sg13g2_fill_2 FILLER_66_360 ();
 sg13g2_fill_2 FILLER_66_367 ();
 sg13g2_fill_1 FILLER_66_369 ();
 sg13g2_fill_2 FILLER_66_407 ();
 sg13g2_fill_1 FILLER_66_409 ();
 sg13g2_fill_1 FILLER_66_527 ();
 sg13g2_fill_2 FILLER_66_560 ();
 sg13g2_fill_1 FILLER_66_562 ();
 sg13g2_fill_1 FILLER_66_596 ();
 sg13g2_fill_2 FILLER_66_612 ();
 sg13g2_fill_1 FILLER_66_627 ();
 sg13g2_fill_1 FILLER_66_669 ();
 sg13g2_fill_1 FILLER_66_750 ();
 sg13g2_fill_2 FILLER_66_841 ();
 sg13g2_fill_1 FILLER_66_883 ();
 sg13g2_fill_1 FILLER_66_895 ();
 sg13g2_fill_1 FILLER_66_932 ();
 sg13g2_fill_2 FILLER_66_938 ();
 sg13g2_fill_1 FILLER_66_940 ();
 sg13g2_fill_2 FILLER_66_973 ();
 sg13g2_fill_1 FILLER_66_975 ();
 sg13g2_fill_1 FILLER_66_989 ();
 sg13g2_fill_2 FILLER_66_1028 ();
 sg13g2_fill_1 FILLER_66_1102 ();
 sg13g2_decap_4 FILLER_66_1150 ();
 sg13g2_fill_2 FILLER_66_1202 ();
 sg13g2_decap_8 FILLER_66_1231 ();
 sg13g2_fill_2 FILLER_66_1238 ();
 sg13g2_fill_1 FILLER_66_1244 ();
 sg13g2_decap_8 FILLER_66_1281 ();
 sg13g2_decap_8 FILLER_66_1288 ();
 sg13g2_decap_8 FILLER_66_1295 ();
 sg13g2_decap_8 FILLER_66_1302 ();
 sg13g2_decap_4 FILLER_66_1309 ();
 sg13g2_fill_2 FILLER_66_1313 ();
 sg13g2_fill_1 FILLER_67_0 ();
 sg13g2_decap_4 FILLER_67_61 ();
 sg13g2_fill_2 FILLER_67_65 ();
 sg13g2_fill_2 FILLER_67_93 ();
 sg13g2_fill_1 FILLER_67_95 ();
 sg13g2_fill_2 FILLER_67_110 ();
 sg13g2_fill_1 FILLER_67_134 ();
 sg13g2_fill_2 FILLER_67_204 ();
 sg13g2_decap_4 FILLER_67_259 ();
 sg13g2_fill_2 FILLER_67_301 ();
 sg13g2_fill_1 FILLER_67_331 ();
 sg13g2_fill_2 FILLER_67_382 ();
 sg13g2_fill_1 FILLER_67_426 ();
 sg13g2_fill_2 FILLER_67_454 ();
 sg13g2_fill_1 FILLER_67_456 ();
 sg13g2_fill_2 FILLER_67_472 ();
 sg13g2_fill_1 FILLER_67_519 ();
 sg13g2_decap_4 FILLER_67_551 ();
 sg13g2_fill_1 FILLER_67_564 ();
 sg13g2_fill_1 FILLER_67_592 ();
 sg13g2_fill_1 FILLER_67_599 ();
 sg13g2_decap_4 FILLER_67_650 ();
 sg13g2_fill_2 FILLER_67_654 ();
 sg13g2_decap_4 FILLER_67_665 ();
 sg13g2_decap_4 FILLER_67_713 ();
 sg13g2_fill_2 FILLER_67_717 ();
 sg13g2_fill_2 FILLER_67_755 ();
 sg13g2_fill_1 FILLER_67_757 ();
 sg13g2_fill_1 FILLER_67_785 ();
 sg13g2_fill_2 FILLER_67_822 ();
 sg13g2_fill_1 FILLER_67_858 ();
 sg13g2_decap_8 FILLER_67_872 ();
 sg13g2_fill_1 FILLER_67_879 ();
 sg13g2_decap_8 FILLER_67_889 ();
 sg13g2_decap_8 FILLER_67_896 ();
 sg13g2_fill_1 FILLER_67_903 ();
 sg13g2_fill_2 FILLER_67_908 ();
 sg13g2_fill_1 FILLER_67_910 ();
 sg13g2_fill_1 FILLER_67_919 ();
 sg13g2_fill_2 FILLER_67_926 ();
 sg13g2_fill_1 FILLER_67_933 ();
 sg13g2_decap_8 FILLER_67_970 ();
 sg13g2_decap_4 FILLER_67_977 ();
 sg13g2_fill_1 FILLER_67_1007 ();
 sg13g2_fill_2 FILLER_67_1030 ();
 sg13g2_fill_1 FILLER_67_1032 ();
 sg13g2_fill_2 FILLER_67_1062 ();
 sg13g2_fill_1 FILLER_67_1064 ();
 sg13g2_fill_2 FILLER_67_1091 ();
 sg13g2_fill_1 FILLER_67_1093 ();
 sg13g2_fill_1 FILLER_67_1115 ();
 sg13g2_fill_1 FILLER_67_1130 ();
 sg13g2_decap_8 FILLER_67_1145 ();
 sg13g2_decap_4 FILLER_67_1152 ();
 sg13g2_fill_1 FILLER_67_1156 ();
 sg13g2_fill_2 FILLER_67_1199 ();
 sg13g2_fill_1 FILLER_67_1201 ();
 sg13g2_fill_2 FILLER_67_1245 ();
 sg13g2_decap_8 FILLER_67_1277 ();
 sg13g2_decap_8 FILLER_67_1284 ();
 sg13g2_decap_8 FILLER_67_1291 ();
 sg13g2_decap_8 FILLER_67_1298 ();
 sg13g2_decap_8 FILLER_67_1305 ();
 sg13g2_fill_2 FILLER_67_1312 ();
 sg13g2_fill_1 FILLER_67_1314 ();
 sg13g2_decap_4 FILLER_68_0 ();
 sg13g2_fill_2 FILLER_68_4 ();
 sg13g2_decap_4 FILLER_68_69 ();
 sg13g2_fill_2 FILLER_68_73 ();
 sg13g2_fill_2 FILLER_68_88 ();
 sg13g2_fill_1 FILLER_68_90 ();
 sg13g2_decap_4 FILLER_68_113 ();
 sg13g2_fill_2 FILLER_68_137 ();
 sg13g2_decap_4 FILLER_68_181 ();
 sg13g2_fill_1 FILLER_68_198 ();
 sg13g2_decap_4 FILLER_68_254 ();
 sg13g2_fill_1 FILLER_68_258 ();
 sg13g2_fill_2 FILLER_68_358 ();
 sg13g2_fill_1 FILLER_68_360 ();
 sg13g2_fill_1 FILLER_68_402 ();
 sg13g2_fill_1 FILLER_68_409 ();
 sg13g2_fill_2 FILLER_68_428 ();
 sg13g2_fill_1 FILLER_68_430 ();
 sg13g2_decap_4 FILLER_68_467 ();
 sg13g2_fill_2 FILLER_68_508 ();
 sg13g2_fill_1 FILLER_68_510 ();
 sg13g2_fill_2 FILLER_68_528 ();
 sg13g2_fill_1 FILLER_68_530 ();
 sg13g2_decap_8 FILLER_68_553 ();
 sg13g2_fill_1 FILLER_68_560 ();
 sg13g2_decap_4 FILLER_68_565 ();
 sg13g2_fill_1 FILLER_68_569 ();
 sg13g2_decap_8 FILLER_68_594 ();
 sg13g2_decap_4 FILLER_68_601 ();
 sg13g2_fill_2 FILLER_68_605 ();
 sg13g2_fill_1 FILLER_68_664 ();
 sg13g2_decap_8 FILLER_68_692 ();
 sg13g2_decap_8 FILLER_68_699 ();
 sg13g2_fill_2 FILLER_68_719 ();
 sg13g2_decap_4 FILLER_68_775 ();
 sg13g2_fill_1 FILLER_68_853 ();
 sg13g2_fill_2 FILLER_68_867 ();
 sg13g2_fill_1 FILLER_68_869 ();
 sg13g2_decap_4 FILLER_68_879 ();
 sg13g2_fill_1 FILLER_68_883 ();
 sg13g2_decap_8 FILLER_68_888 ();
 sg13g2_decap_4 FILLER_68_895 ();
 sg13g2_fill_2 FILLER_68_899 ();
 sg13g2_fill_2 FILLER_68_905 ();
 sg13g2_fill_2 FILLER_68_911 ();
 sg13g2_fill_1 FILLER_68_913 ();
 sg13g2_fill_2 FILLER_68_924 ();
 sg13g2_fill_1 FILLER_68_926 ();
 sg13g2_fill_1 FILLER_68_933 ();
 sg13g2_fill_1 FILLER_68_942 ();
 sg13g2_fill_2 FILLER_68_956 ();
 sg13g2_decap_8 FILLER_68_963 ();
 sg13g2_decap_8 FILLER_68_970 ();
 sg13g2_fill_2 FILLER_68_977 ();
 sg13g2_fill_1 FILLER_68_979 ();
 sg13g2_fill_1 FILLER_68_985 ();
 sg13g2_fill_2 FILLER_68_1008 ();
 sg13g2_fill_1 FILLER_68_1023 ();
 sg13g2_fill_1 FILLER_68_1063 ();
 sg13g2_decap_4 FILLER_68_1091 ();
 sg13g2_fill_1 FILLER_68_1095 ();
 sg13g2_fill_1 FILLER_68_1105 ();
 sg13g2_fill_2 FILLER_68_1115 ();
 sg13g2_fill_1 FILLER_68_1117 ();
 sg13g2_decap_4 FILLER_68_1145 ();
 sg13g2_fill_1 FILLER_68_1149 ();
 sg13g2_fill_2 FILLER_68_1190 ();
 sg13g2_fill_1 FILLER_68_1196 ();
 sg13g2_fill_1 FILLER_68_1210 ();
 sg13g2_fill_2 FILLER_68_1242 ();
 sg13g2_fill_1 FILLER_68_1250 ();
 sg13g2_fill_2 FILLER_68_1273 ();
 sg13g2_decap_8 FILLER_68_1284 ();
 sg13g2_decap_8 FILLER_68_1291 ();
 sg13g2_decap_8 FILLER_68_1298 ();
 sg13g2_decap_8 FILLER_68_1305 ();
 sg13g2_fill_2 FILLER_68_1312 ();
 sg13g2_fill_1 FILLER_68_1314 ();
 sg13g2_fill_2 FILLER_69_0 ();
 sg13g2_decap_4 FILLER_69_53 ();
 sg13g2_fill_1 FILLER_69_57 ();
 sg13g2_fill_2 FILLER_69_62 ();
 sg13g2_fill_1 FILLER_69_64 ();
 sg13g2_decap_8 FILLER_69_75 ();
 sg13g2_decap_4 FILLER_69_82 ();
 sg13g2_fill_1 FILLER_69_86 ();
 sg13g2_decap_8 FILLER_69_115 ();
 sg13g2_decap_8 FILLER_69_122 ();
 sg13g2_fill_2 FILLER_69_129 ();
 sg13g2_decap_4 FILLER_69_140 ();
 sg13g2_fill_1 FILLER_69_189 ();
 sg13g2_fill_2 FILLER_69_203 ();
 sg13g2_fill_1 FILLER_69_205 ();
 sg13g2_decap_4 FILLER_69_254 ();
 sg13g2_fill_2 FILLER_69_308 ();
 sg13g2_decap_8 FILLER_69_316 ();
 sg13g2_decap_8 FILLER_69_323 ();
 sg13g2_fill_2 FILLER_69_330 ();
 sg13g2_decap_8 FILLER_69_336 ();
 sg13g2_decap_4 FILLER_69_343 ();
 sg13g2_fill_2 FILLER_69_347 ();
 sg13g2_fill_1 FILLER_69_354 ();
 sg13g2_fill_2 FILLER_69_372 ();
 sg13g2_fill_1 FILLER_69_374 ();
 sg13g2_decap_8 FILLER_69_379 ();
 sg13g2_decap_4 FILLER_69_386 ();
 sg13g2_fill_2 FILLER_69_390 ();
 sg13g2_decap_8 FILLER_69_396 ();
 sg13g2_decap_8 FILLER_69_403 ();
 sg13g2_fill_1 FILLER_69_410 ();
 sg13g2_decap_8 FILLER_69_415 ();
 sg13g2_fill_2 FILLER_69_422 ();
 sg13g2_fill_1 FILLER_69_437 ();
 sg13g2_decap_8 FILLER_69_461 ();
 sg13g2_decap_4 FILLER_69_468 ();
 sg13g2_fill_1 FILLER_69_472 ();
 sg13g2_fill_1 FILLER_69_483 ();
 sg13g2_fill_2 FILLER_69_512 ();
 sg13g2_fill_2 FILLER_69_541 ();
 sg13g2_fill_1 FILLER_69_552 ();
 sg13g2_fill_2 FILLER_69_564 ();
 sg13g2_fill_2 FILLER_69_593 ();
 sg13g2_fill_1 FILLER_69_595 ();
 sg13g2_fill_2 FILLER_69_618 ();
 sg13g2_decap_8 FILLER_69_651 ();
 sg13g2_decap_4 FILLER_69_658 ();
 sg13g2_fill_2 FILLER_69_662 ();
 sg13g2_fill_2 FILLER_69_677 ();
 sg13g2_fill_1 FILLER_69_685 ();
 sg13g2_decap_8 FILLER_69_700 ();
 sg13g2_decap_8 FILLER_69_707 ();
 sg13g2_fill_2 FILLER_69_714 ();
 sg13g2_decap_4 FILLER_69_721 ();
 sg13g2_fill_1 FILLER_69_785 ();
 sg13g2_fill_2 FILLER_69_795 ();
 sg13g2_fill_2 FILLER_69_907 ();
 sg13g2_decap_4 FILLER_69_968 ();
 sg13g2_decap_4 FILLER_69_1045 ();
 sg13g2_decap_4 FILLER_69_1097 ();
 sg13g2_decap_4 FILLER_69_1141 ();
 sg13g2_fill_2 FILLER_69_1190 ();
 sg13g2_fill_1 FILLER_69_1192 ();
 sg13g2_fill_1 FILLER_69_1206 ();
 sg13g2_fill_1 FILLER_69_1236 ();
 sg13g2_decap_8 FILLER_69_1291 ();
 sg13g2_decap_8 FILLER_69_1298 ();
 sg13g2_decap_8 FILLER_69_1305 ();
 sg13g2_fill_2 FILLER_69_1312 ();
 sg13g2_fill_1 FILLER_69_1314 ();
 sg13g2_decap_8 FILLER_70_0 ();
 sg13g2_fill_1 FILLER_70_7 ();
 sg13g2_fill_1 FILLER_70_35 ();
 sg13g2_decap_8 FILLER_70_53 ();
 sg13g2_fill_2 FILLER_70_110 ();
 sg13g2_fill_2 FILLER_70_121 ();
 sg13g2_fill_2 FILLER_70_127 ();
 sg13g2_decap_4 FILLER_70_135 ();
 sg13g2_fill_2 FILLER_70_145 ();
 sg13g2_fill_1 FILLER_70_147 ();
 sg13g2_fill_2 FILLER_70_152 ();
 sg13g2_fill_2 FILLER_70_167 ();
 sg13g2_decap_4 FILLER_70_178 ();
 sg13g2_fill_1 FILLER_70_182 ();
 sg13g2_fill_1 FILLER_70_233 ();
 sg13g2_fill_2 FILLER_70_239 ();
 sg13g2_decap_8 FILLER_70_250 ();
 sg13g2_fill_2 FILLER_70_300 ();
 sg13g2_fill_1 FILLER_70_302 ();
 sg13g2_fill_1 FILLER_70_332 ();
 sg13g2_decap_8 FILLER_70_343 ();
 sg13g2_fill_2 FILLER_70_350 ();
 sg13g2_fill_1 FILLER_70_352 ();
 sg13g2_decap_8 FILLER_70_357 ();
 sg13g2_decap_4 FILLER_70_364 ();
 sg13g2_fill_1 FILLER_70_368 ();
 sg13g2_decap_4 FILLER_70_374 ();
 sg13g2_fill_2 FILLER_70_382 ();
 sg13g2_decap_8 FILLER_70_408 ();
 sg13g2_fill_2 FILLER_70_415 ();
 sg13g2_fill_2 FILLER_70_422 ();
 sg13g2_fill_2 FILLER_70_449 ();
 sg13g2_fill_1 FILLER_70_451 ();
 sg13g2_decap_4 FILLER_70_471 ();
 sg13g2_fill_1 FILLER_70_475 ();
 sg13g2_fill_2 FILLER_70_480 ();
 sg13g2_decap_8 FILLER_70_499 ();
 sg13g2_decap_4 FILLER_70_506 ();
 sg13g2_fill_2 FILLER_70_590 ();
 sg13g2_fill_2 FILLER_70_606 ();
 sg13g2_fill_1 FILLER_70_608 ();
 sg13g2_decap_8 FILLER_70_640 ();
 sg13g2_decap_8 FILLER_70_647 ();
 sg13g2_decap_8 FILLER_70_654 ();
 sg13g2_decap_4 FILLER_70_661 ();
 sg13g2_fill_2 FILLER_70_698 ();
 sg13g2_fill_1 FILLER_70_700 ();
 sg13g2_decap_8 FILLER_70_707 ();
 sg13g2_decap_4 FILLER_70_714 ();
 sg13g2_decap_8 FILLER_70_796 ();
 sg13g2_decap_4 FILLER_70_803 ();
 sg13g2_fill_2 FILLER_70_834 ();
 sg13g2_fill_2 FILLER_70_872 ();
 sg13g2_fill_1 FILLER_70_910 ();
 sg13g2_decap_4 FILLER_70_938 ();
 sg13g2_fill_2 FILLER_70_973 ();
 sg13g2_decap_4 FILLER_70_1033 ();
 sg13g2_fill_2 FILLER_70_1037 ();
 sg13g2_decap_8 FILLER_70_1071 ();
 sg13g2_fill_1 FILLER_70_1078 ();
 sg13g2_fill_2 FILLER_70_1121 ();
 sg13g2_fill_2 FILLER_70_1132 ();
 sg13g2_fill_1 FILLER_70_1134 ();
 sg13g2_fill_2 FILLER_70_1200 ();
 sg13g2_fill_1 FILLER_70_1202 ();
 sg13g2_fill_2 FILLER_70_1224 ();
 sg13g2_fill_1 FILLER_70_1226 ();
 sg13g2_decap_8 FILLER_70_1267 ();
 sg13g2_decap_8 FILLER_70_1274 ();
 sg13g2_decap_8 FILLER_70_1281 ();
 sg13g2_decap_8 FILLER_70_1288 ();
 sg13g2_decap_8 FILLER_70_1295 ();
 sg13g2_decap_8 FILLER_70_1302 ();
 sg13g2_decap_4 FILLER_70_1309 ();
 sg13g2_fill_2 FILLER_70_1313 ();
 sg13g2_decap_4 FILLER_71_0 ();
 sg13g2_decap_8 FILLER_71_44 ();
 sg13g2_fill_1 FILLER_71_51 ();
 sg13g2_fill_1 FILLER_71_80 ();
 sg13g2_fill_1 FILLER_71_89 ();
 sg13g2_fill_1 FILLER_71_112 ();
 sg13g2_fill_1 FILLER_71_126 ();
 sg13g2_fill_2 FILLER_71_140 ();
 sg13g2_decap_8 FILLER_71_164 ();
 sg13g2_decap_8 FILLER_71_171 ();
 sg13g2_decap_4 FILLER_71_178 ();
 sg13g2_fill_1 FILLER_71_182 ();
 sg13g2_fill_1 FILLER_71_221 ();
 sg13g2_decap_8 FILLER_71_249 ();
 sg13g2_decap_8 FILLER_71_256 ();
 sg13g2_decap_8 FILLER_71_263 ();
 sg13g2_decap_4 FILLER_71_270 ();
 sg13g2_fill_2 FILLER_71_274 ();
 sg13g2_decap_4 FILLER_71_356 ();
 sg13g2_fill_1 FILLER_71_433 ();
 sg13g2_fill_1 FILLER_71_512 ();
 sg13g2_fill_1 FILLER_71_526 ();
 sg13g2_fill_2 FILLER_71_614 ();
 sg13g2_fill_1 FILLER_71_616 ();
 sg13g2_decap_8 FILLER_71_648 ();
 sg13g2_fill_2 FILLER_71_655 ();
 sg13g2_fill_1 FILLER_71_657 ();
 sg13g2_fill_2 FILLER_71_690 ();
 sg13g2_fill_1 FILLER_71_719 ();
 sg13g2_fill_2 FILLER_71_756 ();
 sg13g2_fill_1 FILLER_71_758 ();
 sg13g2_decap_8 FILLER_71_795 ();
 sg13g2_decap_8 FILLER_71_802 ();
 sg13g2_fill_2 FILLER_71_809 ();
 sg13g2_fill_1 FILLER_71_811 ();
 sg13g2_fill_1 FILLER_71_845 ();
 sg13g2_fill_1 FILLER_71_860 ();
 sg13g2_fill_2 FILLER_71_872 ();
 sg13g2_fill_2 FILLER_71_904 ();
 sg13g2_fill_1 FILLER_71_906 ();
 sg13g2_fill_2 FILLER_71_928 ();
 sg13g2_fill_1 FILLER_71_930 ();
 sg13g2_decap_4 FILLER_71_975 ();
 sg13g2_fill_1 FILLER_71_979 ();
 sg13g2_decap_8 FILLER_71_988 ();
 sg13g2_fill_1 FILLER_71_995 ();
 sg13g2_fill_1 FILLER_71_1006 ();
 sg13g2_fill_2 FILLER_71_1044 ();
 sg13g2_fill_2 FILLER_71_1090 ();
 sg13g2_fill_1 FILLER_71_1092 ();
 sg13g2_decap_4 FILLER_71_1097 ();
 sg13g2_fill_1 FILLER_71_1114 ();
 sg13g2_fill_2 FILLER_71_1120 ();
 sg13g2_fill_1 FILLER_71_1122 ();
 sg13g2_fill_2 FILLER_71_1127 ();
 sg13g2_decap_8 FILLER_71_1138 ();
 sg13g2_fill_2 FILLER_71_1145 ();
 sg13g2_fill_1 FILLER_71_1147 ();
 sg13g2_fill_1 FILLER_71_1154 ();
 sg13g2_fill_2 FILLER_71_1164 ();
 sg13g2_fill_1 FILLER_71_1166 ();
 sg13g2_fill_1 FILLER_71_1181 ();
 sg13g2_fill_2 FILLER_71_1219 ();
 sg13g2_decap_8 FILLER_71_1265 ();
 sg13g2_decap_8 FILLER_71_1272 ();
 sg13g2_decap_8 FILLER_71_1279 ();
 sg13g2_decap_8 FILLER_71_1286 ();
 sg13g2_decap_8 FILLER_71_1293 ();
 sg13g2_decap_8 FILLER_71_1300 ();
 sg13g2_decap_8 FILLER_71_1307 ();
 sg13g2_fill_1 FILLER_71_1314 ();
 sg13g2_decap_8 FILLER_72_0 ();
 sg13g2_decap_4 FILLER_72_7 ();
 sg13g2_fill_1 FILLER_72_11 ();
 sg13g2_fill_1 FILLER_72_63 ();
 sg13g2_fill_1 FILLER_72_91 ();
 sg13g2_fill_2 FILLER_72_115 ();
 sg13g2_decap_8 FILLER_72_181 ();
 sg13g2_fill_2 FILLER_72_188 ();
 sg13g2_fill_1 FILLER_72_237 ();
 sg13g2_fill_2 FILLER_72_323 ();
 sg13g2_fill_1 FILLER_72_334 ();
 sg13g2_fill_1 FILLER_72_339 ();
 sg13g2_decap_4 FILLER_72_349 ();
 sg13g2_fill_1 FILLER_72_435 ();
 sg13g2_decap_8 FILLER_72_498 ();
 sg13g2_decap_4 FILLER_72_505 ();
 sg13g2_fill_2 FILLER_72_509 ();
 sg13g2_decap_8 FILLER_72_524 ();
 sg13g2_fill_2 FILLER_72_531 ();
 sg13g2_decap_4 FILLER_72_537 ();
 sg13g2_fill_2 FILLER_72_541 ();
 sg13g2_fill_1 FILLER_72_547 ();
 sg13g2_fill_2 FILLER_72_575 ();
 sg13g2_fill_2 FILLER_72_609 ();
 sg13g2_decap_4 FILLER_72_640 ();
 sg13g2_decap_4 FILLER_72_657 ();
 sg13g2_fill_1 FILLER_72_661 ();
 sg13g2_fill_2 FILLER_72_671 ();
 sg13g2_fill_1 FILLER_72_673 ();
 sg13g2_fill_2 FILLER_72_715 ();
 sg13g2_fill_2 FILLER_72_730 ();
 sg13g2_decap_4 FILLER_72_737 ();
 sg13g2_fill_1 FILLER_72_741 ();
 sg13g2_decap_8 FILLER_72_769 ();
 sg13g2_decap_4 FILLER_72_776 ();
 sg13g2_fill_2 FILLER_72_780 ();
 sg13g2_decap_8 FILLER_72_791 ();
 sg13g2_fill_1 FILLER_72_798 ();
 sg13g2_decap_8 FILLER_72_803 ();
 sg13g2_fill_2 FILLER_72_810 ();
 sg13g2_fill_1 FILLER_72_812 ();
 sg13g2_fill_1 FILLER_72_817 ();
 sg13g2_decap_8 FILLER_72_822 ();
 sg13g2_decap_4 FILLER_72_829 ();
 sg13g2_fill_2 FILLER_72_837 ();
 sg13g2_fill_2 FILLER_72_904 ();
 sg13g2_fill_2 FILLER_72_919 ();
 sg13g2_fill_1 FILLER_72_965 ();
 sg13g2_decap_8 FILLER_72_984 ();
 sg13g2_decap_8 FILLER_72_991 ();
 sg13g2_decap_4 FILLER_72_998 ();
 sg13g2_fill_1 FILLER_72_1002 ();
 sg13g2_fill_2 FILLER_72_1012 ();
 sg13g2_fill_1 FILLER_72_1014 ();
 sg13g2_decap_4 FILLER_72_1028 ();
 sg13g2_fill_2 FILLER_72_1032 ();
 sg13g2_fill_1 FILLER_72_1095 ();
 sg13g2_decap_8 FILLER_72_1149 ();
 sg13g2_decap_4 FILLER_72_1156 ();
 sg13g2_fill_1 FILLER_72_1179 ();
 sg13g2_decap_8 FILLER_72_1252 ();
 sg13g2_decap_8 FILLER_72_1259 ();
 sg13g2_decap_8 FILLER_72_1266 ();
 sg13g2_decap_8 FILLER_72_1273 ();
 sg13g2_decap_8 FILLER_72_1280 ();
 sg13g2_decap_8 FILLER_72_1287 ();
 sg13g2_decap_8 FILLER_72_1294 ();
 sg13g2_decap_8 FILLER_72_1301 ();
 sg13g2_decap_8 FILLER_72_1308 ();
 sg13g2_decap_8 FILLER_73_0 ();
 sg13g2_decap_8 FILLER_73_7 ();
 sg13g2_decap_8 FILLER_73_14 ();
 sg13g2_fill_2 FILLER_73_21 ();
 sg13g2_fill_1 FILLER_73_23 ();
 sg13g2_fill_2 FILLER_73_98 ();
 sg13g2_fill_1 FILLER_73_100 ();
 sg13g2_fill_1 FILLER_73_133 ();
 sg13g2_fill_2 FILLER_73_153 ();
 sg13g2_fill_2 FILLER_73_187 ();
 sg13g2_fill_2 FILLER_73_225 ();
 sg13g2_decap_8 FILLER_73_231 ();
 sg13g2_fill_1 FILLER_73_238 ();
 sg13g2_fill_2 FILLER_73_257 ();
 sg13g2_fill_1 FILLER_73_259 ();
 sg13g2_fill_1 FILLER_73_296 ();
 sg13g2_fill_2 FILLER_73_328 ();
 sg13g2_fill_1 FILLER_73_371 ();
 sg13g2_fill_1 FILLER_73_376 ();
 sg13g2_fill_2 FILLER_73_404 ();
 sg13g2_fill_1 FILLER_73_406 ();
 sg13g2_fill_1 FILLER_73_460 ();
 sg13g2_fill_1 FILLER_73_470 ();
 sg13g2_fill_2 FILLER_73_485 ();
 sg13g2_fill_1 FILLER_73_500 ();
 sg13g2_fill_1 FILLER_73_505 ();
 sg13g2_fill_2 FILLER_73_533 ();
 sg13g2_fill_1 FILLER_73_535 ();
 sg13g2_decap_4 FILLER_73_548 ();
 sg13g2_fill_2 FILLER_73_593 ();
 sg13g2_fill_2 FILLER_73_664 ();
 sg13g2_fill_1 FILLER_73_666 ();
 sg13g2_fill_1 FILLER_73_675 ();
 sg13g2_fill_1 FILLER_73_691 ();
 sg13g2_fill_1 FILLER_73_709 ();
 sg13g2_decap_4 FILLER_73_719 ();
 sg13g2_fill_2 FILLER_73_723 ();
 sg13g2_decap_8 FILLER_73_733 ();
 sg13g2_decap_8 FILLER_73_740 ();
 sg13g2_fill_2 FILLER_73_747 ();
 sg13g2_fill_1 FILLER_73_749 ();
 sg13g2_fill_2 FILLER_73_759 ();
 sg13g2_decap_8 FILLER_73_765 ();
 sg13g2_decap_4 FILLER_73_772 ();
 sg13g2_fill_2 FILLER_73_776 ();
 sg13g2_fill_2 FILLER_73_782 ();
 sg13g2_fill_1 FILLER_73_784 ();
 sg13g2_fill_1 FILLER_73_821 ();
 sg13g2_fill_2 FILLER_73_933 ();
 sg13g2_fill_1 FILLER_73_935 ();
 sg13g2_fill_2 FILLER_73_946 ();
 sg13g2_fill_1 FILLER_73_948 ();
 sg13g2_decap_8 FILLER_73_971 ();
 sg13g2_decap_8 FILLER_73_978 ();
 sg13g2_fill_2 FILLER_73_985 ();
 sg13g2_fill_1 FILLER_73_987 ();
 sg13g2_fill_2 FILLER_73_992 ();
 sg13g2_fill_1 FILLER_73_994 ();
 sg13g2_fill_2 FILLER_73_1028 ();
 sg13g2_fill_1 FILLER_73_1030 ();
 sg13g2_decap_4 FILLER_73_1077 ();
 sg13g2_fill_2 FILLER_73_1081 ();
 sg13g2_fill_1 FILLER_73_1115 ();
 sg13g2_fill_2 FILLER_73_1125 ();
 sg13g2_fill_1 FILLER_73_1127 ();
 sg13g2_fill_2 FILLER_73_1155 ();
 sg13g2_fill_1 FILLER_73_1157 ();
 sg13g2_fill_2 FILLER_73_1164 ();
 sg13g2_fill_1 FILLER_73_1166 ();
 sg13g2_fill_1 FILLER_73_1172 ();
 sg13g2_fill_2 FILLER_73_1179 ();
 sg13g2_decap_8 FILLER_73_1248 ();
 sg13g2_decap_8 FILLER_73_1255 ();
 sg13g2_decap_8 FILLER_73_1262 ();
 sg13g2_decap_8 FILLER_73_1269 ();
 sg13g2_decap_8 FILLER_73_1276 ();
 sg13g2_decap_8 FILLER_73_1283 ();
 sg13g2_decap_8 FILLER_73_1290 ();
 sg13g2_decap_8 FILLER_73_1297 ();
 sg13g2_decap_8 FILLER_73_1304 ();
 sg13g2_decap_4 FILLER_73_1311 ();
 sg13g2_decap_4 FILLER_74_0 ();
 sg13g2_fill_1 FILLER_74_4 ();
 sg13g2_fill_2 FILLER_74_59 ();
 sg13g2_fill_1 FILLER_74_83 ();
 sg13g2_fill_1 FILLER_74_101 ();
 sg13g2_fill_1 FILLER_74_124 ();
 sg13g2_fill_2 FILLER_74_146 ();
 sg13g2_fill_1 FILLER_74_148 ();
 sg13g2_fill_2 FILLER_74_229 ();
 sg13g2_decap_4 FILLER_74_240 ();
 sg13g2_fill_1 FILLER_74_275 ();
 sg13g2_fill_1 FILLER_74_294 ();
 sg13g2_fill_1 FILLER_74_312 ();
 sg13g2_fill_2 FILLER_74_394 ();
 sg13g2_fill_1 FILLER_74_396 ();
 sg13g2_fill_2 FILLER_74_406 ();
 sg13g2_fill_2 FILLER_74_421 ();
 sg13g2_decap_8 FILLER_74_432 ();
 sg13g2_decap_8 FILLER_74_439 ();
 sg13g2_decap_8 FILLER_74_446 ();
 sg13g2_fill_2 FILLER_74_453 ();
 sg13g2_fill_1 FILLER_74_455 ();
 sg13g2_fill_2 FILLER_74_469 ();
 sg13g2_fill_1 FILLER_74_471 ();
 sg13g2_fill_1 FILLER_74_496 ();
 sg13g2_fill_1 FILLER_74_514 ();
 sg13g2_fill_2 FILLER_74_542 ();
 sg13g2_fill_1 FILLER_74_544 ();
 sg13g2_fill_2 FILLER_74_556 ();
 sg13g2_decap_8 FILLER_74_562 ();
 sg13g2_fill_1 FILLER_74_569 ();
 sg13g2_decap_4 FILLER_74_618 ();
 sg13g2_fill_1 FILLER_74_622 ();
 sg13g2_fill_2 FILLER_74_627 ();
 sg13g2_fill_1 FILLER_74_629 ();
 sg13g2_fill_2 FILLER_74_639 ();
 sg13g2_decap_8 FILLER_74_654 ();
 sg13g2_fill_2 FILLER_74_661 ();
 sg13g2_decap_8 FILLER_74_694 ();
 sg13g2_fill_2 FILLER_74_701 ();
 sg13g2_decap_4 FILLER_74_722 ();
 sg13g2_fill_2 FILLER_74_726 ();
 sg13g2_fill_1 FILLER_74_746 ();
 sg13g2_fill_2 FILLER_74_783 ();
 sg13g2_fill_1 FILLER_74_785 ();
 sg13g2_fill_1 FILLER_74_813 ();
 sg13g2_fill_2 FILLER_74_861 ();
 sg13g2_fill_1 FILLER_74_863 ();
 sg13g2_fill_2 FILLER_74_873 ();
 sg13g2_decap_8 FILLER_74_913 ();
 sg13g2_fill_2 FILLER_74_991 ();
 sg13g2_fill_1 FILLER_74_1020 ();
 sg13g2_fill_2 FILLER_74_1041 ();
 sg13g2_fill_2 FILLER_74_1061 ();
 sg13g2_decap_4 FILLER_74_1069 ();
 sg13g2_fill_2 FILLER_74_1073 ();
 sg13g2_fill_2 FILLER_74_1196 ();
 sg13g2_fill_1 FILLER_74_1198 ();
 sg13g2_decap_8 FILLER_74_1244 ();
 sg13g2_decap_8 FILLER_74_1251 ();
 sg13g2_decap_8 FILLER_74_1258 ();
 sg13g2_decap_8 FILLER_74_1265 ();
 sg13g2_decap_8 FILLER_74_1272 ();
 sg13g2_decap_8 FILLER_74_1279 ();
 sg13g2_decap_8 FILLER_74_1286 ();
 sg13g2_decap_8 FILLER_74_1293 ();
 sg13g2_decap_8 FILLER_74_1300 ();
 sg13g2_decap_8 FILLER_74_1307 ();
 sg13g2_fill_1 FILLER_74_1314 ();
 sg13g2_decap_8 FILLER_75_0 ();
 sg13g2_decap_8 FILLER_75_7 ();
 sg13g2_fill_1 FILLER_75_14 ();
 sg13g2_decap_8 FILLER_75_19 ();
 sg13g2_decap_8 FILLER_75_26 ();
 sg13g2_decap_8 FILLER_75_33 ();
 sg13g2_fill_2 FILLER_75_40 ();
 sg13g2_decap_4 FILLER_75_46 ();
 sg13g2_fill_2 FILLER_75_50 ();
 sg13g2_fill_1 FILLER_75_70 ();
 sg13g2_fill_2 FILLER_75_75 ();
 sg13g2_decap_8 FILLER_75_85 ();
 sg13g2_decap_8 FILLER_75_92 ();
 sg13g2_fill_2 FILLER_75_121 ();
 sg13g2_fill_2 FILLER_75_146 ();
 sg13g2_fill_1 FILLER_75_148 ();
 sg13g2_fill_1 FILLER_75_199 ();
 sg13g2_fill_1 FILLER_75_205 ();
 sg13g2_decap_4 FILLER_75_241 ();
 sg13g2_fill_2 FILLER_75_245 ();
 sg13g2_fill_2 FILLER_75_272 ();
 sg13g2_fill_1 FILLER_75_274 ();
 sg13g2_fill_2 FILLER_75_280 ();
 sg13g2_fill_2 FILLER_75_310 ();
 sg13g2_fill_1 FILLER_75_312 ();
 sg13g2_fill_2 FILLER_75_376 ();
 sg13g2_fill_1 FILLER_75_387 ();
 sg13g2_decap_8 FILLER_75_392 ();
 sg13g2_decap_4 FILLER_75_399 ();
 sg13g2_fill_2 FILLER_75_408 ();
 sg13g2_decap_4 FILLER_75_416 ();
 sg13g2_fill_1 FILLER_75_420 ();
 sg13g2_decap_8 FILLER_75_425 ();
 sg13g2_decap_8 FILLER_75_432 ();
 sg13g2_decap_4 FILLER_75_439 ();
 sg13g2_fill_1 FILLER_75_443 ();
 sg13g2_fill_2 FILLER_75_453 ();
 sg13g2_fill_2 FILLER_75_514 ();
 sg13g2_fill_1 FILLER_75_536 ();
 sg13g2_fill_2 FILLER_75_546 ();
 sg13g2_fill_1 FILLER_75_548 ();
 sg13g2_fill_2 FILLER_75_562 ();
 sg13g2_decap_8 FILLER_75_568 ();
 sg13g2_fill_2 FILLER_75_575 ();
 sg13g2_fill_2 FILLER_75_594 ();
 sg13g2_fill_1 FILLER_75_596 ();
 sg13g2_decap_8 FILLER_75_611 ();
 sg13g2_fill_1 FILLER_75_618 ();
 sg13g2_fill_2 FILLER_75_624 ();
 sg13g2_fill_1 FILLER_75_626 ();
 sg13g2_decap_8 FILLER_75_705 ();
 sg13g2_decap_4 FILLER_75_712 ();
 sg13g2_fill_2 FILLER_75_721 ();
 sg13g2_fill_2 FILLER_75_765 ();
 sg13g2_fill_1 FILLER_75_767 ();
 sg13g2_fill_1 FILLER_75_791 ();
 sg13g2_fill_2 FILLER_75_802 ();
 sg13g2_fill_1 FILLER_75_804 ();
 sg13g2_fill_1 FILLER_75_811 ();
 sg13g2_fill_2 FILLER_75_850 ();
 sg13g2_fill_1 FILLER_75_852 ();
 sg13g2_fill_1 FILLER_75_894 ();
 sg13g2_decap_8 FILLER_75_904 ();
 sg13g2_fill_1 FILLER_75_911 ();
 sg13g2_fill_2 FILLER_75_923 ();
 sg13g2_fill_1 FILLER_75_925 ();
 sg13g2_fill_2 FILLER_75_958 ();
 sg13g2_fill_2 FILLER_75_1001 ();
 sg13g2_fill_1 FILLER_75_1003 ();
 sg13g2_decap_4 FILLER_75_1017 ();
 sg13g2_fill_2 FILLER_75_1030 ();
 sg13g2_fill_1 FILLER_75_1032 ();
 sg13g2_decap_4 FILLER_75_1076 ();
 sg13g2_decap_4 FILLER_75_1084 ();
 sg13g2_fill_2 FILLER_75_1097 ();
 sg13g2_fill_2 FILLER_75_1120 ();
 sg13g2_fill_1 FILLER_75_1122 ();
 sg13g2_fill_2 FILLER_75_1133 ();
 sg13g2_fill_1 FILLER_75_1135 ();
 sg13g2_fill_2 FILLER_75_1163 ();
 sg13g2_fill_2 FILLER_75_1171 ();
 sg13g2_fill_1 FILLER_75_1173 ();
 sg13g2_decap_4 FILLER_75_1208 ();
 sg13g2_fill_2 FILLER_75_1212 ();
 sg13g2_fill_1 FILLER_75_1218 ();
 sg13g2_fill_2 FILLER_75_1223 ();
 sg13g2_fill_1 FILLER_75_1225 ();
 sg13g2_decap_8 FILLER_75_1235 ();
 sg13g2_decap_8 FILLER_75_1242 ();
 sg13g2_decap_8 FILLER_75_1249 ();
 sg13g2_decap_8 FILLER_75_1256 ();
 sg13g2_decap_8 FILLER_75_1263 ();
 sg13g2_decap_8 FILLER_75_1270 ();
 sg13g2_decap_8 FILLER_75_1277 ();
 sg13g2_decap_8 FILLER_75_1284 ();
 sg13g2_decap_8 FILLER_75_1291 ();
 sg13g2_decap_8 FILLER_75_1298 ();
 sg13g2_decap_8 FILLER_75_1305 ();
 sg13g2_fill_2 FILLER_75_1312 ();
 sg13g2_fill_1 FILLER_75_1314 ();
 sg13g2_decap_8 FILLER_76_0 ();
 sg13g2_decap_8 FILLER_76_39 ();
 sg13g2_fill_2 FILLER_76_46 ();
 sg13g2_fill_2 FILLER_76_61 ();
 sg13g2_fill_1 FILLER_76_63 ();
 sg13g2_fill_1 FILLER_76_103 ();
 sg13g2_fill_1 FILLER_76_117 ();
 sg13g2_fill_2 FILLER_76_184 ();
 sg13g2_fill_2 FILLER_76_209 ();
 sg13g2_decap_8 FILLER_76_235 ();
 sg13g2_decap_8 FILLER_76_242 ();
 sg13g2_decap_4 FILLER_76_249 ();
 sg13g2_fill_2 FILLER_76_295 ();
 sg13g2_fill_1 FILLER_76_297 ();
 sg13g2_fill_1 FILLER_76_329 ();
 sg13g2_fill_1 FILLER_76_350 ();
 sg13g2_fill_2 FILLER_76_378 ();
 sg13g2_fill_1 FILLER_76_380 ();
 sg13g2_fill_2 FILLER_76_386 ();
 sg13g2_fill_1 FILLER_76_388 ();
 sg13g2_decap_4 FILLER_76_421 ();
 sg13g2_fill_2 FILLER_76_425 ();
 sg13g2_fill_2 FILLER_76_433 ();
 sg13g2_fill_1 FILLER_76_435 ();
 sg13g2_fill_1 FILLER_76_499 ();
 sg13g2_fill_2 FILLER_76_509 ();
 sg13g2_fill_1 FILLER_76_521 ();
 sg13g2_fill_2 FILLER_76_579 ();
 sg13g2_fill_2 FILLER_76_586 ();
 sg13g2_fill_1 FILLER_76_588 ();
 sg13g2_fill_2 FILLER_76_606 ();
 sg13g2_fill_2 FILLER_76_675 ();
 sg13g2_fill_1 FILLER_76_677 ();
 sg13g2_fill_1 FILLER_76_715 ();
 sg13g2_fill_2 FILLER_76_780 ();
 sg13g2_fill_2 FILLER_76_797 ();
 sg13g2_fill_1 FILLER_76_799 ();
 sg13g2_fill_1 FILLER_76_819 ();
 sg13g2_fill_2 FILLER_76_847 ();
 sg13g2_fill_1 FILLER_76_849 ();
 sg13g2_fill_2 FILLER_76_866 ();
 sg13g2_fill_1 FILLER_76_873 ();
 sg13g2_fill_2 FILLER_76_878 ();
 sg13g2_fill_2 FILLER_76_889 ();
 sg13g2_fill_1 FILLER_76_895 ();
 sg13g2_fill_2 FILLER_76_901 ();
 sg13g2_fill_1 FILLER_76_903 ();
 sg13g2_fill_2 FILLER_76_914 ();
 sg13g2_fill_2 FILLER_76_925 ();
 sg13g2_fill_1 FILLER_76_927 ();
 sg13g2_fill_2 FILLER_76_936 ();
 sg13g2_fill_1 FILLER_76_938 ();
 sg13g2_fill_2 FILLER_76_975 ();
 sg13g2_fill_2 FILLER_76_986 ();
 sg13g2_fill_2 FILLER_76_1004 ();
 sg13g2_fill_1 FILLER_76_1006 ();
 sg13g2_decap_8 FILLER_76_1026 ();
 sg13g2_fill_2 FILLER_76_1033 ();
 sg13g2_fill_1 FILLER_76_1035 ();
 sg13g2_fill_2 FILLER_76_1068 ();
 sg13g2_fill_1 FILLER_76_1070 ();
 sg13g2_decap_8 FILLER_76_1077 ();
 sg13g2_fill_1 FILLER_76_1084 ();
 sg13g2_fill_1 FILLER_76_1090 ();
 sg13g2_fill_2 FILLER_76_1110 ();
 sg13g2_fill_1 FILLER_76_1112 ();
 sg13g2_decap_8 FILLER_76_1198 ();
 sg13g2_decap_8 FILLER_76_1205 ();
 sg13g2_decap_8 FILLER_76_1212 ();
 sg13g2_fill_2 FILLER_76_1219 ();
 sg13g2_fill_1 FILLER_76_1221 ();
 sg13g2_decap_8 FILLER_76_1226 ();
 sg13g2_decap_8 FILLER_76_1233 ();
 sg13g2_decap_8 FILLER_76_1240 ();
 sg13g2_decap_8 FILLER_76_1247 ();
 sg13g2_decap_8 FILLER_76_1254 ();
 sg13g2_decap_8 FILLER_76_1261 ();
 sg13g2_decap_8 FILLER_76_1268 ();
 sg13g2_decap_8 FILLER_76_1275 ();
 sg13g2_decap_8 FILLER_76_1282 ();
 sg13g2_decap_8 FILLER_76_1289 ();
 sg13g2_decap_8 FILLER_76_1296 ();
 sg13g2_decap_8 FILLER_76_1303 ();
 sg13g2_decap_4 FILLER_76_1310 ();
 sg13g2_fill_1 FILLER_76_1314 ();
 sg13g2_decap_4 FILLER_77_0 ();
 sg13g2_fill_1 FILLER_77_4 ();
 sg13g2_fill_2 FILLER_77_41 ();
 sg13g2_fill_1 FILLER_77_43 ();
 sg13g2_fill_2 FILLER_77_98 ();
 sg13g2_fill_2 FILLER_77_109 ();
 sg13g2_fill_1 FILLER_77_134 ();
 sg13g2_fill_2 FILLER_77_159 ();
 sg13g2_fill_2 FILLER_77_178 ();
 sg13g2_fill_1 FILLER_77_180 ();
 sg13g2_decap_8 FILLER_77_240 ();
 sg13g2_decap_8 FILLER_77_247 ();
 sg13g2_decap_8 FILLER_77_254 ();
 sg13g2_fill_2 FILLER_77_275 ();
 sg13g2_fill_2 FILLER_77_309 ();
 sg13g2_fill_2 FILLER_77_338 ();
 sg13g2_fill_1 FILLER_77_340 ();
 sg13g2_fill_2 FILLER_77_350 ();
 sg13g2_fill_1 FILLER_77_352 ();
 sg13g2_fill_1 FILLER_77_399 ();
 sg13g2_decap_4 FILLER_77_436 ();
 sg13g2_fill_2 FILLER_77_440 ();
 sg13g2_fill_1 FILLER_77_474 ();
 sg13g2_fill_2 FILLER_77_502 ();
 sg13g2_fill_1 FILLER_77_504 ();
 sg13g2_fill_2 FILLER_77_564 ();
 sg13g2_fill_1 FILLER_77_566 ();
 sg13g2_fill_1 FILLER_77_585 ();
 sg13g2_fill_2 FILLER_77_622 ();
 sg13g2_fill_1 FILLER_77_731 ();
 sg13g2_fill_2 FILLER_77_749 ();
 sg13g2_fill_1 FILLER_77_832 ();
 sg13g2_fill_2 FILLER_77_838 ();
 sg13g2_decap_4 FILLER_77_933 ();
 sg13g2_fill_2 FILLER_77_937 ();
 sg13g2_decap_4 FILLER_77_959 ();
 sg13g2_fill_2 FILLER_77_963 ();
 sg13g2_fill_1 FILLER_77_974 ();
 sg13g2_fill_2 FILLER_77_979 ();
 sg13g2_fill_1 FILLER_77_998 ();
 sg13g2_fill_2 FILLER_77_1032 ();
 sg13g2_fill_1 FILLER_77_1034 ();
 sg13g2_fill_2 FILLER_77_1056 ();
 sg13g2_fill_1 FILLER_77_1076 ();
 sg13g2_fill_2 FILLER_77_1117 ();
 sg13g2_fill_1 FILLER_77_1119 ();
 sg13g2_decap_8 FILLER_77_1194 ();
 sg13g2_decap_8 FILLER_77_1201 ();
 sg13g2_decap_8 FILLER_77_1208 ();
 sg13g2_decap_8 FILLER_77_1215 ();
 sg13g2_decap_8 FILLER_77_1222 ();
 sg13g2_decap_8 FILLER_77_1229 ();
 sg13g2_decap_8 FILLER_77_1236 ();
 sg13g2_decap_8 FILLER_77_1243 ();
 sg13g2_decap_8 FILLER_77_1250 ();
 sg13g2_decap_8 FILLER_77_1257 ();
 sg13g2_decap_8 FILLER_77_1264 ();
 sg13g2_decap_8 FILLER_77_1271 ();
 sg13g2_decap_8 FILLER_77_1278 ();
 sg13g2_decap_8 FILLER_77_1285 ();
 sg13g2_decap_8 FILLER_77_1292 ();
 sg13g2_decap_8 FILLER_77_1299 ();
 sg13g2_decap_8 FILLER_77_1306 ();
 sg13g2_fill_2 FILLER_77_1313 ();
 sg13g2_decap_8 FILLER_78_0 ();
 sg13g2_decap_4 FILLER_78_7 ();
 sg13g2_fill_1 FILLER_78_11 ();
 sg13g2_fill_2 FILLER_78_17 ();
 sg13g2_fill_1 FILLER_78_19 ();
 sg13g2_fill_1 FILLER_78_47 ();
 sg13g2_fill_2 FILLER_78_139 ();
 sg13g2_fill_1 FILLER_78_182 ();
 sg13g2_decap_8 FILLER_78_240 ();
 sg13g2_decap_4 FILLER_78_247 ();
 sg13g2_fill_2 FILLER_78_251 ();
 sg13g2_fill_2 FILLER_78_280 ();
 sg13g2_fill_1 FILLER_78_282 ();
 sg13g2_fill_2 FILLER_78_314 ();
 sg13g2_fill_1 FILLER_78_316 ();
 sg13g2_fill_2 FILLER_78_358 ();
 sg13g2_fill_1 FILLER_78_409 ();
 sg13g2_fill_1 FILLER_78_456 ();
 sg13g2_fill_1 FILLER_78_462 ();
 sg13g2_fill_1 FILLER_78_476 ();
 sg13g2_fill_2 FILLER_78_509 ();
 sg13g2_fill_2 FILLER_78_538 ();
 sg13g2_fill_1 FILLER_78_540 ();
 sg13g2_decap_4 FILLER_78_577 ();
 sg13g2_decap_8 FILLER_78_649 ();
 sg13g2_fill_2 FILLER_78_687 ();
 sg13g2_fill_1 FILLER_78_689 ();
 sg13g2_fill_1 FILLER_78_717 ();
 sg13g2_fill_2 FILLER_78_763 ();
 sg13g2_fill_2 FILLER_78_792 ();
 sg13g2_fill_1 FILLER_78_825 ();
 sg13g2_fill_1 FILLER_78_928 ();
 sg13g2_fill_1 FILLER_78_961 ();
 sg13g2_fill_1 FILLER_78_1002 ();
 sg13g2_fill_2 FILLER_78_1030 ();
 sg13g2_fill_2 FILLER_78_1116 ();
 sg13g2_fill_1 FILLER_78_1118 ();
 sg13g2_decap_8 FILLER_78_1191 ();
 sg13g2_decap_8 FILLER_78_1198 ();
 sg13g2_decap_8 FILLER_78_1205 ();
 sg13g2_decap_8 FILLER_78_1212 ();
 sg13g2_decap_8 FILLER_78_1219 ();
 sg13g2_decap_8 FILLER_78_1226 ();
 sg13g2_decap_8 FILLER_78_1233 ();
 sg13g2_decap_8 FILLER_78_1240 ();
 sg13g2_decap_8 FILLER_78_1247 ();
 sg13g2_decap_8 FILLER_78_1254 ();
 sg13g2_decap_8 FILLER_78_1261 ();
 sg13g2_decap_8 FILLER_78_1268 ();
 sg13g2_decap_8 FILLER_78_1275 ();
 sg13g2_decap_8 FILLER_78_1282 ();
 sg13g2_decap_8 FILLER_78_1289 ();
 sg13g2_decap_8 FILLER_78_1296 ();
 sg13g2_decap_8 FILLER_78_1303 ();
 sg13g2_decap_4 FILLER_78_1310 ();
 sg13g2_fill_1 FILLER_78_1314 ();
 sg13g2_decap_8 FILLER_79_0 ();
 sg13g2_decap_8 FILLER_79_7 ();
 sg13g2_decap_4 FILLER_79_14 ();
 sg13g2_fill_1 FILLER_79_18 ();
 sg13g2_fill_2 FILLER_79_23 ();
 sg13g2_fill_2 FILLER_79_29 ();
 sg13g2_fill_2 FILLER_79_109 ();
 sg13g2_fill_1 FILLER_79_111 ();
 sg13g2_fill_2 FILLER_79_121 ();
 sg13g2_fill_1 FILLER_79_160 ();
 sg13g2_fill_2 FILLER_79_165 ();
 sg13g2_decap_8 FILLER_79_225 ();
 sg13g2_decap_8 FILLER_79_232 ();
 sg13g2_decap_8 FILLER_79_239 ();
 sg13g2_decap_4 FILLER_79_246 ();
 sg13g2_fill_1 FILLER_79_250 ();
 sg13g2_fill_1 FILLER_79_291 ();
 sg13g2_fill_2 FILLER_79_319 ();
 sg13g2_fill_2 FILLER_79_366 ();
 sg13g2_fill_2 FILLER_79_372 ();
 sg13g2_fill_1 FILLER_79_374 ();
 sg13g2_fill_1 FILLER_79_402 ();
 sg13g2_fill_2 FILLER_79_443 ();
 sg13g2_fill_2 FILLER_79_449 ();
 sg13g2_fill_1 FILLER_79_451 ();
 sg13g2_fill_2 FILLER_79_493 ();
 sg13g2_fill_2 FILLER_79_499 ();
 sg13g2_fill_1 FILLER_79_514 ();
 sg13g2_fill_2 FILLER_79_520 ();
 sg13g2_fill_1 FILLER_79_522 ();
 sg13g2_decap_4 FILLER_79_582 ();
 sg13g2_fill_2 FILLER_79_586 ();
 sg13g2_fill_2 FILLER_79_593 ();
 sg13g2_fill_1 FILLER_79_595 ();
 sg13g2_fill_1 FILLER_79_613 ();
 sg13g2_decap_8 FILLER_79_641 ();
 sg13g2_decap_8 FILLER_79_648 ();
 sg13g2_fill_2 FILLER_79_655 ();
 sg13g2_decap_8 FILLER_79_705 ();
 sg13g2_fill_2 FILLER_79_712 ();
 sg13g2_fill_1 FILLER_79_714 ();
 sg13g2_fill_2 FILLER_79_755 ();
 sg13g2_fill_2 FILLER_79_846 ();
 sg13g2_fill_2 FILLER_79_888 ();
 sg13g2_fill_2 FILLER_79_904 ();
 sg13g2_fill_2 FILLER_79_969 ();
 sg13g2_fill_1 FILLER_79_1002 ();
 sg13g2_fill_2 FILLER_79_1017 ();
 sg13g2_fill_2 FILLER_79_1037 ();
 sg13g2_fill_1 FILLER_79_1039 ();
 sg13g2_fill_2 FILLER_79_1076 ();
 sg13g2_fill_1 FILLER_79_1113 ();
 sg13g2_fill_2 FILLER_79_1119 ();
 sg13g2_fill_1 FILLER_79_1121 ();
 sg13g2_fill_2 FILLER_79_1176 ();
 sg13g2_decap_8 FILLER_79_1191 ();
 sg13g2_decap_8 FILLER_79_1198 ();
 sg13g2_decap_8 FILLER_79_1205 ();
 sg13g2_decap_8 FILLER_79_1212 ();
 sg13g2_decap_8 FILLER_79_1219 ();
 sg13g2_decap_8 FILLER_79_1226 ();
 sg13g2_decap_8 FILLER_79_1233 ();
 sg13g2_decap_8 FILLER_79_1240 ();
 sg13g2_decap_8 FILLER_79_1247 ();
 sg13g2_decap_8 FILLER_79_1254 ();
 sg13g2_decap_8 FILLER_79_1261 ();
 sg13g2_decap_8 FILLER_79_1268 ();
 sg13g2_decap_8 FILLER_79_1275 ();
 sg13g2_decap_8 FILLER_79_1282 ();
 sg13g2_decap_8 FILLER_79_1289 ();
 sg13g2_decap_8 FILLER_79_1296 ();
 sg13g2_decap_8 FILLER_79_1303 ();
 sg13g2_decap_4 FILLER_79_1310 ();
 sg13g2_fill_1 FILLER_79_1314 ();
 sg13g2_decap_8 FILLER_80_0 ();
 sg13g2_decap_8 FILLER_80_7 ();
 sg13g2_decap_8 FILLER_80_14 ();
 sg13g2_decap_8 FILLER_80_21 ();
 sg13g2_fill_2 FILLER_80_67 ();
 sg13g2_fill_2 FILLER_80_88 ();
 sg13g2_fill_1 FILLER_80_107 ();
 sg13g2_fill_2 FILLER_80_132 ();
 sg13g2_decap_4 FILLER_80_150 ();
 sg13g2_fill_1 FILLER_80_154 ();
 sg13g2_fill_1 FILLER_80_159 ();
 sg13g2_fill_1 FILLER_80_168 ();
 sg13g2_fill_2 FILLER_80_194 ();
 sg13g2_fill_2 FILLER_80_203 ();
 sg13g2_fill_1 FILLER_80_213 ();
 sg13g2_fill_1 FILLER_80_231 ();
 sg13g2_decap_4 FILLER_80_236 ();
 sg13g2_decap_8 FILLER_80_244 ();
 sg13g2_decap_8 FILLER_80_251 ();
 sg13g2_fill_2 FILLER_80_258 ();
 sg13g2_decap_8 FILLER_80_264 ();
 sg13g2_fill_1 FILLER_80_271 ();
 sg13g2_fill_1 FILLER_80_297 ();
 sg13g2_fill_1 FILLER_80_315 ();
 sg13g2_fill_1 FILLER_80_324 ();
 sg13g2_fill_1 FILLER_80_333 ();
 sg13g2_fill_2 FILLER_80_346 ();
 sg13g2_fill_1 FILLER_80_348 ();
 sg13g2_fill_2 FILLER_80_353 ();
 sg13g2_fill_1 FILLER_80_355 ();
 sg13g2_decap_4 FILLER_80_360 ();
 sg13g2_decap_8 FILLER_80_368 ();
 sg13g2_fill_1 FILLER_80_375 ();
 sg13g2_decap_8 FILLER_80_381 ();
 sg13g2_decap_4 FILLER_80_392 ();
 sg13g2_fill_2 FILLER_80_409 ();
 sg13g2_fill_1 FILLER_80_411 ();
 sg13g2_fill_1 FILLER_80_437 ();
 sg13g2_decap_8 FILLER_80_447 ();
 sg13g2_fill_2 FILLER_80_454 ();
 sg13g2_fill_1 FILLER_80_456 ();
 sg13g2_fill_1 FILLER_80_461 ();
 sg13g2_fill_1 FILLER_80_466 ();
 sg13g2_decap_8 FILLER_80_471 ();
 sg13g2_decap_4 FILLER_80_478 ();
 sg13g2_fill_1 FILLER_80_482 ();
 sg13g2_decap_8 FILLER_80_487 ();
 sg13g2_decap_4 FILLER_80_494 ();
 sg13g2_fill_1 FILLER_80_498 ();
 sg13g2_fill_2 FILLER_80_512 ();
 sg13g2_fill_1 FILLER_80_514 ();
 sg13g2_fill_1 FILLER_80_531 ();
 sg13g2_decap_4 FILLER_80_550 ();
 sg13g2_fill_2 FILLER_80_554 ();
 sg13g2_decap_4 FILLER_80_568 ();
 sg13g2_decap_8 FILLER_80_581 ();
 sg13g2_decap_4 FILLER_80_588 ();
 sg13g2_fill_1 FILLER_80_592 ();
 sg13g2_decap_8 FILLER_80_597 ();
 sg13g2_decap_4 FILLER_80_604 ();
 sg13g2_fill_1 FILLER_80_608 ();
 sg13g2_decap_8 FILLER_80_648 ();
 sg13g2_decap_8 FILLER_80_655 ();
 sg13g2_decap_4 FILLER_80_662 ();
 sg13g2_fill_2 FILLER_80_670 ();
 sg13g2_fill_1 FILLER_80_672 ();
 sg13g2_decap_4 FILLER_80_677 ();
 sg13g2_fill_1 FILLER_80_681 ();
 sg13g2_decap_8 FILLER_80_691 ();
 sg13g2_decap_8 FILLER_80_698 ();
 sg13g2_decap_8 FILLER_80_705 ();
 sg13g2_decap_8 FILLER_80_712 ();
 sg13g2_decap_8 FILLER_80_719 ();
 sg13g2_fill_2 FILLER_80_726 ();
 sg13g2_fill_1 FILLER_80_728 ();
 sg13g2_fill_2 FILLER_80_733 ();
 sg13g2_fill_1 FILLER_80_735 ();
 sg13g2_decap_8 FILLER_80_741 ();
 sg13g2_fill_1 FILLER_80_748 ();
 sg13g2_decap_4 FILLER_80_770 ();
 sg13g2_fill_1 FILLER_80_774 ();
 sg13g2_decap_8 FILLER_80_779 ();
 sg13g2_decap_4 FILLER_80_786 ();
 sg13g2_fill_1 FILLER_80_790 ();
 sg13g2_fill_1 FILLER_80_812 ();
 sg13g2_decap_8 FILLER_80_817 ();
 sg13g2_decap_8 FILLER_80_824 ();
 sg13g2_decap_8 FILLER_80_831 ();
 sg13g2_decap_4 FILLER_80_838 ();
 sg13g2_fill_2 FILLER_80_842 ();
 sg13g2_decap_4 FILLER_80_848 ();
 sg13g2_fill_2 FILLER_80_852 ();
 sg13g2_decap_4 FILLER_80_858 ();
 sg13g2_fill_1 FILLER_80_866 ();
 sg13g2_decap_4 FILLER_80_893 ();
 sg13g2_fill_2 FILLER_80_897 ();
 sg13g2_decap_4 FILLER_80_903 ();
 sg13g2_fill_1 FILLER_80_907 ();
 sg13g2_decap_8 FILLER_80_917 ();
 sg13g2_decap_8 FILLER_80_924 ();
 sg13g2_fill_2 FILLER_80_931 ();
 sg13g2_fill_1 FILLER_80_933 ();
 sg13g2_fill_2 FILLER_80_942 ();
 sg13g2_fill_1 FILLER_80_944 ();
 sg13g2_decap_4 FILLER_80_949 ();
 sg13g2_decap_4 FILLER_80_962 ();
 sg13g2_fill_1 FILLER_80_966 ();
 sg13g2_decap_4 FILLER_80_971 ();
 sg13g2_fill_1 FILLER_80_975 ();
 sg13g2_decap_8 FILLER_80_980 ();
 sg13g2_decap_8 FILLER_80_996 ();
 sg13g2_decap_4 FILLER_80_1003 ();
 sg13g2_fill_1 FILLER_80_1007 ();
 sg13g2_fill_1 FILLER_80_1016 ();
 sg13g2_decap_8 FILLER_80_1025 ();
 sg13g2_decap_4 FILLER_80_1032 ();
 sg13g2_decap_4 FILLER_80_1040 ();
 sg13g2_fill_1 FILLER_80_1044 ();
 sg13g2_fill_1 FILLER_80_1053 ();
 sg13g2_decap_8 FILLER_80_1063 ();
 sg13g2_decap_8 FILLER_80_1070 ();
 sg13g2_decap_8 FILLER_80_1077 ();
 sg13g2_fill_2 FILLER_80_1084 ();
 sg13g2_fill_1 FILLER_80_1086 ();
 sg13g2_decap_4 FILLER_80_1091 ();
 sg13g2_fill_2 FILLER_80_1103 ();
 sg13g2_decap_4 FILLER_80_1114 ();
 sg13g2_fill_2 FILLER_80_1122 ();
 sg13g2_fill_1 FILLER_80_1124 ();
 sg13g2_fill_2 FILLER_80_1129 ();
 sg13g2_decap_4 FILLER_80_1135 ();
 sg13g2_fill_1 FILLER_80_1139 ();
 sg13g2_fill_1 FILLER_80_1149 ();
 sg13g2_fill_1 FILLER_80_1158 ();
 sg13g2_decap_8 FILLER_80_1187 ();
 sg13g2_decap_8 FILLER_80_1194 ();
 sg13g2_decap_8 FILLER_80_1201 ();
 sg13g2_decap_8 FILLER_80_1208 ();
 sg13g2_decap_8 FILLER_80_1215 ();
 sg13g2_decap_8 FILLER_80_1222 ();
 sg13g2_decap_8 FILLER_80_1229 ();
 sg13g2_decap_8 FILLER_80_1236 ();
 sg13g2_decap_8 FILLER_80_1243 ();
 sg13g2_decap_8 FILLER_80_1250 ();
 sg13g2_decap_8 FILLER_80_1257 ();
 sg13g2_decap_8 FILLER_80_1264 ();
 sg13g2_decap_8 FILLER_80_1271 ();
 sg13g2_decap_8 FILLER_80_1278 ();
 sg13g2_decap_8 FILLER_80_1285 ();
 sg13g2_decap_8 FILLER_80_1292 ();
 sg13g2_decap_8 FILLER_80_1299 ();
 sg13g2_decap_8 FILLER_80_1306 ();
 sg13g2_fill_2 FILLER_80_1313 ();
 assign uio_oe[0] = net1374;
 assign uio_oe[1] = net1375;
 assign uio_oe[2] = net7;
 assign uio_oe[3] = net1376;
 assign uio_oe[4] = net1377;
 assign uio_oe[5] = net1378;
 assign uio_oe[6] = net8;
 assign uio_oe[7] = net9;
 assign uio_out[2] = net10;
 assign uio_out[4] = net1379;
 assign uio_out[5] = net11;
 assign uio_out[6] = net12;
 assign uio_out[7] = net13;
 assign uo_out[0] = net14;
 assign uo_out[1] = net15;
 assign uo_out[2] = net16;
 assign uo_out[3] = net17;
endmodule
